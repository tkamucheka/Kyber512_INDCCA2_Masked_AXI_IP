`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/01/2021 03:41:37 AM
// Design Name: 
// Module Name: State_Unpack__mask_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module State_Unpack__mask_tb;

reg              clk = 0;
reg              rst_n = 1;
reg              enable = 0;
reg      [ 31:0] rand;
reg      [127:0] s;
wire         done;
wire [127:0] s1;
wire [127:0] s2;

reg [4095:0] random = 4096'h0107089500180639032507240aaf0452022804a108ee028002b100e102ed09290b190852048304f80be104b206fc095601f204230b4903bd0c830583070008ee00c80013063900cf00e70a6e0a40035b057105c2081406ae0cd1081208fd0b7e0c4104a70a6d04d901050105060c01fd04c808f90076035602b006800cae000b06e308d5082301a509150c54014b051b007c0b650afb08bb0c4209ee03b90c7003d9003003a609890a20066503d908f3002d0c6a03b708fa052d0adf00d201c6021b0781024b04a0013006a0058a023e014604cc084202120b63081f06de0686024409670b940b5d0682011907ad010004a90b1c052e0bcd0b9b035809b105fd0bf40b2a00a3081f000b06330cbd047307b20bb407a202b704a9079407790bed033108440c8e02210b6a06a700ce0b8f07960ae206a0052b076607d7006a0a32042d06a709fd037808fa032b073604ab08e501c3002d062a00b70c89088b07b20754048a07c9099c013f041501f400c40290066f05be09b2010e049709e507fe0626075d0c190c3209c506d00bc10bed0680084707a601d70cbe08870c4f04a606b005670a4005440ad606c805ec0625050c073b06c707af018f0393000304400515008d03f8015b08e4098a032a0059027f055e0a8202350574026c01bb0acf036f0c2300380316045c03310a620b32098305ea092f0bb600ab0a230acb0959;

reg [4095:0] SK = 4096'h0abd08a7065901ef092d09a40b00051508d809020cbc02b6004d06bb021f07cc081b0987023b058a01a3038a07400b0f03d8099708cd082803a003cd009301700b4408900cea08d7003601a90b0b00220bc106d704c6037601380c180490070b016505fc0a59008d067c0bbd04ea08ba06550413006008250838007501640a2508be0c6b0aec067c02cb03610b0c06bb01480b7f037f09dd08300abe0a640b56061f031f0afa015404ba05f808eb0a5e066a0b710bb70af800da05810a6a030f0af50381066605a804dc004d0c1209fb021201ff0815012e084f070806bd092e0b1507aa0575040304da0c97074700790c84015f0adb06f8022c008603a903d4063703a80b170ba20af10a0b0c350894047d09de06bc02d508c10a63092b03c001c90657001a0572032d026c0aca02a9015909c10b4605c9032d07e3050f039808780ce607dc0763033005e406bb00fc01eb04d00c760306017308e708f1093503ed053f06a003080a82088b066008ba02d90c33016800d10b930231048c042a040d0a40039f043109870807035a00d6052006d5096e0bae0b4e03bf0b08042809cc03c40737042d00920bd0014308f104b1074a037c053705cb03d4002909f40b8f0bcb0703062c0a5204e601070c990a8a04c003e407d6004505d008c5074d007109e801bb017f0bcc06db0602070e016602a601f907100c380c3d055f0059;

// 09b60012064108b706080280005100c306b

integer i;

State_Unpack__mask DUT0 (
  .clk(clk),
  .rst_n(rst_n),
  .enable(enable),
  .rand(rand),
  .s(s),
  .function_done(done),
  .s1(s1), 
  .s2(s2)
);

initial begin
  forever begin
    #5; clk = ~clk;
  end
end

initial begin
  #10; rst_n <= 1'b0;
  #10; rst_n <= 1'b1;
  #20;

  rand <= random[4095 -: 16];
  s    <= SK[4095 -: 128];
  
  #10; enable <= 1'b1;

  for (i=1; i < 8; i=i+1) begin
    #10; enable <= 1'b0;
         rand <= random[4095-(i*16) -: 16];
  end
  

  // $finish;

end

endmodule
