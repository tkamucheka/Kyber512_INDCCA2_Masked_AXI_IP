`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
DGyv/e99m5LREs0VEi6Jl4RlcDAGZw9ScYtzsqID1kkVYKQb+tJyo/oKljjNla8cTngdwz+D72Ql
tHGdEFtbAg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
A5nVmQT4jX5rtOo5laslrLuf7jTnq6hJwnJfREZDyZ8Bl1ue+OgkVeisAxpBVI2fAT1pAn+QnHWr
0bUekWFkOjPCqNtghWYxZ20bUlSoJu/E+CFdyZAoe/z20Ug/FNmt1N5UIjvmc0VavCYKin+zuQtZ
rT+ZjpDCmgnaCR/uhGA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
SaCjWjj7WCShovAgcEi+zWlGnR2i0HX6RiLilkMc15YWkMWsX8eRaeHUUjlzBjhdPJ5HD1txSKS0
DgH2vQwbO1nRAbcr22JzG89qvDQ/uvpBWSxjMwAVZIz4riHIBY6mvJtJS4uEz3miDM5g2mKE5YfI
mtmwYzxKKQwOwL1Q3BugPIuRYIR3HSQOBq/no0l64+89qK46lTs6b5qhsoKdOHUCpgrGaCFVPox7
rhmcSBYdd8LmAZ9W41kHwNRcMH0l422XGyrc80pmpDqZUlQHAK+w7k82mPVUcvl+IVDGzW4RI01P
blCPA0pIgSkfuG0t2BnQqs2eF4aQy/pDlEICRw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pMvYbJU/C+WP4fgnox3tgW3NogGesSc0qsStq94uMKih0/YVeJo8jouzfwnQe+vQao4u9dhM20dJ
EWTVEF3u95ZLeI6vbrfj5fx4a1NlRmKqLt21cw/RB/H/lVgFT0XgMv921k/ZUBS5yGwT5Ve5dciH
f0IkS/8ERcnuZ/+W3nZPz2HLnM5T143mMV4OKShkWpn6nR9+bqS0sMe3AWXCET6mwRlKQCZQAKEf
2lbK7qDZf820jdndiCOTJYC+JYzbCatQi9yXkYQTQBAhYYaqWW8xYl0YhsGSHhZ3o3Nas8b+/097
2ETsglmp8hjyupk3l0hgBEFU3fQtcvpiIlLmRg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eJCjQ8EoJFQbooW8+AcUEn4z9WKAZNsV3jEceqBx1ZUeF4OCl1l+sVqRizSDh9d0h288Xy6590Oy
d8XKqZQTH7kbIW6Pcz6iym52ttGj9C4VmWBDFr3ry0x/LMFvbT3z14PISxUfez+fTUkaK9EvSCNd
eQBL3qex0w6mgPPrXFRQxIBE9QX7R6Mcfgs/d02PvYsN3e8VilxrtFQjRTr2jbMgdbZdCgfY2BG/
3vI/SveIGIdlac8Llom8Jr65mI/jrT1Y2+J3N7vFah3E494YglGPhngvuiX7RJw43yVMM+m21ZF8
I4oD1FOa3gxr1BchbAvZ42l8cQOa9gzF3+jjCw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YE2XCADVIy3Q3WKcZ2cfhXf0u166DNGuwZEGTKdbvfoqX5uMPeNCooFA0HoUjztCIK/VZpmb33Ta
c3JEknu+ugzsETMcWZz3eIra222trQX1V2R2hq1Q7FTyHANw1KliRagesNTD6xmRCmumbVvKlp2h
BGqQtG8FFkQPGyhmbk0=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GQQua8yHd/po5lc5tOkxup4W+r5iq0c+m4vDuy8ji74YsDtUczw7GEFX+KUSRT1O9yPBl69BkckM
3rV20MrxG4GOyXsW4ApcXrkJ/FE1mj8z3ZrsTyIElKPmtSPHbuICp+38ML0Vi0tnuLSXi39lRfAf
VnswEo4JBbjv8xHKLQtuWB13x09ikcPa5HLBDfBmx/o7lVNQh8gvTJoUjOckMVafNUGUh2oUQeSH
ilkDSsIVhLHSo1xW/x/PxAIOd7Onp363/oT74qmKxH7t9mkK/5Afy48xGGvTW1UHFbzJP9XRNSZi
A/PDJ6odxdWhmiGg9ZuqsmJ6ahHaCX+eIMSc7w==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 71392)
`protect data_block
s/JJIyRDRSX4lKq7oB4nbZhgmsHn8GffORCHtZArlQYxdz2HMlQOE/mQDot7S9xIRan3FOQNIkkb
LM3fcFZCkUk05BnyZJHZ4NK9UydNwnGH/ObMDpqMxcoXa+wnBS8Xl/hcxtAquw0prrodloo+G7PY
7X96CEEmIym/maqVhIWM1uGlTa3FDn9pwqrLuGPbPcUtMO4A66CCFNmR0nRvuWRqIf+Jis0JmJ82
adYSNXYb94wTnv7qh3aAAYRRXeJ3ZOO85wIW56YDWPx43KsfsrR2/sBfIQQ1p9Tc6iT7WuN8RSPe
5sGcJ/RA1w9q1Pvzclra4ePe8gCloRCMOOt7ETI2FXAcWpE3bxI7neA3WdVu1yRZh2iU3NpKukGw
TMGzCEgZXPpMpw3XDG33fXuARvSf5i2YhsRYZOHPz1DMLzsdfKgw2VkyLqqrXJ43lPYBp/3jkKsU
aMgGhEVse2vIXFGrgeGW5OAjW/xh+bl/TWRbU+25UqcaWVo9+/lbb+SxclOegTqDqj6ATL5ZrArF
1RLwAEUjhtw8aJjUEusEHrnMqAmsba6Y+7UNHlNv92z62nSgXN2pfkMrujzI+0cXuV1OdjATBdtv
R7GLVpadMpzRP4PZqMsUBBkr69jRjaK1U1FM3382HDkyhd71JqLT2QLJ5sR14nQDBJYQZvR2Qxo8
h9joBhixPsjKaynjcbO19XRBUXizhnZG7SS8hrW6lUNJeDZA2u/Mc/fP3RERwoIhfOGOlSA9piur
hXWF07f85YB9YoiAlJQAyrGUfcYh+vv3rBYZmeSy3rkhiXi/x5OPRfuKWC9LEFpDAL9Hq+cEVAGI
5sw7j7U46rAUklr+Ani6vGSAXr3zgUUAgWaWW0+G6/Kz0Yi4Q3ctZXdIXLNmYz6Znn6mU1kjU6iR
ZMB4kL5RPNhUaS5XTN1zYTc3a77YTPCmBnWougnz6FAC5BsrY4PuWDQoP/K+3dybKkbiYJ0ChhXp
W/LPyWMDJt9oXWB4/cQ8irxpE+rfyJ/Dg2GO2bflqAK/AFLpgdmNy30fogY4frSXwM4iMTXxRf7o
7/uvFqzeWyigjrTW2zbwWAD+HHQm8IpBnb3IYkFc7RMD0HoJ3/YE5etTDLnl1ZoYHAO0/l5N46Iz
vnmPsK+0za2BruYOFJ3t6coNjHc2mUFo/Z1rZgj6PA68WvTmOCaaEXVjz7KS17Jwjfycuifwg5HK
kidj2qVt8jM6UJ7bkxQrwps5U83whsve7EPS7Fn46OjE4WSfCjzCSp3AIGTWQe8zVg0wkHlfG3Q/
aKy3nQq6btEPnZxBZS6tpziUiMwVXOqmN7IUy7+T2ofzY1JOHQOokcaWr9q+HYnrlmSjzLZQWlsf
nhLrGE3lBKIAl19gAkx/KeT7/AOu5iID7tlvOYq2f2ipiS4kNZu9PMktev5TIKczIKPXG9pbLRz4
1jkwd5utUgdEVj2Vr/5a7XNhdfe1zqLWZ6rYhUcbTk8CHUDqIAyP772nPff/gNEQhlPQBfYJUgZo
LBl7t4RsYTbDmuorBJg2BcSt1vo7q+a8/+o7wFw8zUU5/Vclg3atoKj38gW6/48xFTldQD2qRZKu
+fU1+4bAxknoW/ebSE6xljQGTF39OqLdVyft2cQzA5kMX3p77emKkIwaZfyDhTEcnuSGczcfBz1f
ivKdi6uQjaIltjZraI8iUOxBHkrNsRll9cbF/FBTcMn3++TZOzLrE4Hx+nZs8xrCbXvcKEpwf23b
NTRfhRrbpxAzWZXx/TbBMuhG592TJ1lmDJfw7DaCQOkgY4C6+MMkQ/W46v5fS1lZmcQyBcfAjUra
wEffFgQi0FGHSZzRxpy4wzXLd6l4TFM5O7gDRbqQvoJ5KVgcST3Ztqu2siwnCDrOZf8fQuzRXKMw
/rpEpdmW9q6f8f6Pxuzo5cZ5/6yRbWXgQigMHrVnaZ/7e6areKE06IW4JHwaOkoKlvu7GcEYcrEO
cOYkxJHo3RzF795a4SdIy1deRMAyOs5aS8nKIMRVZwDPt2YLpL0EBmyVu7lHVjcOTCN27GiPl4QR
VS5r45G8l/Kt0BshTSqo7MRU42alpXtKxXCG/hA3jjo2OJhgOvv+WVFA8WqAx5k4UqBVaYSbnSIR
fXxFzqPFYzK6zRmd1sc9wIZsvrnagNmxKl+w4MF8z/VDue3P2oUjxnyVC2In55lJ8yS1mQKxm0fV
MQx27+cQo2UH5SNj87/pf9fSxQF8DuPpTzkQd027kjSWl4ECo5/asG0IFcwauD1mzNuX3SYW56WJ
a7h1wwCmOTS4qsgyClwLHI4RMoDaSmK1aduYGhtIBqYbUKQ889nJ2FbEqXjRlRasQl9yWFfkKRq5
zullDvusLe/sCVTDMUgHzPPnpX0csZpNL9zvIXWv0FrgzBM2oiRuxcpVcwd84wf3mvBHOoKi/Xke
fXySFubmuIkwcnLAeKLmUbQadTjs1Q47IFByfpODuWC+WDPEbbK823FxSvT45PpB/OZdObZPBhmL
uHXL6EBZUEdrZvtCopFW6Wk7jJpWvzKYAR4jEX14sffrARzkPOS8uiYk7hlsJFms81klTEWYswz3
93E7LK/5kmbjWOf4D9lm5Q82Uvw7wECrYGG/7C/DSAtlsjcQ1NwzP3MAL5SfeFePbJ6t1KGP8VEw
g4SzZdIKda9yMD3MDzVcqzHKLjxbhVTX/nrPVgaI2xHm2rO1eDv6G4KSvaAWZZ3dtI3GzviSlpuI
U4R7h/ff3hwm5mMFx9MAlE3nm4O9MPC43FRIEUJ/HLlC7aKy0AXklqEGONCIY5/YeAVa6MHZsRcO
YTflYRwMvHCCig/qM4EQKyah1iqLTw8nVcku9EKO35WaoYd4yYRCj1ddKmIH+yZW7QMG0okZblox
5G4ObxLaFQQRGxkc7X30/nugopk20AIAaY/kesvp6ei0XkBuBIx50CNR2DY5S0uO2eYHRenQjjKC
lnWzSsoZ07oCF++HsDl9Tz3d5goNAEOxO8BP1BGe689+DPN1ScPLd+i9WBTaga6wwNz0vSyBujWc
pCRK69Rv9DGKPyV/05Fb9uW5yJni0er1jWtqKEsIRVrbmkhIQFlIFWYoB9vdfyrDLxQ3mvuiX1eg
4wtYVy0P9JdrcexlMMKz69HhYPE7EehH6cjZql8fMTGSLr2CLnVBK9xqG+dbTZuKw9peDp106+vv
amL8+N8BQvqmRSyQcSWSaWkeY0yeOI6Y8LggMXEdw7TaafnO9bZFEG59cKDmx9RAxK9skk5hkpoI
AbOaFxcJSlnUDnU7ciiz2BsJU6UykP1FMLqJsc3ASQKzwi2VaYKcu90OhnE+pZyI/O941E0IfhfH
hjO/m0tjaMmGpIbVSglYfnl/ggryIcuVzSaC9vht3Ql4XsGevjFZbQSN/6VX+/V+2LgiN/sDDGn9
EQUcBmp6HiYP/HrCwRU5r3AX5Bh4dFfRvsyj7kAu3FVcLQpompdImJ93BXCigPYZiHZziLORF7KG
TvvoTC7yrDRZpeuxWlu6R9KM1Ly7YCkvpt0UxDxy4FZwzjTJeTRnqkbbsNxXEwNAQ5Q89wsYBBRK
xObShQbI5Owv6E0Ae2brYdHI+TNMAvFi6SQoAVqgK/Nt2M8znBkZqu5paFd30uXpgsVhjuvWINXV
RFceiha0F4DxL5ffhrZi2JeCrJj14+8CjZjydGsMUhhECNDnmw4kejFCidvxVlUIUYG1l4mYp4ty
q8qmhZVMntJAefaT4RMacfQCW0kwK+CWla/rDzO9OC1gch+BYF/EGF9TR1gSpeH/x3Ph1sCdnlQE
b1umZNMZVL1Nr9PsHKe7yomTP7D6IZBgv2MIKLCjadSbAKHBZe82aP8aIvhXj5Zjs5BJV40ywV6o
ZqansVnwYiz+OZMJ+PRAteuy30tXw8EZOjEFr0pGqgDzbCR2nJOiPrGEaIelWZ0YEsK6gUF2+Cua
h2t2WbqC4NJWFUOQ4QgeXHWOXWZi9hP/CEQWOiQOW6PMoz0TO/tG78LZfEHpbbNgqw3ibFY6e7lL
wByhBT+hO0beD+V1T/fWuPlOmJLT9+/CFMoPpkrGzQr4sNLRh5ljRW37sb0UhrYY7sKow9MCkwzH
AikCxd0WCyTSR5ICY3aaW4oyJHaosbCwvh2Y6Dl5WlAB7mtOO9MOEioUPVdsVTgbI1PyyrOoltLa
3lu6vuepBEI3eSAe7zG+nwgHk9tktNwK4425Mg+gBou6/lTI8X07bsmL6CFK7vsfTDAMmVJaN0Oe
Ql/UBEu+Z3TR7GJA19y/6ukugYlQfQl9DlMKPIYWB925qtOfaXh8sfXoFqBnT9/Lkw7/fJLcwDoL
agVFPokOu6/3yv/7y5N6exp+NepGYONCTpiJ54AMuAUo+5FAkuorivtgr8yUsKuTfUjHUY3PpdM/
cPxfSP7N4ey9O4kx0iNQicGHWia/KVHtCP3yKpyDgCdRaTItlcZfeSicNPLdbGVfjp5wRXXKi70M
/BtiAxgWCMjqf5gMFQDl2hTTVJ7fde9MMuhZo5lXunFvfeNiDHiWjeC6496hStqzCTjFwgRxB/t2
UFF3OnlWgvh+YziiiTieZI2F1aagiynFxESDj4vkx18WHbsWJFfeaFRZa4QGyFoDBkDkADe+CBN6
1gE9TeVWY6xWS4j39XY/Usf7CHDhvpgvM+9+1b1UVtLq75e2QWWDGwnbl30VvNuQQFUjZAuQ26cf
Az4LFo39nTzAcJEFKpKvGTUbkuJ381HWgp0HEbXXM4QwuqaduTP/JfHTmHsUaiYBW/aNtTQLeJPn
c0ppejetTPzbh7QvilCN6E2ftEMued1EYKm5tWSo927XS6AkKORbYm3SHRoueTg4A4BDvvoxSssO
ieeyyYD/KoH5gn1zMV8Jbd4849ydPVHEKLDm3+ruBOm0XGu9e0uTeQ5GQVVIrE1VO1B9TCkeecXX
vBT3dd7rypSO0w9yZy9RpWnZgugJja29wigofda/SIgmUu0xbSdqRXXbB2x90ieyYWwxNGpyNxp7
Ywq8bUS3+vLC7yw/RlPVNOxiUpMlZqXjpcrbKWYryBWBkL0NNhg14wwois/OII1GtqosG1Ii1bCa
THqiUGykmaRsYg1Vd222BNEa+brogQOH5HMaqX10sc6A7yFNAwmJ0fvJ8mga+2a1RiyZ8NcN9WYi
nvQyDO6aCb3MvPU/3pQKRsKSx1CYn2K7URGhFHvYKWXoRIWPw9pi7Sdx5rRHtzGaHcqFXs0ARRC2
NNyZeUTZHbKcOVcOMPtoHIazWGdV3C03OkPyMBw8f70TBcMVEDp6e2BQdvK4DT5oLvAfSjqM48Dc
kpQVaF25qq00cUocMmtxWF5Z/Jt2OzQtM6mHHC4LRbM3EvaMsFkrmGGOP/SRVRBZhiAJbL5tXG1j
F+7/JaV5QEhPtGlenmztOXFHb5henNhaPzfw+2eQWVmMDq5W5sm5+t75p/Y7OsVw9rWb4rwkPtcV
WuqJZdMIO9/kvb/KQf//7LBOANJrVc7Y/9ih6sC7Gneme9eZn45HLJfAeiiLHQaInVv4D3X8icgP
S/aRlQqQx4shuecml4TQIYxCzTKstLztRPY3gvcwvAnFUNOqwRjMt2j2kK8EvBhyIuVXvpj5T5gL
FK+a6x42Bc+0zpc49vgNQOTBOqeArJfKS4qjwRba+Veukz3HLGtVNRBxD1KbGHR0/bRoaHa4HaN7
teKegNkKAVP7ykCJqxxtSwerJiVJs25ArwFPuGnkjwXZuFPQYPPh2kV0/zheGRi1RTWv76GGnCbZ
rq0mq919+vndDc7NT6i7RMEMGiRVgdPKHlvCxujZMbCVLtgpV/DAdNHmnQJddwUGrx0y2IyQw/IG
VjQDtCQFQ4ZKz0XzGqMU9pSwwllVdER/8ZY9d8l1dEyyv6HpIwu8yUdQ89S1wXKk1D+kX1uFX7nX
nddfV0ptL3dmK76pHPFzkFvU9hRhtKjPf4Hc0CMHKaYxrAaSPfzAk65qkVuvatABp8G6vlh9dx+5
uxbcsAlfxMeO/G9KXoZraVfCgzBq0lzVQ/Q4yOYA+2vGXYQG1BdTS71sZHi57ZiTjbrRfIyjWr4Y
eI1b0is7FU9TfSzae5V5H+GTJ6KvvVegFELa/H3zNO0kObcu6+d6cHfhiftTKw/lnIhrm2iOxPxP
jpADBfcxQaAdCyg74/2W4vTIjCNDsHi4oBRTabu6PrhovmB6Vw4/kLrF0jKz/NR1sPMZEqs6Ed14
vZtOjdaEx8ZsVoptBil8xXGbmHSFLIOL41LwImBuIFG7gDo2hmGLGqqS/Beesknj5xOy2z3J3JjF
IBMYgY9pThp3Es/Zbhsf5FVRT78RJ0qngaIRZJDNuJyOwi+pR9MU+Qo5956t8bT2UdfFKLj1mekb
J5metsq8LLmd9FGEt2OWjR3hppBN/XhOMOTSnAz5vMLMVTdiiG1dQvgL+ihSis62zA5GxRRc2pc4
MzTr2xhQuFtZdWW5NZEcw8xpUC7Ul9glZDudnOezLv46TrsCqaatKaFUjgwJKag41o61vfK5GLBO
zxSsbXD3I7aLDIb7cdzDp/Xu9A7mA6PkJbAsCsIhJKUaMd2UoYOaOTFzbn42KK1Xk+NwzA5aqutc
/LEr5RxyKqMbbTQQ07aF3is7smuaAoHEsmLqsy1mOoT/4MB8nFIz9kImLtiTU0dDbRZveo0puUpe
i+iWBDXC+/TuNXgF5ZbPW4hC3/f1mKV8ZdGmhp0WjKGBc5b6brxTWu2QPBbw7aqTJ7JS1Zm6x/WX
20cB8uuWOBxtljnYcKqYUfW4+J7DmwNWz/K7YrsyAcKRydIWVkdIEJ5KKAciykHE8kxAkvOUtaEa
DZf1KnnVuxGBl0ghbXmG/wFIsbTnBkIxd1ZVOkAWDpZRozrDSb2UrknYnk5Wca22Ms9DfXvNNjbZ
ouXGwErAeq0EgPOshqR1YhDIqEhAllrFzE8wF56fLoIdnN9V/SHzO79v8udklODOCXEIlChyYt+k
9t7UwF/ydBz3Pze3Qr/0IO8wo8tQoLMb1U/ZT/HdFTEedhhTERY8q9qsBHLtqfg05kY4isfWqdM2
QKLogVnnE5+UU/XlhbpzokefzVw9mJdeNTKNw5woLcv6OuCI/if8lqyUXToFhkwLPqxxXNy8bb46
SUFUQ6DAoKZ2kpu2pDWd1MMlpuTVojN4CVFO2zfFyFzs5oxPGKtgwKXKpK2fIItpCtJ+UfvnHadU
z6xXOMnlk+dJy1oqsfiFXJtG2BwSCGxGiJTRvYEejxxEufSciqoRyZKaY/bSUcT9BjhLwifwSdw3
mj+Ncr1Bok5quSLjgW+ykAt3WiCSJrdLNXfj/wkAkb1fQZjeMORdD7KZmAGnGCmD1eDQlTRAqOOo
z+Gc350+jEqRFeF5QIWtEjPRMUDFOcBC7CW7h1IcsshzD+iKY5z1RwS3mWbGUxAaWDWKUr/lpS3c
WxycGaZy/nh6/FqmdmxTJNzumJiYCnTPj9MV0VpHcUZcuiLd62CzoyVJyWUP038g1+7dcl6hv0vA
LH4Z1DxsP8ULxEG2FavF7a+B+EE7sdtpPQ3r3npBu+RXqralkCGpFhg45TlQXymcy7MXwjBYO75W
GKjM6b0DcPoWPlJFxoFUoTGqBxHX7ADryi18UIQs2Pm2tGTMbwHN/zLxlA43aH8Qaxn7Kaekl4YH
8ECgEQW0L9gaL86O8qA+q8ypRcD2Ie2xYecgLwignT6Bgq7WXLZgb25558zMJcYcQ05QKdTj5bbP
JTmcHVvLNrdSsHBwGUhI6mnbeGjtfCvSKS+nvLnqgEqgcwPxLne8GdXPNqR0R90Y9gh36Z+g7EMh
COUHCLKq9YRI3hmyEeSowsL3H0wUUdKK+MSSZTagCI7aKvdOkh54jkwb9hElULyk5Lv3ZzwP2/Gh
BT9b3o+2lBPbNzRUQ+TaYgx/Brs45haBuPufp4Zji7BBl7ahVkW5ULXH8tYfd9+APKMKSQR4Dos8
RZKJ+FYTYXyVY1m/3Ow50TAovxcBNjW9o39vEcmguJZMIMNefrPBJ3Tk55ePzq6mc2iJ27ZVTptb
sgx1ZlcOhueRrYKR3LOovVg0p7oe4WNDAS45N0ZjKTY8z6WPlj6UZQdiaFUFf/MyPfMYUQXAhmFL
GppSmA4EkOZAQAaQHaL/wEr6Yj5hEvyuDKV+snX7nml3OJnCGh7KWaRSqk4wWJHLhvLz9Eam/Rzh
BxdD5gBHl5OgkNpO/qx97/YGMu4jKoA/3ChZetJAfBvn/NztK2PalRTYS5TgERdLZxgclw0JVuEU
4L+8YLoHVbg/VfueOQW9ZCeaEEhxk/4CaxAGAJH63pYAcuS2K4B8gmWps7c3B/s9lJ0G8leX0nmF
YzpM5CMJ5CpuVpkJ/hFZ8lks84GxWLQzPXif6blLcqvxgVUXiD/7M+c+tnYRdum2gb5wf4nIEGSn
tfzJWPhX7jvVPezdjNpwUeHgcQL2mnjYhgcgCgwlCV9MPpyFEAsjnYLGQInCcf23JslRypLqwSEp
QEtUPkOG9Uj7sSz2vXrR5aUOOKKvg8vmy3HbHQVI2IXQujxR64ZnCkchmbRNYxNmne1mAjQZNv66
2a/85HfvrBDFarDALvMamiAu1Zi4LKyGqzA+ffuXq/6CRJ/UudH1LvvwX0KE8Mq9G+AYO4lr0TB9
eP6sAD0IjkwvGGkuGArP3+sTyj+0qMkzxES3Ms/oJIhJYbibUM1PgBO/dPTFOAsuKZ+4GPeYwfkb
B958FIcU3AU4JMPhfVgIRK8k6EPh7vQJPMhQoiWqkkBx8hTabF7A/UEOWj+5CGzbsb46Q7zME77w
wn7UjPryOjv4OpSUHYUDXwo+wXaxsKCrJa/wx6MGFnHKi3nwQHANdYTeOh6lkZ3uTyiwgwiLQzBV
qaxyJSA7WispNGQZbiD1E3IVC0RUZuvPL6TcuzpHDeAAmXc7bQlxahysi4B4/+tXly/JXlk8+p0Q
Rewii9kB+xGHvKZLlv/9eDDnClcciGMPIksdYcD5+2NtJTcjHMC02E7FZIgw/nKNZlFek+I1hqcx
iDKKZU2bVkfdQkOaa5hegCW7rO/7ZlZkiem8RIYMlcMutcDrT/erGJEP+euvVUDXbIpC+EylV0aj
0U2FDOBO2iOtO+51y5/BaNibLsSHNpNiO4Wfnup0/nbx8wp64i/nGTiyfEY1hwXOgbsiXJocNDGn
ptgipqMpCcFhZPBhwDFqDAAE8q3nPRuzPTR3mxva6YNARO0mzf06vKDFb6W6X1EBHbi313o3qj7s
EblP0UPU8vDSfIaYBBPZreGjU+tomUyb8mxO6mb6jKtxlMJWC2VzrxVGK/VlO0E5yWahNAWHLC8W
Tel9jz7DaNN164NjSIY1KDxNphHuMwXyIkR4eEYH1lT9ulOkg9U5x5x5QfIF6XlcQ6AeGMKqzm+N
fJCLAjo2oIq7X5qmX8mT5HBtLBxTDrxhUk4QXsFWhDPw4ul8LVD5hhRQiwtuGnwUMjFkZuE9UUf4
wG5+km01sW0mewUE81UH6ferG41Ictam5bN6W9E/WY2LBKt/Mz+hmFC4MwLU/fvAtuceGUVA9Nn6
zv4cftdMhE/GZg60HVmu2JQOY1aqFNlPoL8mYeNkMyeND6wYeX4IO+rH9blZebSp8UL3FqQKyoaz
J+mGOfxgieO6FL2QY922qTCP84eUiIwE/2D9O8ekB26NYZXs3Uz2i2CChUy8Uv+pU5tsJMRJLaV1
dHTJFRgtthD5D/ulD6AVXg6PstW9hL4hY120Za+Uvq8qgYXrsnd04nQf1hVB0hmCEv4xe1fj8w0r
O38/lrYG+FhMFGMEyYCp8732WjhNgftGg/DcMPgxPhPZbVntCGB+qt9D0Aff6GAiSVX3gVCFPW8Z
TMpeoDTFVQ82fHZUA4t59OjBcDyr0Rp8DxYlnZr6uB/7LO24GFskF3swfAQv87Bd2w9QINtONrnT
1YLW08qFfwR+SSjto4pVHub9cv4f5l6lVv/4rmALbNfkm8i2X2HCmwUxnXaraM6lHIk2RlAeevL7
Sv603oxa8h0iVGoUw5MwVIhNAWRZknEFmPWgFA4mNzJv3H3Tx4JU1+wzet14lm0dkM8FQNvLZyO+
4LL1n1kbHeouPRODkW4u8A1IcAhYbhlK3/0qxoI7nrInPdkqQp3r/H5jBjNLZmCB2/5VHlRFD5+h
0IWH89DNbzHGLHDG4dYpBra21iTwvzN/ZnfSbZ+fgQsBj6b0Om2hmo1cysDtOviJMhJTW2gGhzuB
jUakziVGEMi+2MQJzFlTgZptK/pOWHBK3hd9oVtuWYg8vIdRl704BefLmxxdRv9TPb83MhjYCsob
x7cwkoTNFWXgnnQFlz5A7YEb/+CadVp4ZUznMu8QvuyozkyVrXvgaJJIGhkddhqkoMFMYyY0mtOu
ZfmvuCkToRPgX2OnsezHmx9sDJYe20p+JLWL2YrD0We50Upjrb2kRihEbfTiP0Pw1XMw3w3uWm/X
C8SSy9VkZywBNQ3GO7faOpgf0sosVNK5l2UtqQwZ9IqNAQQS/jPB/oNKtF7CqL90HtlJlHVKx2pu
T41J98CFAhpCeQ2dtuKpfvcXBVCmLpXBflW4qyeocPFrcBXeLB+IATxZo5x6cUjP8SpBv5RKbKx2
jWzlgV5ezCjOt53/SZPn0u0nP7opH/Cny5VC0F6Zei1fo7rY0/gx5enbynD05TDWcvB+cLZRmIUr
ze+If3H3dyK6UaE3KBrPUTHOvWFFSPY3WYCgibqrjNoNZaH6bDeGd3WNcOqntN7V2lRZgPi+Xmsx
wnW7HirA47cyn4Vs5GcaP3o7aMSp18WF/tKeXCf37qFWlZA2VLJ63DbwflU4SNaUM5QKD0GtDiBZ
vyT2tsXivy2ZjDvnpYW98Q9Vfs3Q5WSAOmfBpyosdnqY8oINmC8HoFPMhIEjB//gbsUlU5xJGa0R
PkQDLsdMbskIxVWWNyPZbwcg63IBUij5tz5DKM6iGAS/a46WANNjs2p6Kwk4+NmQdPkPvCt2tnmA
rK0gdjYQPeEeHNmUoHEfUwxulScSEWXDHORDsHB1jtNWLAJVO4epqDNlWjHhAQbskTPxX1MITuBm
r5kg/TcMfguh8bwRGGxVJ/OjYm0TAHqFREcoOMSeCZw1ujhpZ3hlGCVrAMOsHZLP25FDAOCqfMiF
wyEr646fmNJJoI6MsyenpVazZiDA/fx/YKzmgYxAYpJIJZn7i7tUVYWAhCQQk0UbKEyl3L3IUfPd
MyddQ7Y6tsl4PQWkB7/N9moDfOcRzfbfoZe1LvohsNQyWA67SbDnV26raqjGy5r1PcTEOxp2eSfe
2AP7D2W80QBXs2okd9JSTs5gMcQdLQNTllwK14sCxitw+37bDqyEuLaxvR/k0klojfS8dT6z1Zrj
PwfXAjEMD3THvx3LfOl3+m0x6jA7nOZv4IO/D1JIVt/JP16p0ZH4kIPoct3UPQvtLVvv/4KciXf6
Ekb1Tnxj/+Att+WBoHS0C3MYsovPFwPF4Hl9FcEq3txLKH9ZnKyQx9QHcWP4cUnp2vsKJGlEX/7Y
jWp4G8gm6fEZbdFbpNmUGmveJL6nfKsWMTFR7ot0ml+HZSiX2xsyKAgc4jRsDAMxJ9ktiJNnYEnf
00vQ68vFPfRq+QY6m2mZ+THbM4oJyNe/VUVHjKUHBA9VaJ4YgDVDGiQZ+valHEdLVj0GiY4DZU7A
Is1AYz5yibtgYB8ldr92qNtGgxbMDh0MvwXQDuuGxjFLAOgEfkR5ka8bbHahXea912rYR3p6W7KB
ZVFlLKdocuL5e6Zh4eqEyw7upleTA1S82aO4jVJFIk5RnddJ66wFJcgWKTlSoviavMlVOv0l4zrd
6bNs+Vvscnm5B2fAWHkZUI9venxCLS/427Ab5tnVveIa1yFe3cZhq7NMwev0Ang4mrIZ5oz0Pft4
TxfCwI2EP9WbQX1zLntA5zSgOvpZOIk9GioLWgOJqNFHAnr64soPvyah+7Q6WMJSuE39zhmkcMw1
CMR6AFt1QPeG4d0WdFkAXhVRriS7pnMrkP4zXAJ45ve1EbYj4yaf8kfYkH50PDUt+n6Bt7sIiiib
nBY+wI1lDDNY0jTBH4nLrfQOBgIbyvdfMrlkZpmlWPqgJ2Q3nYo9W3lKb/aOGaTm9O7Nkdr8zc+T
DBIE+1yK1UrbjB+4f12q85t3ckuugEGz62qcU2CG56uVvyMi5/BJmpS0Df8Tfsg8WyuEpBbeztiV
7Eaiz4Gvzujk7y4+tWjl5TCD4lbVYjvouGf5fr1bhqGHac77oICgsIj+uCdAVzTtPmxX4K7WdQYO
C/oREg2/J5Dc4LQtcQRM8SpeIiuZJy2gktk1RC63SNtL2i9vje8tQakF7QnnB53e80BGuh8c6Uut
vOw9/IMGj5rXo/IqR5s/7LxHwQKSnOGx73mcv4qw10nzi7V9wPGsddS7OwtGQ0Fh3uOYgPN1tJhX
VoKcXnU7ut4rkAk8WXC2LMpOlgVi9U7pnHwCS65KAecg045dL9IbZ56ANHgPiYzGpEO9J2Fv+J4u
pmhKTKXhk43W8oRhN8e0J3NOx8GQ9tYfY2HCXSbfGtXv2Tj6Re4NFc2ibk5KB/cIyTbrFVTfCFit
AYebBjk0VAccoW3ZGpDPL6bzDYVOwRcjvLPd8Kqc60Td0hhecUEkkLqUAy3DDQyHBo5yJ5Qkl8Mb
jLLiZLL4O093gx9YCorckDiFcdlL+C7kyxX8735QJwTJwSn1GmF0lDrMII92wIWLir9x/JAar6V6
ZYTfeQfyVgjkznGXaXKYGcCeUqxrro5qwP6Mjm0sG++TArpdNIPzyB9eAEqo8bueh3iOLypLHCBb
gOLxGDbQnMM3VmCTZcAIlrzYnVs6ECQWUgl/msajvAThs3w0w4+KeNqZIK4IYi7QeQYGUfeqGfhe
ZgS77nCepuSaNkAVMOVrXs79ud/2cnd6UvVzmqWkCtJR1po481fL8EroL8GUZ4zHCGerfw6HIsge
/ieZ+/5vi0uLv92DqsLfYtCIbWLkrsyMIEsgRvb5dj3v9cxRWOw/xqskHPg7GNXh2cUY0iEGuFp5
nJWexcXsM4PBOTljUH3pqMuo5iXe8stsn/l8Rcaheu/DAUinq/KXOuI0HwSHg5htcUnFZ7If5Cbd
fCVu7C+tMOJXcILM5NU7kRb3K45M992Ad5lE6486KSGua2KKPQuW4sU+kg2MR38n6xp0GLwbFkkH
gr2fuFr+P2qyqV7H2lOZGQM1MmM80PxzxoJsKKHfyGBLTHLGE9uJkBn6YIPLtDh34wnsY3Jf7vVt
2yA3E5IL2Q+0UoJHjt1Su/63+UD4kzZakiXV9CzgYqehFjMp1ZTT5k8K/lg8O6LgY6UtqV7j3Erx
Zcx7teGdm9D3QMGgJsyAn9Sco7NHVUxm5OhE3F3JKIDZ/fbW1IW+9BkrL6FkdxRp5sBofzYEaxMS
x0Z7QmahlNEiyQRvjwnjKN3UZQf2OC4RPTEpGTJc5VeydK4C+SXbCQPUmOf4Eg1cuJTB2qVcpDsD
/K1APhHC5aN+smPDRw38erZ5o2FSQ8sGXptkE5IZ3x9rJ1hkkSXq7ERfbcwS5GYK6vVcwBfH+Vl5
c3wMXDv9Z1Uh0DZirFRgO+PLVdsRT/NP7GoFfkNi0BAkQ2gcMzCztvgEqjO3WxrtFP0eYNqklhda
AEU02O6pBRD4sDogoOMdzz6RnPNJ8HoNdoaC6W94IA5sHuLsk/FpUmrJTKCNwZxWd2sIywM4knr5
DUbMrrOvhkgwC4EsrcGS3syVNfQ8fjM1LTrH+FRSxLbLgfrDXTD59GEUnSAOptyL8JA+JapUNZPU
24iWYp70okmMYL3lWMZwp5ZsD2HueD0UWEqNkGpNYp9j6S0mcDivILyeBNtRCM9UPK5iAqsllWST
KmrJoevEErRpwz+By0l7mwHnTNJgAm4YmnxHz7hutbzlbgbj0xRHSRoOtq4tyP4P/TqX4iK2MD2j
2ftGOET4MzoH8K16yIuTJ8yycyGhAHPkeLUqx3YOwaLFgVImwcpgchvsFbysAa9eH1VEjY/s+yTO
FCA2P4Aoxp+j8wDgT9+ukt0CeJxB8Ne28R4/jPPO/Uc6G854YJyfJ+UMBQRE6A+EII4JUz8pdt/w
QAkc1zHJQGlRpJeFA2le/MMgJnabk5OTx7vYo2aNhzgOzzX4zBK7rVEhHXSYFFzRvSIsJFfURdpB
FdM1LkZAY/nzwv64ZWPr8SopgQv9UIwPjphced1hmK/NtoLbnbvyqoz+DwMYBmvthiEgZEm6VKSK
j6Ktk1Hp5S8LiVHBrh3Z4qjxzs3DZzzU9hzAEF3navjdc0ONvDbtmKXpRmKMTW4ADJ0GPuEZ2mWd
akWbMmdLkUHPNfIToilTLfINLajOdzR/9rhahiyyDRbORA0/nlEGULbRoU+6dUrMV4K90KnH5Yrr
TjcGZLShpeolJl3Zv76zPuKN+mw6HYt8RF8YWEm4zj89dS/2QMOZioPnapIWeebLb4lp7USxHXka
Y5YvSw3Ex636O9XjmCCNmgH8IQz9mBOyCe0txU1bSbSKsctNMoy4Pm8CmW1RD904+3aac+mg3Yiw
rTNMwm8DvC5/qLf0z1USF2MxOBrvGMxmsxd94lkH+lYIlUwMFhfK4awo1NsAJF91FtvguPsB1jk8
PqHpKVetwqKxc7hsaR7dJQnqxJtJMLZgJL1p4giD8VBs2VGaw/4VfnXI4/ZAGb4OVslaVqp/OqCR
+fU8CRX83rBS2f9x2FMqr+wlYna0pdwjSPUp/7N/7lgdCh7CTiUMandAMN/XC8fhl140YbZIB8Q4
zjGjM0gcUxilBgKRThv4lxdllTLNPmKi/ggbQxK7GwC0BFZQq6nBn+Z0oUdS30SGpzJ/X2vI9jvY
C77VfbMLyZuGuWHPojm5HQHTs7pIpJYlWPcH8TtA1H3ZfCRLyeZ306wryL9y6nm0k51stwDhfnXS
4LbkTpKXVy/8wvwhYIdCO1TwoLiJpxuvVz4WOuyV1iFpED61s2boOk7omILgyECyWUtXfmKGYaRL
hlzLQRh0RfYgc5zn976Mzv07q2kcm+0GqIJD7xesoWBae2aqqbRa3l7vcGnCW7biCqGsZHrRPLK9
XA20LkzkZwv4H/399FxC//prrmmEAifw1DEwEL+VREQF+RS2S/aC5TpIQiq57KeOo4/OhJwArRUw
mzkkW6u1q/PzwUhAAZFPSKm4oLEAunW0hmXGYdeRLNIr9DO7VAUglhLtm1/50JPxfVYzMgclW5tH
L/KNubJM+KxFUtm1/XABOovzyEuyLNElJ513eXUsCf06mjuBJZJnIEyeIBrGrVwChFXJBAfBXkcZ
aUXQJyDFblIsYc/dLDzbLSvTgHF5e3cD71/YuQLv22UmS754p4ks8U+fkB0svx5Umgo/L/eivK2I
/vuI9d/9S1fXSfMvMqSyxMRUtBlG1l1hbJCH6EUk0pUWtmM3uGq8D7vbREZxJEI5yTzZ/QJMOhpX
Yk7vutuWlH3W2rsHPm/wWUPySOPJOtIHrAHEEzlLWp1+Za94R+BXW0r1fm2KqvVlLn2hR5rde7+V
UO4ZQcX2kfkwWTpr74bvRh8kWK4ViTXSgr6KsjhFcMFiVzugXwJLcko43w9H3uonXC5AOD3RaOX8
6DLXNvXDHhghFmr74yJ9lYVwaWoTFuynjv+o5Guon3Qe5PrzZoZ+2UBS8ztJlBSxFdTy5y5s3CW7
dpRrdxcFIygXOiIp1mEYzGFgPA3S8WFuqO8fIGfGZQMF1Qduf4hFm7iTbARg1BSzEo4oqU/mFE/1
hwHzNzeCv/c0pUMpv5S/MUimWzc6CSHaTePCyEm2qlnBLfFglrIOWu8HEAmQCRkPWkb9xk0LZWz0
EtM/qiCk0sxgMFZmFDtGT9/R3G7BFOJQWkjQ379dvgcp+U7HdShzKAm7MPnX5WnE/bgZZEC1brla
uqQ/4dgB5drjHe5gi3fqX0pCu9R2M+LYTLd1hw/x5mfpYx0yUX9dfIW/DyqwC+Q2S3q8PelgebxE
KPHkhd2xbDMrzqVOqwUUIEmoMDtnOiv/9WLI/ELCu4vc8qJql3Y9T4p9n0T8++hGvuYccTXOeLGn
1uvB8vmRKhEYKZ8lSq0LwOA61UU/xNJVrc3D4uXxZE8XaiQvPyBzJW/UcYLmp/gzDaBAKIxrLUF8
HlyWvf/2snfE48TElyojtpJsGNlH3opivXKIcIEftDPJpmBCXYA6qJNdlq+DLPU3jTwCqd75z4UC
c8GJGvlBqGXm/Arl3CyzRxXP6bzzogXnRya6jE+sjWK+Dd0jLfPcUFKuNtX4zM0eMqBemwhIKDfR
qOB3oMDymvnmq7GAudACNtB+XWHYGeb4ZPFr2j5Qt/p7yjy718WauGbmGSYTPQmLD2cAXx0LGchb
lUL5PKMNhAr1Fm9i27M5itYze9+Pgjc/J7pV6e9cvqKJDca+YP23JBwIHzE7u6AwXbfSFIk7pXBT
X8bcusalUrUh3KPO8W5SSI5CtZRcsZU8AsEo+tpUOco1kD3IPJWRJhw3nXDHUHeu9Ia/786lcz1w
yCSUeQ9yCLqAdN1rdEt0kfUWMpKea3UpZnCeObROLvZBJdoI8cS/sboiGCc7pVaw4Ai6gxhdkQVD
NbAi6uel0jpF5hC7ZzXuSDzLWntRVR4TniuhYov3DEtKldQTEu+KGkOYq+odTXO8sAHz1gg8Z3Oi
4BusK+0Ujup5tdRxTdcmqE7mztuUrvHd0pKG9wktxn/3G6+uZbbpu8LKT7BbXq5VkAcPyrSkrw5a
qRMP6sISUyukQ/q2IniGoT49f/JuS8y2O19EU1xKjwSkZS/PWNxXmI+5mzx2L50pCf0+DPi1b32S
KP9V5JOrVqBadDoEt+O8bxe6QaJt/l1KECSXd84X63CosPXFNbrYa1S1s2UzDDA1A1rByfZ6egXQ
j24xc9Llk4N2A/pG43wCeImiiCN8hks8g7tWnHMEN+YW2W+TYFwEDiD+5IP9zBhgusEVO85I4mQm
cZD3UySQ2xuWLJKHolOkouisIncRVjHgwPQyWRm4rGXaVH1Qwf7d3iJ0ik3i3LrmCprLWWqpS+ED
t33K9JzgNLRCtSSMksJ5lpiMJQbVry3DbtEX1YdfOg8Jzyufbg8ONiJdJCVdC6ffl954NWzX3QhH
XgNNs/FSphy/zBsXGhFAyUSVZzsCrmEcnRWrMo+9DOfSLQL3pVXvNzsqA8fQ2FaTrztVzb96/Qra
Kyw8Z2hT8Rx5bLALi3jI3u1yvSu9xYaQTN68if3Iv1DM7csmx5GwmOcjOzt6r3Ib/lIEMzGY3AeG
SKfjG7iCBY756mNNuZXvXb935bhWCggBtjAW8LcKboHIuKTJnTiD1sFQNukkbcM37QBbD6Bo2CRx
jzIFhLQhWeD4wjqFU3HWMuTfm8/LX+r7v2hboR4G2qZewxuHOZ6Vm9a2gs5M74mkFCBjCFWAMPfU
8MxzHGP/PbcpauH7+wtFAzonDs70R3RKikg5x41DWd376cfZyL6fqTk/0hApKAs6hNmJJB6AByXi
mvAKe61zMR8+VSCsuc+8Mhs3GSs2HAbWRfySxlhSET5+cauw58S4fJDiT6nmcvpafttX2t9+crYr
+uBdNTikFycH4AB9uI6aFXqEEjtmJCwWbZC1YCUEeYj8qSsVVxNyVDoC0t0kV10WNwNTRPH7W4PF
RnQEmYvGuIYJ3Ujmpx+MlIWr+2SSMntN+WXjVH1520FK07Jm8l4aM6C7tkHxRmwZjvMWDBG/GTeZ
EZEBw1G1gcNAxtZd51mx+8vJvmpTLinaFRAPu/EUPMA1mheuhwVasY5ZGcPgVpD6BAI2KlmQVkT7
Os6eWOVPuzavR0i/MzIalv7epEJi0lw7pTVviurcJBR50G0H66E0IAdSAKXMYRSsCKyt4D6ah262
48lR4bU2wxIMRJ+1aWUdpJ0jmruDSuOZ1OUXCo8QMBLOEkGg7Go6duVgL9Vy2I+6BNeY+MIwFrqU
gMMUXa21edtXSj0rhRkGd0HpUqkXoWssX1/UH/Ku96vUU+t2enK0Ucf9PemcRvuYS+xATXvWAKsN
ISwV97v3kx+VXzHsu+WrcrYBXMp+q3vx3GWqXyHomKJweTqtimCZRp7e3WDWMnjwDc6ilW82To8v
+TtHyUmuIkCQcJm0MDdvcLSoHLjGU75zud3NlWGkrCIREfiJ9K36D2Fhw0Wqi60ddeCorHyNy+GZ
JRr6BHAUip2jQ/0SdMVWpz5cZ+xNvyO/uEp/krEe0duFdNwhyhqrHaNRy/sE4E1XLHSjaANoA64A
H42346zojTnDme6NxAcQ/6WkkzNRVMTO9fQ+i9GeR4sXszYs5YS/d/ULrC4QwjaHi57+ImJ0svy6
bkzVT+3f7HJLjrd52ScrCPSx8FHqB+tpV52iOokh1QVb3JMaZTokuZLfz28bdVRh1zCF8B67nLLa
sH38gspmfYD2N1dHzLIq+N/iPcwQ6oOFnZ3aqOmTiP5dXzSSd1fZKuXpMea0Cz0FwxYv3WwTJcmA
t7e8EqGxRP4OGoKhTQ7fTdLKU2GI2PSJgAsmMDRRDx40M45/6ftJ8SjvcaZ06sqifj6meyOIoHxF
dshTK6ZoLoJNGkq4DSS6KxPzjtxHuStjOxRV8UMrQlPXNHwu7CZMhZxYdrrvNLaXHStHX+1xX64j
XCBVis7fMJsOMB9Eg67pu3eJHEhDDJeoR/EXyFgi0GyLlQ6JRnrd9I2+brkXLTpaIzgqjHwr8z0b
KBh1W5IU4C0QTRfHuR43yEb60GT9moJYBBZ65wl6j70q2132wdR+2ZM/mUkEzN5ksluUFxyVCR4C
2FqVt5HAtZ4PXvAJz8QHi0mNPZ9nbvQ0H7JvZxx8WMG7AirJMDYVX8e7M9wvbN/NwEfX2YRY4zA4
7YBbRF27vxOK2+Fms01kMazZgCowf4mNchmR8lknEFUKNpOGM4fg87N1UQ8wu2KVxCxxNKWp3lwF
I31u0JvEg3HVkOPjMqAgH0B+RUvNbBB8edV7PizknmZTTypM8X/x7ipjevMuuFc17ZO2KCScYUWi
Xq1kHaGaTd+iL4O+zvuc5H/jREEHhsbPUI/M4iaexrme9GQtkqm6ORImhV0QpdbO6rty2/l/WyK3
ssJpvHEVCWTX8N8qqc5WPShVN+dVHKJsoEip1M2OWwjfxAPwG2ulGL2ySAApuEe4wF87QnY/2qMZ
1QdZX+0zd18dK4sAhr8+CH6KxF1Kh9ZKpoT3ZWLmvDL3CdRPj2owG+Pxn0dPIB6nBa+zCEfPsuaj
2Jr30o8DP6TNPpZy7s6jiLucW4f0d78BcavqAdql+pmo8mdg7H4gG3+kSoOJHbx2bNBbYasMHpnD
8hMiEXew09XWRlzGGWXUqcq+Xwvm5T9uAVtYZi7JAgY9ELSf8mzjxfrTiwbOMNyhRfYdC1kDaayY
E6OAN5MFqqlNRaqO97iSQOFVURWbPtFJLyJnegDX+xt4nzS2wNVcQv7jpsp1sYLbqPuFVECrd+Xb
xDLgOIu4wQmakukWMRJEtSYDqACvZYRNSEjB1lLQVGyV2J7+bhS1mXn+IpJnseK/G75iOFaH1hPM
HItxUJ5b+x1/lGhcJL5zjE0gsu7UXNQ4kKPZFutK6/nQSYItt59a0D+NhaMfgGdZLlFZjBNLGwzb
rTkuifLnx/MrPWc2gi+HjQmBTdpVkUV12vudCmvMx1esvyFfXNFY3RuCCqdtYdlqAYW0gb1NfVgc
0azIURIEefnHz5JUAZHzMtNepdin15/qvnvhpldK3Z07yAYPyhQ+ceCGeJGo8Y/pddIk1M7+V76p
MHgYiKDOhpa+U7RZHTf5W6HmY9GZLREXWaag60hqEdNLRlJSGHSMfSIFqgzvDTY9ph0YCESvGapT
8XeVj6wJbbkuD8mhrfJbLJ+bAoYOJrOxOWmnnoX7MhKj8NMVXRgieSfSn8SFeNVbfeLk7Y1CSahW
cCYbt4fyXzhgVjI8CtASNfKDMGnq4AGutC6ZnwjsI4mKEUnb/PqvbRlBuY/VnnHNmXvv5v2xAPMJ
WtMbnPR88yUjMXFXDsC53mmtBKJcQeWENdC69X02Sl3Yjib7VBKtN6TXsu6xfC4Rc0hsADQHPQTi
UVV8nYEKU/09kYhsdMpQkKyYH0B5ZyE7YVEvXypnj7zT6zrd3bpfcKgbePERzRIjhfi68D2MJE/J
i+zV8VQy4zM2mRHgPlVxCuY6dNrTi2OGcE2GO8ksS1OCHSqdenvmooPXF90Q2P7VChO/eKC48Kvm
KUErqfn3ZaXL/bKI1Mss+pRZTiZhZ6coMlRuArensz4jrByYIcmdJWHGcMbsBzKRk7SLzukXEZsJ
IzSS0+ZpSVuJmbdgzIGN2PsK3iKdLfjYHuFrtphuw4lPEVTwz4sza3JGCmzk/esdCgxnBXOuYadw
hjI13U7PP4cXiBjqbfG5Z8JeiZTrdUz7cAypH1U8ysbrP4s1It64RnqHvMkYHFC1Y45hjLTXGpbn
u9DcNPWZm/44+ItC2FfreqaA81b6hHZGjujgrdlwASW9+73RpFn1bp8vNx21dFQWpatUhTqU2Wq4
0Eiwjw9KDcMYe/TdwKYCAe2acsrLsYn+yFyuOKU+FDEtmPDgwSb2pCAwALSmtK8B0PLD7xaZqJW1
2Xj2cfIB1k6JebFX7Q475Rp0gcSaYByzGFQPBjbRJlpP82xpMPA5Fdp1Mj1KKmRxofO0q5zYWqi9
LQ51X+wnrvvTXF42SzdLk0RTcMQhVtUC25r57n/91hqaCAh6ERoBd/44AP6CosWFyqfZgUVSeqkg
UahER9vrZcau57/5f3Fsv+Ri6/l0WZ46HTBFUVmGTEKzCytz/RXD1QijAlM24mQGqqEz3TAu2pR3
cMb8CQFG7GlOmgvmMy9N0i+L2WkdqWFshW9Z/zHJ2rA9twvD+i0815G9FIoIgFnEbPyaOtG6OkEA
qDYQXrpPfCe+7ti7H8uuEbsZd+ghHZiPG/wR+jD6CAQB1XkiIcmj2kC6ruaUGx4vCDSY0JGY6mDy
TkmmdcYrfjE8wxyCopVdeEiSixmkNl9KC6Pima1jcA4q7YGpbzrycAcIBM0HB5ERsCrgiyWF4vYw
i1E1/sOP+doUHKg3cW/qDE5KLe7vPvY2MkTvvWkOPyEHyg/0GEeQt8zRioQzPyWKy2MRGkS4SDPu
be4xuf10Jz1iRYPkOdpEG+QRDAzpkxAoSWCbVPHqnlbzso68RkYF9OnM1QQyLxg/2mP6ECKBpW0W
GSk4e4wlsEZMsohVF4CIZY4P0LK14BCPEDto5WnGqGplctosQ3jsGfIZegqSXq272P5tNhWfHS63
gdvAgfIioVTXBGfz2hxJY9z4g78pOafymnnJFa+hSNX809o96ATL4hjUU9yjJqkHzEPuc07YqIrq
AMOrEFeCbMwuXrACn+z9zPM8vim0iY1AR5AmSsdddoiOq98HQq5A7EjRGa1jBF85Ze2IHwLELCJg
f7H6g1wWV3qU1Xg15ZaYC82sebHGkoAfEgAQO+pGG4g735+GMLaqzZG+GfAbnLRbVHanb4NWqDV0
vxASis3vTqW+nzqwOc708tFAJkL261smadNVZYRfrqFqTafjN1N0EYY9L9Qu1TZB6yHMPwNunHsH
lonfimxBzHrcjuOPemMZW7HcJO5JS5ercfvbMaKTHEibwp/pXNBi4nqyl1YjSWN/nzKVbn2BQ1es
CNaqT4RY1PjEzEebWM1rN4YtMCFUuFtfD/A4fTFBeSzM1JuzNmCCDi93LJ1Hux1OCElpm20Y4PsO
32PFJsh2WCEJ9GymxlPS2uAA6E9NjEJFbhMiGqG1M0xxwjGgz9hr6Kf+t7DmxpYK+avZheZKrf29
6lTFCRBToRgIPrnuYWZ/OoNnx7heoIls74IBWBp1fNTXX7t0J7HxzvLxJxS+ZYmwgYvWSvxS0cIz
cJNEiph0td7ohEYjcVmzG1CRoEH1y0FS1vuLR7V33xUDjHFplecoHkO/ZKeD4KDWl9MZmF7j0a/8
4DkyIjS9Ptgv5JvpGd7Sx22mFOHr+vq/P2aCi0aSRBQM5XxiBoN3Ro/gAVmzf2V+tqfBHqE3Y4y3
91nLp6KZakIKWKFhfqaL/vd2UstVIqjb+ne4TcHwP9k8OWVof1+KNwuBri1EfliZEW6e3XOf7MA9
kX6gul34DDhHoY0zeyDuVFqkgEX/lEy/nkl6EJrO2satovFnBN3N2z1vDe/2qpXOpeoTfJnU94UO
pECY6m0X8E1qxZ2xdGaUvJ7ahbMLJDHE+SmJlW+gJdubv6vtzEr3S9WbHFxlNRfMZHvxB2fpeSQA
FqP4MbWfjDplY2uU8RTU1stq6aUyg4Pei5sxIK1qaYH4cFAWAXmTQlZoSRRROJAbrr/+ERKB4++s
jmLAKmwkk7aZuhlwJJShoSw6yJWu1XvS+POuhUXxTzOLAcVEGUgxik/jyMYa3T8t9ABSeEywwrNG
8J407w6hOKCjWIFy75FhV9R9bKYlyyCGQn9STDXkv54TsrSsAng89UDMSJ+6o41pjCvpvEqs/reE
rXTuo3LIBCBvKv0WWS7dlZ4r0mYbJyD3vW6kV6cjI0kUv1W+bUrN3ql1L9gBE2MMLwB6mDYyf4Th
gizKkvzaxtn18C/zROJvqiybe3VQVOMrU6OANvRqTqOU7aOQqcs9qGZqazy6JrPcIVkKq2c05Wj6
7X+LmO8qrMOI8V8pR9dQzLuleIlmybJ+2qeUpBAVv5Usf7EOxEGum3C0Q1oDkh5TFQJCoNe2HVNX
RXQPbpXQmNdm1PvTmx+8I6RTlsmU/nuIzbCGBj9jYcjBZuyAzgsm5siHXRYQVTt+h/vJHhUWNjMB
NRHy4Tir2ut/r/Ywp/tSNF6yrdXyYi7DZhzLIe4VuCBznoYyRfNH5/GCQgG8tM9E6w5bNOw7bK+D
xn+AOReJDiGxbzmFNWqr5BLt8VIO+aq8BEUycqPXVtzky24QkHOkHwXFqQcxTUkybWpeFCx/UEWY
Zw3sjhJg82XIrbuwEzKS/2QgWG8vL6ecjvLDN/Z30ve3nBXB4OqYjFYtgV2XGlBDj1JsCplts/N5
OfSy81HPPs8c66QfSsSHIn1P3/Rcry+tlUJV5ePpuy3ZOgg9hs/oqfN79J32RC3ITuk9jZPyDe0a
ZerYPcQ/QxVWRAkUVUc3oJcFkax6t6z8ksv2Alhho0IQVECmKmFlrpKiRXA7g9MQLYSwbJvPj4t5
lNOiYnPOu57msyOoUCLmLt74j4ByocBsKUqz7qlMpbt4VefR1iOya//0WSfV2+F1cm3VZhv9Ux+L
rTkrqTCPk4k/kbpcmcbzhEkGp8jUrKd1P6Fl/JcYKvdrSaa1PytaaBOYf4DQBtcIoGUh4ixAyc6e
sPJPtLHiZTpmnzxHsuUCHrYmzjYgbO2ZdhYA1L3u6BlxwFhcWasq8uuJCFYSELdQmwgxoq16yGEO
lhBAcvDejb/RGNbTUg0PkKrba8FpdrRvMInRINdjc/X45AmPENqD8DdiVHgBMvQxJPVJsG6Llsj3
q1L6NX+diJ8z3DvtNRiEJaYCFelkbxss7Q3ScL5/HIdXKwSYF15MUO1+Q4nBs75RX9Ldq48l108f
XVtgzV1encZGhpFdODsSFpit+wKcp6Bv9dKugCtGm+LaI05iJq8+s08AV53qfTs0t+Z2eSPPwZbT
/kag34ix4w7Oxcktn/+373+kvOIqfcZGefiXS84aLkwwI8/79R9HJRuX+YFZAuztAd8H0YngDNMg
otfLE9UDdb7umw8FchPDx9O0Hhyfny86XD548a9cdxCi93ZYiuUo+DZ5MxwrjtJnGXnXtsvavjW/
uPRNA1Er9SY0CFErqnniDi5f6cX0IhnTDWmzlVgtLna5QlR1K61qdVWPFzPQvLB/hogLCYvC6j+g
KNVVe/mtD6GDLeXPYifv2i//PpAi/YqFXs4mrNK44vp6E/aAPDd3K0U9Qbmz3VbnTlDXW/Stn/pc
tLjoZEXKqVEUPPrp2cPyfjkI/9gNlW/t7lHKUK302YimnyJq6+sxBW9YlWP6S9NQMbhpJyvGNHnq
3+LfK5MnARA73cIWLYr6YeWQEPD45QvKlQV3IQWNrTxIeyYGI3wYaUhyg98RmKP2vUvGkxHnmDr9
ML1MXhcAqFkRGmCO0xzvShFMLZ3sWUp38R/quEavGDEUCqDCCUux3BvDUQ6sQ+AKeGMooH9/pl9N
2DZDr1NppGMV63Rg5uOBBz8XzKPSEKLYFVubIwCHTcnm/9L7x2V8mdW7+z+SBJLJnYdLrCESaqLI
7itFUygEtvjk29H5iNcRHneK2tkuBasBuGLwrnXgQaW7pyv6SBHD1ACUNdvxaDcOWBCMMvT3KsLL
GWUc3/24moEJRIPWF4ru5B9CZEwUWnPVPDm3OxL5ukGU7rl4DJ3/4rcU5DaQh7i5PaHAsliySucN
M4EA1H0PaD03Iqhgj0PES1tN1gSKx0dGJe7ZSiEG82A/SHBZMxpmQNdi+z9TQmn3fe98lJOUpxl/
bw1SDCOhd/ZOPyknEtnPBDGjSuRlaPPXsi8ZdxIWiIodPqpkcoG9ixuWYMQ3829y6UFRYtvbx+gU
TIy83ko3qavP80dSJg8hm8UPMBMaBwhaVqTgiLORRjH2hpvSmyyGtrrlErokd7mRbAxceOOlz0PQ
5k7CJ079A3GLokFhD4lmEsJhmr+FTp8NCV2NhiHKKE0lxvqV9qhIzs+lR3NhGuLME0Ipa9nyzR7n
YWea4ZIy1nUIDr3SwCkV370YvuwXIHUwA6BPOYgjTYNHsuUQb5sgez3r5wPT+aTdvlyK9mmqxLz1
qUVUYHx0286mLv7R1i/39ojQan9kQtzR69pBlTSV0wkBg2HeoH2fd7YruaZl6Wq1t3OjQIMz2SCT
va/lkY3DX+D0zTnav0w9w/O9yINXmhKCJj/bBr27XpAiCFKoxvb5l8PNFZEXpM7iQ7HgX8a0Fa5Q
mN+AlaOtMcKCgmLnXFApTXsKBsqdJeF2FiVzP3e1M+X9ZzXWXdVh4J+NYRJMBQy8wN1h/YvdcKLJ
FlUo3Ko+Xrexn63fKe27KhCvv9oGw6q083s0+BbEqFycjMqpqv/FFmK1zgTcIf1attfH+caG2naj
zzOGOXMVb8EIxlFJNV22tItUtLpCmMB57CrlsQd17jABUs7Lko6NQ+7CyrjTHSu7IMO46uNs0/qq
sCu/mu9A106w+hKnu8mNhVtUX0gediJNvMwNwq88MM7xS28Blp7TvE0+QIusjteMm3lI+UykL5CQ
jgQa1w8jv9drHpwCkysgEdghqnPt24wlVAoKzjXjmmMK6PzwhK3wDmd0ly6gN3ZFStj7/0ANJS9t
EAqoMXUd09Ana1Br+Xjts+gyWFfhlD3yBEL3s9GXSzJ88Swgo8jes8gJu0ennEiY7LlsXmjNyXy/
wkQ0KYnRjoZ49wtY+guEBaECSimY5ik/8YY3gztXDo++q5ynp1s8UfJG1N972lu90jSd4dNcDx7A
Xn18Y+JPdxB59kiAtNTodgy2cOeYyVRvZIE2Aznixb3KA9FFkTE4XpkLC3jd9La96xjecq5Zrf6j
K6Ef3BT3vm8sztZfOYrwCFKvCuJTIfOJjhranUanLZVbid5sQAeZlETww/PKGhEFY/uCxaRA+J3W
REtm11tYEIyvTSsW5VPFu5f49D/Ieauyg3UDArbcEUaNvDOnmr9WNQpSDIZjOHN681v/qQaiXOv/
mCPjJQNSTjQm7jhwK+Sh0vVmyrQTH+Roslig07aGrKL5bhs4qvwU5htzn7YkkRN+hisIx1D/I3eC
bL51H9Q0dk2bt56t4IqhUnuBXZlxhfTd+AWEKMd8v+zhKhgzBX06JqBijd4FQIBhX8IbD1/rwicr
MGZ3ea6PqJi1IPt62SMplx5ElvHdafu/vaVlHFxtFgT5HcWZbJm7IRGV2TNC95G+SkwHur5Dv0OQ
x3/mfaeQ7vqtbDtVsRef4TEi3JsaaoW2gIRi578cZl3viYegdtr7wgyiz6bPTe8beVr/d0V+Oex5
Ck+EgRvDRoEXIMw8KxzvIA1BJeW88/9dF0ENcazP021vB8gwhzAz9DqMgB/WjfwtlofEovLpvH9Z
crzCdxQ7nnKky5Pyzs5vUqAisHUa3881lKmmbCxZPbEqLbkpZUeQY8Wki/QTyz1w7c30It5Hb5Oc
PE8SFRi1AIvPq/+EUH5qgj82gpDqPpGAzJir1dtZv35D8pUlBDWE12i0gGZ9I59hRlXm993yYuvv
JPEfsK7rr9ti5/AeYpY5A0kSpshQkHBvzbhNvnRQe7ku5OyO3zmbOOme1Eek5YgBmnuy8ZX+PpzC
99BIHAfaCTk6LcsIKH/094ey8UghrPobiSZ3FfKE1n5vyX80bD744oGb7VjkSuZNHR6q1VnjcD0q
mZIlyhM05pWp4iYigron2VVXa+WL5Q6UAh46WCtV8vxNrzrEyBNNf+aSQoloESRjd1eSFh04eOzE
+zzVqbp4VQkUnUtgIC+4TKizrGym/hPjEnm26U+yAfn0gk9/KYGmwKS9dCfJHfAs1DJlV+Oh9J3T
0XdKULBtA1Mv4DvzMT+DuF5KGXSvatZXPhMeaX4pmbTyZY3IBVYot3X54v4Yw+kvCZoiiNpzh5mG
NDaLfJGijZgal5CXnDivVQ/gqkifjgVVn47waRm3Cill/EhyYrmgbdKx8qOVD39BVTnqMwuigcFY
kDto+CswDNKhnDXd0BFUJfaYpcIBhVNjIRipSgaerRXRQ1+uSeNrQRTL/CKLheUGHl+H4WfF4JRh
HjY7OAQtJZ5t5n2pU1/Y40hJ24WtIIyxvOQdjIkNRHdCGSuNZmWUmHKRco0qowhHjfX6NEPijAzb
RclLtAgVw0nZgmWhnYf8HMpZaFtjj83P3U6/H+o7zqv29iCznMJh+WVxzSL47dVum83pdqq33Zpg
ZB/PtRaKYYHJfeclyd1sLzRaLSv6QMQjhq1ao6JW1TfbwdcDA+03v0b0nMYv5sBv+khZF6NX34iY
V0mn+YosdjwUUGCQbFTlc3+gFkWkxbIqNX20ed0BVGeqrP0HbKPjl3R3nus90GgZ6sqQNO6TO/dy
yxoTEQTg3d5JwbxglzulSqj6/j4+JVt7LhudW7byjAjIlCTBmgfJqE6v5H4q4ZxC0ZlGWhhsHXzF
jp0dWefTuPAg+WBXLgsTswSRY4AMHFaRwPXJyFi2fLH/CWvVv3nSN/9FRQEMCJjbTOD1ez2q0PA2
tBiA//0jqUrMoQpkH6gFML64r1+4Qe17Xu8EWu/fpJdytiHrcTP9q9k+gyii1aCos40knZ1AI39L
6S2pobeN2QJdARztVSE3kRCJ4RMllw9WmLvBlChcKFX8nBEhvBFp4EbHjxLOT4OqdsMgZ3VCEFcz
Qfvah5XnEvRFfTkOsMM9e17IQ90tKtEYiNrzhtX9SRL/erHy+6pdjP+k5ihYY14uEyBsYJW1LwQx
YTzXMjf4to2lFkwhuhzRT5+gqnZvBOFo+Q4JisTH+lJid1cqEdcCJJAZgFM/Y2Bq7/X4SrXWIYNg
9LfpkgH2pL1RADENzbML8g9ne9QqHWVx38+8+Pwf6m7izOaQaMQZqNJOhpM3hgcoOPIpkR+SvPfK
I6blRmIMDpgCw5HPIpNKvJFXHFXNrJpFuScbSFgRou764LfAqYSlIS1uwKDkgg0VhfAAUdwHGyL9
yhLBdAVF0oGJTpJYV7JRhEonPJvJNUYP/nVYvZ31vXhi8NB6mylmQALRCBngVRKTdMQE8mddoK/P
OL1eF0nRatJJPzdZTurYPv3U/sbHfVjbOj/AhC9hViNYSKW5r6q0+wAkrBfUGH+el62y8036N2oN
/AB20b7I2isdTkrN8aBY0vBSl3JzY5lcLkiCmcH8+4YsW0W2BDrTWPBSNmwCBP4zleFNy5mgE5Cn
7U4O8JpJH6XeLgs//8RbzE0yFGedDpylTqFxVUvKqTN1h3XLNL0zIZq7Q0cXjbGPVrKaUyWkhbJx
0GlVyj+1r4MpG+h1Tugtij4VCfYHZPPQNLigJoUKr4fsRb3G9hZc2pixcnvNLL8YfJmVgR/a3Pi1
gbrNH/mmIlS4LlXWpWqztIF5Nm5sZ+nTZwHeNUz87AYf7qt9lny0nOFG+INpfcRC602vrg52cErZ
FAmREHRMi7QJ8MMcp01M8oCiBvYqC3+tu3YKkZ0qA/VZ/mB7MpOFMxiK7LC8/JggUyyyVCSC8P9e
Bd5xvJSt3ZMyhgGBpZJU7mj1/b96sZ1b21e17uTXtecDy4/zOe6wITtzGzkZ1tYjT30z6LBdkAgN
YVBAgJkU3Zp//Ma1vR+NJrB19QNscV+c58lXaLEQ3gd89P0NqZK7PsM+v8eeDBL4YxxezprCXF0k
xrk2foLm5DL6/1JWZQmxSprtPIrC/4UYtz+oZ8CkadoR3J9ym9eWAB6jiGqhLTS85jJ7eUQs2YNz
Q2um5gwpeiDH3QYBGs8Wa2NbKCaviMQZHvPDmW//Ls/rM3lWzrqn3XTZH5e53ivfEz/rNKVuS2XO
2H1Qtq1voppTW3e/Z7Wg9pyVJZaf+RYqCTs1JXpCtdTpPHr41UihoX8fxEKimRNcrdGS5kJuUMsh
AELO3qbERO34vOpG1y6V652yXs9UoTLk1J3db589IWGyRjR+Ev91j2I6oAJ/PQlxuzBTxGfGjq1W
V4SKanWqgRHj0FX596Z+t+SDcmrJjj8Pe9S2bhZuVepl2er8eiYYZqvncQyHTFZtYKP2ypyZ1ZUw
mhjEWbPn6ndN6gXK53lCgw6gQ5uZXtQk/D18TwxTrtkxciZTfCsz700aG32dccR6OC4+pLPqPUJQ
/mJvwAIWS3QhzUyHJSaYbEk+1DAdM9ACFROaqVHn2lyDftOQIRSyD5ZkvSp4D7fiqScuMrE3fHrF
AV90sthVqrzhgEe3Ni0SzbVOZa5IhpDwexDX4PSUtZrQ8zUorEbDmE9/sECwx3YOKJHvsKNa4R5z
9bNOZ1K/VkfW1NojVT4G+llbswvyh3u47K/7Int0iN617/MB46Frv8VPxzPGEa0o/sUA3/uojdCY
a5a5p2Qh0cvH/Mtip6B8yCJ1UmwU0jW2GujL1Px0UXQZIMuzL6RQ1eyrzfeTZZSxjUgNg/ueRld+
rI8h7TClFVpcVkkRbmg6SELSta4TaOiNBwCZoJecsRNdlVS6D/htZBaAy2GfzHgL2VCtLbar2Gcl
AE4u9+4sIvg8jwqBCZ8pWBRs9jTgYcpInFu1VCnyTMj/2zUJGJ/T/DPLrxO+PdZSniOB/6hCNduy
P30P5XOheiuBq//ZnzVm4c2Zgmmbl38hPUSP4D2Eko2jT7B4U2q44idCtt7hrsdP8eCU8FO9TQUJ
ErbWt4IVmWgxW4uzQKYS8ldhd7jq+pGPxvwCnaWfANxuT46pxBzQm/NBM9gTQxOh2R5lB4gb8n6/
KPLAzCBgAtdLIuLECGlleqnOeNNVz9CqvWolDRhWH2kH4iM0M7G1HKatzAtc7wmvFnx9SnUlZLkS
vtsvD7Bb2thRN6PRkZPs+UHgLm+kA4VRKAw6ITeQQYaVVj/lU1JpPJogWu+HOMiMXWQwZbcnVbIQ
W9qi3ffKBPQsrLOATSYVJTu/LkIh4O3mViMSN51WX36CgA4fpX4kXlYxY6ye2A54x1i31JdSFy+6
B/Sb1DTwC1xLkpHxbHA/sCkEKfNz7nkKgEr9s1y1PuQh3C+uU02RCB9NKVqwRkRq9gc/IRh4lyu0
xcJCvt+o/IV7MDUihcShxjQtN2FVKY/7c+xU466p1esdobo8Re+Ke4uUmublud6pXQpu0o7LUvFd
tyY24jFdSMdKZbTvMIiPOIGnWkLIxCNsfGWVmKjpQ+Ksj+f9B1LQJN4pEVD+vT9zL+e7JGmaVzqE
uTjjn/P7iG2mMu48OJVNUASkFEJ6k28MuiD9EtXZWaiRRkc9vzvRVsw/mKjkVx4mhL6Vq9j54oqR
SfzL0PwlAvMgVptCQ56FIopipzv0MD1Q/GJmONWVVRy4li7/5RiYPTdRSXvqfSGBUhYWvARy6Ds1
WUvsIayjpTq2AeAMK2WAw/22dSumFmgH5RrgEP5Z3lEqqKdWyHVfH9o+Tg8B08W2mv5ftwJ4gkGd
/v8uL7kscczabwz0WEbn2GUVCfQ5bARWcNh4uzHs4Z8OiTdgySJ3BNSqcX1dvxlSdGRbkzW/diQm
MBlvGQxq2PInD4EYdrSuo9NlcgEo6sfFE2NgJVSioiBRkbFqo06urL+ZYYD0JmF6hrgY/rR2KBGg
D9HIXUfIDbMDSCTb8a3u1iMbrL+kLVADhvQbtSNk5o8IsA9rpElPwPJ1c/H0aQn6ZdgT4Vai6gX7
2XBK8AQHHBPvDgZEcNInv6/EodA12ss25kuyqwXUQcKJ+Mcvmd1ogSg9MH7ambXu1aObpGExKFm2
DhhJdkaohy8PkzAqt+NDT0LRtXtbStI047uKfP4/9DgD/2GsCDKK/cX1XHBv4b435S3C3l7qldh9
BQ5xC7BUHVsqnv81TGhe2HzYWhBPVegdsODHO4cRw4zleQrhk+pna/etM8U2ljb9qD7oaTEjWitC
xdexIDLrPX+Liu6plW6eByCEFbG/JAEbejL8JkcowQ+5qVT0m6gAFGDYsa6dtHis4WnsY0lAp7k/
W0TEDEIHd1MJzOKIw6IMIsSAZLe1yJ0skvvulNn9dr1HnJxtPxBOSOGwBOE4zWujNE2oJEPCnZxZ
Ra5AlxBUhCa4Sj9NBdlv6uiKs31dqGimqhwD2VddEfel91Rn7dzn//h1X8HFMffRx4KyD+CbAcyG
BiCF3HfisEqzHZ7/iWRu5Tq37qgCuhRYdwV4JPxN1IpqgoFl/miCg7AO4ruJrYXyIceUAb3O4v8j
Clar2spgzYEKeViZv5LBo5l4WVYWb8ci/aR9gk5DL5BMxJm6z6xEufUsx5V+d3rcg19wcK3Yaqy9
lUMj1gpawSyZDkd2ufHlJZsSA8tlcOxCvX8FbAR1RnZzhagfIwoRflbfjxOkvTNjrK6Gczvjp0SX
RFsyLkugJFQ14YZe3Vq9P0YxzaF+CaCowiMMKlL0b1L5BqEzXGU0+8MxiXuS0vCOL1+5y1fu4vSI
XhYsBzaHyRPj8H1eTUt7TWCjDT2sABwinfyhs6YA45qEsnO7UQKHMihswWcwPwf3Zu0X5J2PfTgj
qBbBP22z/oCEHNoCOueQW4m441AFwSqURKP5Bl4FDLyCuehUzrnGafqc2RFAakRiMyNC0saKOkk7
H8OIzMJy3efcEgwxMuygzRe6Najm23WXpW/TsoAWx2dTAmnuOGSDnTEkEbr33IhzsWf67v7eIajL
MTpIWFfWFp35CCxw0W7nYKPtmFAsKi4h5MXEv2AvcBbJ6iO690ilftldC8M9Mhzlj0NVR9jwihG5
TpWZ8iaC5Q33Tb5HEgeoU77YLj3AsprUWAdIKZ0hyQCVOPHDOWK522PvLFWF+uvsqsJxx9mil5+2
YxUkPsvppWAEVsPH/vlNp/Icb9PSMjwr0VrPL3tU5kevQpKB5v0yaZ6YsbeZfahdB9ymcHnmqUnf
2mf48kwl8NZjjr/t6yIV7R6DIVamsy8jlCkBEXAC1zJNlIZZNvwmX0lFobFpeR9oy0FOnZcSzoeG
LKGJT79pMzKz5Iq5l0uW9ULMSbd0VKmHIX5D0Ga0okQ5AFlTghpja9IN1uAlCJ8KrhD9lsKSmOo2
RQqVrlu7gZAPq96Rs2ksRx9jr40cGSJkkqEEcc1RQ0obtiDsWKE7qpIPS0s2AFN3gowWrv2Kc3Lf
NS4Fs+O2oxuuNgmxrzX4XzM8LHqkW6iCby2clNIapuBlG0SGvE7dYusDc4kZ3HM53//YNC4SqjaH
emsd3kUYFVfw1A4v+UiwbZiL5VhdC9YhDTExwYpnN5Z/AANonvXHbJ8mphthqmI5X70sD1Q7tKSv
fNq0TwOExj7ibHTxYhin3h2151PmyukR48CGvHukZCmDn27c2FqXfAYlVBAxSjgxxJoYEOSR1av/
XdCg18+HB+KRgy3KT//QptW/rqIcB88mXbWRHDp7EZ2R7sIhwi33D1mkOI7/9d8quX3nv08vvA0N
UloKu94Dov1iJq5mdUcqK2cIbkgLWrXY8PvHrluwJ3AxaV+K6SJSGyyJWA9/ZhO4mtGQooDiQhxk
c5MWSOpeoxBVbhL5C8lSb4zyDHdbbJIPQ3W21dEekMdWw+LZhmqR0G4blZaEqZMBJRT3M4fSj19t
UFLnTbAQecfqYDMpzem3tECE814xROVE35mz04pE3HhlZIrFzkU1/ryxdZKnJu31nYj82+lTL1kU
l5DIEvG6OmMFOB05bVAMLBphRc0Yp0kh8C84SWb/6qGERL6fe6eFnnVyVhj/PmWzyr4eC4PvuevY
4ZK4TmnXv1LuZ8JHhZCVGJ/5zNOrgKF9/5R92IY+9DQGoPj6X10DYJHtPY07iu2upGibptUAwgoD
Oi3hVFrCmxKnlQ2iPkNzYwYvLksEq39MzGvSZxl5mxLDpzYANoG7yDCdxTCBT56Jj8TpjU+pxiaJ
CV6YcgWz8WDmqpFhTvepe6VkCkSUh96htw+NuBPkKRqmOtH0Ybsj0T+jGnrl3pstpwOCTXayJGIT
cfj1uwukKiAsRPxw95PVHw+DkqD4S5mF8lqE5pkPvxTY71t/3bSKLo/wVdLMyEKYu6N5zupY17Tx
BvAsp7IdHDnfTiar6fO32RZ8v/1fFhac7239JqiSPmLfzGCFxynTNIpAMDs1Pa0hXgTtmlcIBQsc
SLhMMHfCExf+VnEC17oDxM7iFaIuyfGsondRAlEWOf+jZaErSrfwMhiAIIWUms07Ip3pLoMXajG/
VCeHsB+dpPNfXeoRXLpOuFnWF+3UPCmw1M+0Y/t2yPa3tOeJC4Iu8p0VFIjaepe0QMMhWOSW2Hbm
HwlErWZlr1GNZXLFP4902pTP629xdypu8BfMEBlvqfCu2lQywE31k1XwmPpUaCWJYHdW27N+Fgq8
tn1A7QTRrG/QWQKwRss5jR4aAfpucsU4Ui4eoy5D3c/3u2DBJ0MbHulnllJMAdph3w3mWUQmw4cO
SmS2x+FsY/D/a2woka+pP2SDi0olXcaXTncsChFxE3PTdTsj3Wij9LKw5tJrXHvSHXPZtQ3sl++E
8RjReiMfAET/jocgf4LN43nusU6eyLyh+nLA+qlL6aYj6T42uMQLZdhA54Jqj5kxLuhWYznpd+Ri
ShEmNhNWNZPjWy+Y3p5P6BlshLMGCiVby1DZwW+QP24Nix23hjLvhJailgGWaN400aLj5spM4lJw
pS4kUxQKn2lPTu3HcCdiS3J0bQx54m8M/p/IbXWgWEOmT6HxuKbLZ8MBM0tKO3fTl3lv4I8jfWf0
QbrpcH3fJl+g2DbTS/yKwt8DtFsvvqLsUORg5ucvLP0iijNJxhKei0Z8gP/yY5fK8mJyg/KLHGte
6KvkUgGywk0ZBTj8YRcIdjVOBxjQW3a+enM3MMELQaxUmXQgrQZ4QCVT8QcsioRCnj7G7mLHVSip
Q129tmEgg+SyHZ0Ni+DX2hHLbWX55R4ymKszvk4/DR5QbsDx7BYJB/tS3uyiOrcFXeRywrJre6AX
fxt3OfhWpjaXJdF0Nx4zPlUUSCW79Eo5J9Jx05NZQGQxeCvl71IgGX2ntD263QOiLH8ygBIJj+wj
9uk9oWLHn5d2NO5FJ8Apntev6fsek5cwVBpfXgxmJQPKy57gBEr0GJG1Q6YqUhg3ZTFn1ZDF3j//
GZrPyPM5ZJ3dxVKuNJh11/aIoHME+q/5/WE4p58WWEkZwzgXGZyvfBLQXje0yWIZKdfYjmnKkIH3
WTldE2mghG2cDhWTR3fsKssouDEmp+lCeU4YElHpmeAgFgkyJi81KndGCRPQ+bhzCV2FxgRtLUrU
ZJdHfGqePZJ/ZJ8hFiAJxMCxDtvvEO8UPoH4gIc6fjqjrhF6WKTqf6AR/R6TU1XSfeBP5WN0SzBu
CD3PTYxEbuXM7D+MjKU1RuZvrLl8cSLTP2GqZp/7V0+BOYCVeUKbv6/avdLyCWMF58Kpp9Fd17q4
xJT7ty85j0ufnrtUeg/KGM6mAhBna8LJKtRodHHHkcuglygVhL5pFGDMfF7kYA5Idly+aspozP76
CVUWWJsYFw8m5qHTtqKjrrisnxIExjiEU2wWtuumgjQ350VSncC6zIZ2f6c+ZhM6NRNDvvkxF+b4
HNHeTGcuhoYUGD+my01KMhvAjo+7wriAJ7zdI2TZHFw/2vTqt3x2bzPTu9gfxBg71LL3UkoOjMLl
axs9OLYvAy7yVgdyTDNw/ISVS0EkQeSb7jpxr0dqUr1YfmsHsGajuCWapfsPhhFjsbgy6fWa/LyM
jxRuVzEFY+ZWZWjPpwr/urT75syHiyXMbn9XBYiCTS9eYAzkcb5ZApCZGqr/sr8BnflQ3bgoKVpa
I4Brx0Uk6EaFu7c6ayw3v+U1xywD61Nz7nKqkz1214yjhSNh6Yl7wLsshY3L5oypCjehjeF9wCvl
B13HRMTh7Vr1wIzShxXR8PpKsF7r6MdgqddQuSo5meslZ//rqLWxEOmdhr5cpAVMzul1zp29mtpK
S7CWxpQhamoIvj1IcpBd36ZiNlQBbX6Kev5GCJKhMbDsShWXxJXLsObG61CuPy7oYpPpWY38uVZn
r4aEKmumrlabtc+88nkAaLGVuY7R8Butrzj+NFK4o3M81c/2RamNB4+IudVp6OqDHiauXuGKJRjY
tkulftAXLZ3+rI9XZtbp6upQWV3K6F+AfrNfFcQenA6YxUaG11h5ubSyFjMhRZbnxMLcUEOqSyun
E9SvGPwVva+dSU9LwgMsiZ9LY79xptTYCFW96ztxhh3xNv/sOmpnQX1agxKK3iHXX3X+meDy7jGM
/SdHSiwSTUsP6e/Lf5Xg/wYr5JD66Ka9WQ5RolG7r6zXFcCyFviav4I47zcsw5HuoMHK1G7hKzO7
GAEnsSTVfMqZXqLjtKwy91CiCMb7au4ZzNXT0szxEk+UJrIMRcv3qnYYVDyqBx1lgxy7Z8B67xDA
jCk21m6/GmT52X3p9zACLvXnoP0M+mRVmpE9CGeag0Y4Exexw9YUTzCM0wXBg9Fi91ernbB1XXfY
JyOqLyY0QW8mp4Ezsndy1OgJ0yWsi16A2dBr0ShZx9T53DuH2cEQoTYCfXTC4H6SmwXZhafLJKom
RGuOYi7HzePs4OO9ZB4dVaEGDkHxMFyAUngtSw24q1naNceZv1O3jB3eiwkeZSTaGuKwANAV6Zre
j0oBuR1IBHebwlezfXaFacAJjAyJwrsyGU8d/DvMrJZYe+4ZHHj4EZPp5iTYSVWzmi7R1o+j7kBO
MFZrUz7gUuo3WZyEatrGvkcaBHy7/5kMAaNVoEUigSlmADOH1VPyv5eDgGu/854XjfxBRHTM+yH8
Ui2cEbq3nx+a1IINHbmueHiBOzEWrsnUIpQ0+9whPbOX0JvtzJTh0NR1Cn86DORhdJHDG7+HuRry
UeUrHyzMCWPEGo/Ax7XpxA2qKq9nTbw5n3mrxMm0N9O23ci3CGnachAkVSEW6k+TaQYpM8SE1mwC
9/A3dY8ezFf3uH+tZ29WS29IgNL9g07+NLSOmy/8t8rlDlxVT5gVatlE0X+cYQ+VzbVd91G/8gQ3
t5uUXi3IzY44pMsBSrPpH70OS8EchZptwABCq9zCugvaazr7SamdXCFoMP4qRaPK9Wz4rU9pONn/
tIZM6VfmGbIvkbPk6vrdfcurSuOqoo9PScViHm0mMWnl2J+ws04/pUN//0RBU2BqeHK1hhVJYeur
yZlg/urqXybW6E5T78cJghBgL6SYynSb1RDTmayFVuxNRFU59qmZePPLGlTssuBdolqJX9GHtenZ
sMo1HCnP6b7FtXb0YcWyULHZ/ZmYZGB/CaQ5OBi3g7SOwS3fUsH1SO++JteAB/HPwe65kwocDoJr
an+JT57XmSAkCdr3Ukn6FuWhfC6NNk0aoiICNiWW4k9R1j2bU857ocXRcZNRm/6XJWbhNTmHSCU3
XoykVkeMuulQwSg41JmOHhfCZ0nbH8v+hkuHx6eIYP/9UXsuMuZgGwBd5TsT5n+OjESRzAYpTmwm
kteQaq8LnLNFobm4BlY6U8/89Ir4+IX+DNucdkeMOPiyiTOgzNXRMevV4xsL30NKjUl3RsrSDWKr
pswDLNfpEF+H3SmVik5rLayCEkHvenGKhqT72uGk4Lh+M9Q4DwuGotQM3vL3szsJ8s6qNXWv6v2t
pjP5qXT+FVq38+1pyV9zAzS+lMFcdQ0lulqycVdj28QX2buff/VIRnmHooPmzOJo/AIFGGvntQDu
5fReCN5Yszho5ZVJnU9g6Yy/qfd/nvosuHfAZDt+JPqCsGoEaCKZ03xSVZhnLwxD4v7fIYn4ABEo
x2PQbMKDesbyU8KO72v0N9R3VYBTibDPFtNXp8jMtgy/mmy/S1n9WzbLKkZ4K6UAi2Ti6lNU9ALb
Cqudk/EULvOq26ofm5ATowrdxZ7qgvY6IFTj1jjV8h4ruK7gM4r8lNDpg1VEsxnPuwEnHV2qbz/o
7AkOv5Fn+HhdrAlhFCqxKF9ydXODBZ4t1HOpWPLtQSTz8SjrwxNq8pVL4BYLJhN2BcKTCA/oQ2wq
6Hp7R4zQru05bGFeLc9L58RdilTt6RxhWruSiWS3xc+wgt9t1uMXVYAOw7SO1l6oMYZuKeSxOhAL
CCWby2a7h2rJpymbvXB49eadiLFwi9BPvzhM4odHeaZmyi4lgD+kfazwVghE5nBuKpsZe1ElCB0d
X9RCnA8ut2mlB+dsAV44b+0mmcOwYUiOkKd0T7h80hdS/XvqWFDJvFtGzKZDk04YVNCBO2YiNGUP
PD7A0F4/A2G6mDnq/VPhXTUAFwAgAMK9b4+V3zrn0qBpm4Kyszrn1X2Zci5/l5VobeSOX7mF/PG8
vjiQ034oXBKy+74SNIkD4hB2nIoAfg2C3LTVEYeD7/usRxBDRRBdapkVl2E5K35Aen1kruvJjy6A
zneh3Apts53CrQ7gJO2mVtMJpvSMuUboVdoQNblYUtj/oMW3BeMCx//QinVxq2YrKLNkZ1TcK8Fi
w9KU2Tshj32dNh3LKIC06JyWvc3RPxqyLqejU+gUGodVDqnyHApK/oXCE8l349sDQYxOaoTV7GR6
hZwylEmF8Fsm9vDdd/w1NPpUJ4N5ET7Trls+j7ZXJ25mcFUqQzoKXBGIXTgmLzPa+fr9KJzIp9OA
fG3H9ARDfqMY2EzLdF7mKFK4T9xkB1qa14spNOajsqxpx7IT5ayNHfzwEYr0qk92cVY/bTMcNTGj
ulsNeMHyXuIYzc3rWqJF/gLE2A8tRmmfgZwFSRzWEE2PpdWl0OLO1KCiKHj2oi03qm78NlulULAJ
zkDIsINDNwQ4010SmB7n6508Cuhh9iC+acjCSmDCK2wPhNRrWvtEKyjY03PfEQ7cEsnE9jMOEfoj
mDo5eh2Nvz/j+FOyQG8IhOAvDq4bVG4Bo+u8GshqRJcTENcyF7F6vmF0qIJRRleVz01Q2eVsylje
TVzubD2zGehbBIyvXPbcpvM4vNm7Pv2e0os1ykcZfh7N4zC4ldNnbH/8UaN9yWUWAFsQTuLmJ+Cf
Pol6zzgPrZ9SJVYRwPVxtmKwQDYadgoSQ0iRHNKsIkcbAeRIMwT7xOb4QZM8j7IWKkswkxBh+Ap2
DAa/YxEIP2OOJuzkvVaZ0gk/LDukJZUKEZk95dPNkjw5KWh0BWTM3wqADiybGjYlQTt2XxOUwsU/
qVzdOV18C2wKW7I5VqZc5lf6amlb6iomN7pvsrwkq9c8PlizmJBqUpkTstVsGQJhibfaDxFgw6yd
I13geHlYrKmew+uKkxe6c9SpPFQT2J01qN5ug6svDHf4aJkNZs7B5Ga+KSdhSdQZ0y7xIcrJ7HLr
h7hTZRoQ8H4KG5LWpltOZ0FRCaftETkSnnDFm9p4wEYWIMNyYoJafPT9+mxEyMhPFfbncsnhHBPf
Cdq3d4So6/3+VYUb92OAa5rCV9BuBUUE1cvsxLn7Fr8VOIcY5LGDKDS2zPoV37zJE1RKWNqEZqk9
O9mZpQ70ivtTBtPsHZtGEPJxBE+LQaOrTWzyBqIj3ZQfgrADn4SLsE/hNfnkIz5TkmGEdt23T6GU
LqBPf8NE29TiO7/FNA8rue+N2Ac39mPHennWeh35QyiibH3ZHH0dsJ99JBgNuf4KZnJFCY8wB+y1
3QyEzcc080XPU9cGlAsXRCmr5I7kW8lZmXzO+bmowMqyUyLjJsirV2jqPeWgqr2Qk4ueIeB9j/5m
y+G2EXxU5Uh6D4GekVw8LXB6AFpPcqFX6nldPsJmVi5cXdO2LmDhXU73LTppjAcheknjFC7Zckor
QplvaTif2dsT5OazouQReGqlmopRXoZGJucimcjjniZJtpcxFdjj32LMvFWo6F9pYBFfq/FBZvpJ
NvZxAmlm9NmtO9d6gHqTeyyAKePWRdkreScBF+FnCeg6v27q76s5Utjkk+oHCKb+Zhq2bEUL+MdI
lOFZaeV6aPklhXWMLNTTR3fjOaMqfCgbuUC6uBen0SoIfkGmF2bIuC9ItJO3rcUrZNseHWyI+7dL
Keo0jinIgkXb075JRANCRvFD6tv30Uzb8l34ZJsMkh54kTk9U4oyBHqBTZ1+TeAtQnYW18+5k+Nh
Ti6iCIAOucnyUMmzcnlBiXi3bgITuh0vhQ/JsukUiVS7fdFSYJxIobbIA7LpFNyHcJQSEQ6SAzoB
LG590xRGmWeu607ojw+2euJ9NPI15bMNuyHNep2JGvt5t+blacKx6Nb/Nu/uXOJUYYNOYMwv3SkE
jWlWS1qnbFft78mQHxVm2Ajqt/ALvM6cR8diE1f0p0TGDiB6/TAf52joR8fePJzFlHBJPwvKf4B8
Qqs2q7IDOVW6v2AeBo4x0Cg9duqgQ6ATF8EDeLloTNYbYyMJTallJMK/uBYlGrAI5E91uBFO4/T+
jy8tvYm2xJvjlAxsOFj+9bzU/ezDW74i56cTSpJwhlKm8L00LldYWh1oZ0Pna/I94Ian7p+aU00s
bLySpDyiupvRw9zdeYkL4U8OXGjoNB0zFdYJLYGp4b68g0TSFGlCAwnhFx6x9vEiG7OBmvOCCzL9
Kvkr+9YHcPuYTbUnkKON9Su8NXDyfl610QdjCldplG2lPmT/tyyIGLGAKWIWlWWiJfi1cr+EKQWv
h59yTVkxBZJ+CmqzrXEmdNUSXUW681S1LPMuU34/l7QwrDlCPwJMMVaD4E2ZwOOxZSAizdNDUl0g
aCrruhNI15Pc3tV2rSUaWqJZZjUtK8KVw98JqKNQj87CoovdB4T/CAjq+GZ8XwQ++ukNpez6PUem
9z5nGyDEQO5gmQfQEGeT2H+kn/cw/35HYLHBlpPrW9+WDtHCw5gsiXe/FIsKyChaZTN/hChZl2aC
vrlvYXJH4dc3DJ6fZK2yd6jk3m7b+OsBAyK6eWgzrMtH6l33RwStoMgZiKAUNiP0+IQ2DgwqfYsY
K5MWP8+E9xUif4jm5n1EsgTYPJW6DTaTx6gzre892FpauPK/CsHcesEYge0ntiSsGSDCbRdYrn4h
bw6D9ohnG9HW94FKE7d96hiomkMeZL7tjAzvYxv5oLRJDiu5kNfmH0ffpiYNUgtMrOLcNOqhfWnM
LEthZPIA2MVnW6/7ypdk+Loj1aGvqeX6JRpE5ElSHNj8bDajsspkKJU2+4OTKo6/ytSKB+9iO7Uv
RH1lz3qF3RFXPIOtO2Bd+Wf/JeLP8uWmCQSpKfbssWOFgAXLs4TjOICGyyWp4Q6pdOV4fnS2DFQb
ITfPQRhB40oLKJ5VdN52DbGxMrOxvLavHYvaNiC6xCSp0fSGOWDJPE4qULvKnpw7o2PMxnSE/WtL
9GjjxLfogD6aBaRdGLq4mE45FZHf4R1HQmkJ7/FiKh53Ups166XWGE/fZwifo5ioV8RjBhu+/wm8
26L25CVkzzw9+k/BKA9KKivEXsIS5D6G3Yl1oqpvwjzMwQB74OSMALan4TTujsAqixEbL/AOOyne
yBsQ6sBbYP6ruRBZXtMKAGQWckh5Bs3izcqK54u9OYpl8XIOjYCxbdt4GuXQ1nlTw2MxkMrfDuic
dj8VcqgQa5LHmlatQqkVye99l/vCe8EUO47ZuZ6P6Fa/RFhKeZqbX7zdFkAoyOX857X0lHr3KX4S
6jQtRZFSBxiirP8BwQxs5oz//xLng876Js9s48HaMvO4pFWwvq8RThnZmYEFqeU1OHaODQsBA+KO
vSUKk94EKMePJwl6DLbL2xjsQ/dGefM7v2UvSFdCieOoK/V+eW/xT1ldBiskELTiCb/kVJ7R6eGt
e8TMv7cwivtuA4GVbJl1gMDJbVGEfZdo9f9aVUXqsCqVCTh32SUuXYW01VEJythCQqbiz3ogkdvA
Xdv5oN21TDgDaqi1x0Sm0Yms255UhbLudIvUbbjKJcEWz1uPrW+1Lvb/pp1EO4vaBhrwE1kzNWny
8Kv0ZidGIJQIgzdJT0U2TvYPK16U1a5Pt63/sT4MoYc8+u2ZqMmhAS+/ninVuMTdVWLSiD6CcNLj
J0hhRDp1OuJI28XgvnmAT2qn+A5+bbfhlwD03Jon7L3NBK0yC2KbN39ngE1jTC5KtbKEYVNLSJtG
+2A3RT1uKWomGmA/ZkNwhr7s084F9qPagK0/OeZleuX65XqqSmgumQa+jtqh4z75e3Dncc29v9tl
ZcucopF5df+UFy7wD/J1TQdA8oVxPJZZ/fBqJ61bsdAFOhkBUWQkCz6LkJgQ5i0AHVcMQC9b6tOY
gERgDk33G3asDl6ogQLlVd7bcTJx84i1b6ndWTwwrxR/DgNw+wMv88Lu/Wwg/WN9OMRY+UcVNIq4
nMfbi0wZ2Qo1w8OgBlqviVjrC6/iytHEtxFIBrkzakJpPFI2uHrlk6pKz4dwomo/+fgwU65j0Gl5
e7jKjBBeRzCHJSd5n4YD+KW23vJhSUIqSIIWxEP9xZYHnXqcboaH3OnHck6Qp3TnEnRB9S29sKjf
y0UJCKgaiqdBN7cc/TzK+G+y8YWXh2O1bVWImqY1oZCZguV0A88hESsOc4ZKFQWNg/Ys82Rvj3tO
i8S39gXOrik679vW5LJb+F2/RKEJ4GOpTH5+fBdzojArH0qBD8kvtGD6EeYjqe9Oxl/pv1/e0e3u
MmU+Kef0dRqK5Xe7wpEXHcgWPeW1HipdpMqn0oV7Okfc1YslCel1ea572FHadigiPKWpKgeA5sLu
MWjVkeJmDl5xEaBKMhLvYIkJ4csFPBGBxvenlbZ3zulAymnxU3mYP0gl1ukeagVjTRUtDuHSpTjO
tvchGITlE1ivMlNRIreQvaWQQHks0EL1aePgDm/8nxgcUkp5DcKmVYKP8ZDRklliafW9ykg5t7vW
SkDS2ZilnhOOpg4DtlzCYETZZXGsG8UM0Pn19omH9ghhW9lCgJpVUyRovcZLxLEbpzWb1cdG12S6
CNs4Lwoy0nDgbDtghu6l3pCIooHn0T2XT6JdL4eJP3cL91oldDYFp4TB2UAzA9ctlXahkh/jCxUi
tYGzbZhUdO0VRl46ditYRldokQ6upxsROyDHWK8x0SGuuVKZAMwB/BTPS9KjVRhkdGZMK5HwmW+B
L5F8KZYAXywB+0mSximPjmsoX8yGE/xP3w7MWVP/wY6EsY6CqOLNHSql6aNwJTn2kuYv+uV5GUYA
2ekBL6brQvE404lDsElYp+TcZFUvb0Qhan/CvtVhP6/S6KSx55UP0jhGgI0b9iVDY4lzdqR8upus
jQsJ5+nyNxOo481QDg/wlRacFzW/cdDzMc2fX25EiMSzg116/3DL4DHFrTxtn9Y1571IN6hrFZwK
Y4coPLAN04ozsJjTgq0MFvJ2G3cq7DsYDlYMj8KzOvItAsFh3OV0XYj/mUpYvkpsoxhze43262of
QR3hExSN1+1f3A73NajH8p7qg/w+kc+WCgtQH/jWAXKw6grRzfDr6adPukIzez2ZddzZKHPG5cxx
usoVuzJBy/PAmbDu/7V3r+cmyDC0R/Z+DYX81iZZZ+6hTVol8PSwAUbvZgBN6CPH77U11IBDY51b
/yualeuennfgiBfs9wD9frlxWuMEMY6GgHTiTAeOx5VI92d6yrn2VqeVwb3ufCqN8qL/gKOGaC0K
lURyfukRdczuPzKbQQku0rmY3urLq0mOCVGyjS87bDY6vaUy/2nges2iyWXlKLOAJq1y7gOaUz0O
i8MXw8LciIX5LH6iscZq9OykQ7Jxct5Ky0/Z3ao1rE2K8RnYHmvBRKeLauh5pgLuAZqJZ3tadKWa
1DQyOx13w97qaimFjKJEHjta2zrxtiRAItIL4f60r8yEugxUGEAo7gTthtbSi3nns5ul29rXyMmE
lhTGnHDyV+ErrMy0I0cWhrnkUwTDQVXrFwShtGkg95jPzdRHNE7+OeLP697UFrvpeEtVMJVfoOXs
Hpc8c3qFa2pcbK13HbpCOdIhMyojf5jNsQpp+f2ZMBmAiwT/bZc8vTdRgrI0+j62cK+TmsGQ5tbj
wrHMt3HdCiqH50zVy7a7CKaT4AZmhlmzYr7folxs8lKCYpe2ZbwNY67lwkLnn2R/q1YgUkbKOBLb
l6Q7qEItDgHw/TUI4puUv9fQlKrUl47Jyh4Gd99CTKXYa0jY75oupTobYt4gjaAUmVRUtdu4MdI8
AKhV/SttUVcv4Ka8/cDwo4EPdE/g5cLArCzpIUdsh+xtJLuz3MfwzoRjp0l9Rvmy0MPZrLx3PnQf
mlBMMmyJsUiAWY38p3HruBhyZBj8hZ8j/tSkvFWJa0b9OFZZEeZ4HfSMm/8R8+/JodlR6wRU4OwO
XuHQax+JTClH+iSRsq65YxVWXDaGkbND8KmrmH6eZugp9QJT42mDvN9Wh9WNIWzqbJvlgkC+obYN
j907pa+elGLTvdTcPrT1fclC7wlIcE1uDVLn2jRgMQvKRMO19/5ejnoCb974SeA0MCGJGOeL7OtX
13LYCCIJV46KKzDczpHlZkyk5RX8p9qTGV6E6E5GYF/T0sztuXMgk0sC3rvUBvMpAZWB4I/djjAf
MIJOuG6uSJn1j9lBGdiKCxfSah2flJhduGN9k0FTXHiNDhrVF+wQSvit60BCHj5+DOBCTYcK8TWv
ptKUWjKOXieUAD7zFGuv1TevfF8leZEXR8eSeCjtmwOTXidz9ltNfvDWocF3Yzmdt0ljEsY4nAEZ
UX44QiMmQRP+7DXC/lUoyRwQ+vkE9ZwqRrCorAg6p1C9HiTqCGJNC2KWQkNqZtvuOSsEZW9gGbhF
64wCyq2uqFxaupGbLN6zQmvy35hkose6XR++mkxT8lU6bzcLIDxKIkCtFIJ9tg66+HEzYDoK5rVW
NxTAi8YUVUgpxvdPEvq7U7ovHr5ZT7CyGAo+BJshfRCyk5dtlfmkFz4YNWJGyqrQ3G2P7SS76ZCg
M1dq7RSm5AGl+DlTyyOVhgbvGwRh4ubj40vQ4u8QInAEzDrciWLOUKvARfq/2XKj7JH31bRrOQn+
5PYobBhd92utzqDwS4DcUy9sLdbwo+BxdKVIv/8AKL63weIh3BU1G1v3ljqCyTIha+OAQrhljGgG
Ic89tFc1tcFQ8oO0HCtbO4+x8+MIQRx7V2MrI8o0IyGCz2cot9UR9JroR+/O2XPsby5lWn6qJsjM
or0c7S86ZrdrzMX+5BKuihANfdB4ytJTZuXa7EznOgNjBKE6vMwq/YfxIe62ZzHC173buPZSpgr+
kTM3VL4ea0YRYM5vjl2ZQaNtIVvXrJ5rUvX/JEH2Ls3yqjftD2+XKk8pneo7kLmP6j4foutFFR8O
YwS2RKFWkYY8qCKf8XA7sx1zEr17F9sxXNpnKJiPsNGj1RbNPI1ANfAprCpMDXW4uVfexoEMutlp
PE5nHAmRxOhW+lQF23KF7JatfwXFBrRhmmoUQ+/wYpu+rdGe0iuBUsVzeeUsNkg+9sBw0/nxktgH
vvw83qxMien30ORzfkJjKwE9kFIyuVBo5SX1nT8W9tD1F7voXTmnmhIUeWhVEY4XNJ349RihOsGA
y89JiNUe7DD6UyEK0T6aXX4/kMM1zwCA+3z4hnxcEd0zmZwkv/L7VmCfoPMtkfNG1g5D2BGjBsyP
5VoOp9xr/B+yYUUnhd0lF+ipPIFoufepS9gvEPF4bwg61WH0CNN73Orf8ZuiEpp/uCHE5BM8/aiL
QPYuvTv6QmcIrxyS0skyTq+NKE5XOsXEHIsHbinZFjcONtkFTZENXukjga+taD39pb5vShFMjJZ3
+Dg23pt/rpn/sZY8DDfBFm09lkjpUH4AZEfmqsOE2gT2FjSZZibXTyukvylfwvIlzpkOcPp57syK
vWfrGUptG0fkHxMBA+Kh+FrI5b+Tv5t26zae7NNvLcAe+yOBd1kin/2bxw5qYdgvXq+ZjvUvdGi1
alGmVOX+OdouD3UeVuGT3+wzpz423iBfcFDAEyN9T9qPWp0eAMBnqNGbQl8nVUpme3CYWQ4OPi7g
cYT1giL43slFUYxeqdreN2/PBrcRZGa13km4VAsEV+/Fb+9wDKVT6CVV/H2oJNjggmkqgaXJSj01
VTaEPmTiDQimxGO5hP2/b9haafwNX4pVaXFmecYyN/JbgKNujl2Oac2dJdAjlwNgxDzPHyCyx8yO
Ow8XNUrmKVpmxRrHFOceYH3OKNOFTKnkXECTUnfILlfzY93coRdLvmgaxwokUgkodRELB8fZqzDo
6hJ9/Y3hNaQ2cjKBgitMuHvpDyvOXF9L6v6tFV8UadM6eFK6GSpVSjV/h1Kn/eHW/tEqpgJFKdjV
pGZCkkSgkBjLj5fyBIIOa/xJp/9L0cltkaO/Lhp4eJRk9xuuiflvEq7otGX2a5V8wOmbpMwZsE9z
YDgnxWu1IQQ6eEX5jhsEweA777ygqW6eirVE4HdpxEdhHDcdRhnfjS+LLK6ZJhyeR8NFkVCqZ2t3
fU/IAeEStWZjEnsjxToQKFr3EBgN96D+QftRVP6hvVdAz/6Yyu2Z0oiN1gIkOEIDR0tpy8sbCKTz
TCBaQUJ9EWvTNRl54yeyOdiZjHCYsk7uSHgN61eDRHf0YwXKmK+FqWEsyV68CKJo2joG9d5OsnqA
NPiQPDEATznIeMWqP9hCTMvwVhho/Xx9K10JTRY/2AW8DAsBTJ/OcK6JDhTVUKkgjB6pRHpVL6ju
wmcOgp7lo2lyFAqvWAP3JLO77GgSsg7CTdLRzorUPk5PuxSGdeefXuQhU8gHVf3qSDlxnzb4iTOb
/nPrCiGbYBoJzsuuCjSjvhIQHl4JwZwqtt3859pDmUY3Hmp1yHqS6MWAODf/3S+NPiYnZ73uJmzo
XnEvkaIMfZXsA1QWSkwQPu1liVmxOxkD96I0A2P7aOdKiBxU9tUSU6MGcHunPC+7hRPXogZd0/pF
KJlmuyPJMX0vTMFhhzCO/OALpUP9wT0/NMfQA8lk9pPpjN+RWPTulT79NKJcw5JRQ7D+VAQjIYa9
McQ7jyIncMOzbQzGjkd2UxL8iyADPqCDmfi1XlLIYbcShGD8VuRbSa8fgbwhjdi8TT0iWQoBQmPT
KGoAR4t0xK39szsl8fTkBh7h9O8zsR4bX4hPqZdms7b67e5kS+oxoS9dIQ6NkevC5GHvAti8cEq4
gMjneg2EF7d9Dj22XJOuQt8nfWpTIAyfGQllGkg5vhAWBkUu6s63cKdck6CoZIvi9W6Y+TeP1pki
qlu5CvVRewYmxByUyVFHNCmerMsjGteJvjSEWfGVEXt1vHevQxRBcF2qb3i95chA+gCugqSXkAhG
sMi+DCKr6DaLUyzdyF7eZBPuh7a1ROkeZQTO18k0GX9Cy5AzULzrPg6EJgBfX8xQExL3E0Akmopy
VUM5xYolTnCBz9MEiOTcPJG9ez7S2IbQQIwr4Cz2aRbPpN9mehbIfJo0bOTHUKg9B65MWay1ew30
6y4mA9azYlLsVBkL+2KUoMc/CX5IXzVMk6DUQlEQ3ey+9ehPL3YseXWgtP4lYhrfqGvGMcxzoUIc
t0SmgvicQ3Js7prgg6yepBHiy83iQCUHqDPYvYCOeKobXxMu3hs3mg5X46UXS3PaQlSvaMveuJkO
aKMJZXGVkgOGOVaFQ+rWLGptUdWi0eTvnUE3W80ErqWrnZCUpMEKeP0FvhnJKOuySJQ2XgfMk0cf
nGm7cX+Tyw9K4b8kxZQF6v1OzfdpGEK+KNPjoTJqXnsGS11V9h6CLEg1Ud/mxLux6Xi6n1JHokF5
W5BE2TO/ZQeraAV0O/itM7D7YHZpQOBB9zVIWuIpCFVbcAs3XuvwYcmEeqq8dFVEThBwVEYWuaSO
m6kePaLjbx3Hc6La1TIcQAMmQsUDJjkZEVbkwMudPUIeSHBEEpJshyS9PhOzJe2l/E/Sb0XmgyzC
TzlXBKrkfGZzk+H+keVb+lpmWKh4Yd1rnOQ3TwYWv6HMmoRf9CA+fINGbRyy0s0l2j8h+6joRJES
7X1KznfVb19tW8rcBjF3tlW+lxx+iumV8W6jTMc1IOiCSGS0r9kEJb7HhFyNGhCWGqO2FYgdaRPb
fH/Q13wXIbHAe/JtJsCjBZtx3fSBbsXPP8XHmROMkPvAFkCW/9lqXqRYCP6GDsTE7vIXTmyO5dUW
nu/kiAjwuRtVdnHgNe7xcS41IGEnmZjCN/aNrI+WCnruq5/Em9tRhKTYdtG+ayosJKiyrVjw1mQ+
BFlzXQ7I15qnxPDE9A2iRRc21V478csO09ZfjGifVKiWcRHFHHBCnIWoncMf84uqudDm/NWSoQCK
Nu7onPW2FIAnln5tf9Anx2WQCfGSPCgyWmwWabJNT18Iiv3YaYvmAxtSt5A5v/watK/zBeth3+64
qhp29KJiJmEldXowv7gPGVok1I8MXVKMybBlRSqdiugGyDFBWXX2cgPWByK37AmjpbJcEjzN5L7Z
9pPdzOrHr2bTyGBs0vZ9MYpbR9pUoGgQ3Sb1k1mrJGa29by7e+7xPegzdMEIFMEuUDKQgkRka7dy
kBHJXykHwkxGTmLQj3pxzo0KSaJcd3inGu7EdWgjHr+uyJqT/Vz6Q7OfSjZCPuWE35OVBl9kK5ZZ
jJrVlwi79t4lCDyiVG8potXvRP/AXQb6zY/UXPpZfF7IUI315XqL5IIUaCOIx+9XMa+tqfxjd+MF
bCXOMFeD9TfkR4lXnglaqZUsl6pD4tl68FX3R4xQQ/QojtH2FasRnP6R7wP4G0MA0cx0mOBXNhs+
79E1q/j97j6uSzCN7jLSDNbL0EJe+4a0mezxsnrN0PKJN3X0olIUkl6U1rKrllRmhbMjsphkDWsn
9mGQhQ9MrGL6DK3fiM7ko0FuUCSRaW2531CwdC8lmxgqzDt9J/BmGE58C91HwvHSBFghQy77CPKz
Hku776NR/P9YaDtZs6ttiJzVRDatISgIhPs9q22rj79C7cfjLh0tdfcgh79ws6b6U1D7BQ7hXqgN
krOgYWrRONDDduKQfcC6txDYhA2LhnwZG6vU7PPBM/OcTq4/U5sUcWWchtNYUh4er89JZOr4/iye
wWPS3VeAypRd7OcNCW6jqp2kSu9T7grZgB722QOjz/VeP4vEShkZx1r5/fvvD2ZHeJRcznytYO6U
ZAJS4dX6T1KsGl5SkWswOkzJ9F1AW3xDFkki759YQuATrXSfJRUK1pOaB3qmWYVvk9q+XVxjiGKb
6zbboZQ48Rc9RvrpVbU07mOZUvTYKNAmGbrP3Pn9yxV5ZLEaNFLdEeuYRdJFggigeWkjRLQMMNXl
UUa1X/Wsp/pgSYXBkOxyZ4mL686BlIL0eA6Q20E4CNseV1RRrkoBSPefefHXQa7sBSaiXt1f7Nme
mysCXOWjja2QhjBqf/mZaaW3EyHsArTb0Mozp7J4lxCn2UJJmSxH/LYv7xx7D+vd4r87CAtq+zMX
ricquQS+kGCGoQK/VMysaSPOLuYyQm7PyGSccaCKA5R2rJg2KNYb0BksQh54xwl2jHG5/xncvUSr
7A8HZD/UMVSRdVUuO1fSMieBR45HOFQJ/yRG89IHPFECs0Qm2CXRfqMnJ0yImFa9L3gmILobA8K2
Kkh+coYFzrxsqS1+F2yIQgfOAfHxLM2TXV7up+VBNPtP13X2Z3+i+kRRFf0cFyvMsxgL4/Np4GC8
Pb7VOA2SMYnDty+H+FQ11pLJMRSvAU3dd0E1/23JFVWXTr4A0jw7k08MdCVmdCo315w9G/4AckOr
AHx/GYdCfsKILmIn0/Tp7DYlT0AbQUdU4qBIkiERUdJYgKX0t2OKpN1zUCLhzvEVwQzfxdgySJNw
2OEUyXqu5+IkoVvuNWeBdItqdtDCTFKlE5UCYRh2wVyRflJFZx5/46C0Gf6idytd2ZAUWp5XlO7r
RI+W7ibSf8gTxHV89M66atLrOl43smT6IitIYMQwxvoZbDEq3p3tvYzSV2qQ2gk0wMEhyMCkzoid
eT01pAf42qNA2Lyo9MSdnMpfTO/gvM0uPPsSsIC4OovbLoLTtYr3ma5D8eNnPw5ZLRZ09dv4YmYZ
GEtBZMx6tPWEP9v1+OJSEgiQvjuSDgZlXdpXwLy4DjzF3bFSSG6fx+EZlGeCJhDNUdyv/dZ2Fm9B
34FRikCexWRsuhWjtBrodHDskyYoun6paPuZPg8L7j0wNXivmqC9sJjlfXT/xyyyTFENzj7EUYFo
parYwzgpy7UMRCsyqlD0WWK0ZVjflzdIKeGwEGThRYCUUdWD/Yu5NxC6isCY4AYiCsZ4IGTzGx+X
MHj1ImlWFK7Wgp6J8HDYyWxys6DbEow9bP7BCpLzunxPsiNXFG3bM34tsT78A/9xG3q42IEIRmyS
nWrqqlZVmG+ntmIeVdNLS5WLAKZqxnebNFSGYpg2ax5EwV916olzRWV6g4y71+egBOhDfjtq4Rnn
h0Gd7jqu9NCnATHRYBMA3Ss+V9LPPf0+jhA8B+vbKL4fOLqo4lBNZE5L+6lYuPU8CXV5g3slM2La
pWIS+wNWkgrLeQPiZEuIEX67+r5rRFmtNR6SnKLe73VcalGTNNVzhR7nvWYVGAwqQP3QlxEu1kPK
mmhUbrtFHJHRdrC3dDeNNNQ4gKbcxwiIgMXa8OVY8yLyw2APgG5RgMEpWojDnjocYfkiubTAiSAt
BGZ83jsFHlwJMNSNIuNmyqF1uZTgFB3aOdNBHL2SuPoZ45gLCd2vtYmKBbHaw2QQ/W1WVdN9hwVf
JgSme+MfcR+5fyMem+iyXZbI6oUpbFAgJgBYD9wZETAS4rjopuBCcdR9a/Ub12fStYjpBCyES/ua
IpzxmePR7L5VIyiqxU1GKFoYZRlLWmaZtVbVOowGPvPzkcNQs74Vzp5B2Ax9jXNUNaM+Cn29jrwl
5ao9vuoZdmbb4C0Jm2CWVXqN1q1bl5ViPMCxVGrEwXRmP0cqDINYjbP97YvKDOSswvPhj7PvzPvI
KTkhaKpJfndTQwXvTs9HkQ9ZtrqxAzZVqYz5DvCrJf4oUu3ORbxRxMRjbcdBOaY9mTY+JCDAWFav
g78tp+jyNsliUWAupBZrt4QJCRZd/T7mnJThLUlqnljDJrAlJ6FF2Lb9Ym77uJo6CWDr99giPTn1
aZZj9cWhXr+ZiJsqwRGLn5vtyY3Z1GGHRvGpqJHtAINTxVnIo964rPhsaGuDJdJ2usaeubbFfgGQ
+ujBc2KOuxCsZj9cJUoFTeLX6VmS6+XFH9fgYUgDMWK7FUY3QX3GQ0k2dqritoNvkM8v9VmyLFQe
+PbcSR7UaL0i8I++LRu2I6QchtVENl4KLrmSDf7TW3f+gq+oyZx+zw0HEA7+kciwDkq7d6mZ7z2h
Kamptnl493UboJ1M3FtgbcBwgNTuwOfqQcJfauDodwgThy1GrEL5bEQlQyTPhBwbMLbDMrEQOBrw
9N1d1q1FeN3uJttGwtyfwpTs5OUjvqGTpXn+LK2ceKeDTiBJPwG052Qhn86NLHnIq7EKUywaVLt7
q+rSX1kwImP8/fyDcnxHxsPwZGv3Piq9Nn1B2wyWu8x57n/bSgVa7xmZRLGdJ0cz4qe0WCwSSjZD
0WRyis0AjSspoEyBOxzar3xKNRB9Uyo8Qgprt5R7UOXGtRVJEJQVrfUQ2yDxn5dApJwjBjsnsYb6
jto0IotjL7CYNP6BPg6QaBMhulWQWY+tUi/dvu8Y20PLoKk3LBnjFab1at5LTt7MiZAqkovSXHzc
Rg7IEWOeRfE2ppucJ5ucXQNmCvHUoev7PWaAP7cV686LEhsimWMso8qkh4ob2922z0NGgdnQaE6u
dFF+MBQRpXbWJJepw/7+7qwXgenC6MYWD6D0Zu2XmJN0M8/4uVgGo12fOoaUYU6PAASSbc26yhIz
vsf5m9KlbcapohR+uw/AF8TARX5dtB7TE/jxaF92DMSP78VeZ4urzQ5waVhf4NXL+SSI5b1WXKWa
LItmc3UMqkLFabjMfFRZDMb0Ywj7vkJ1se/A6l2++wC3/RHTyK+pxomVxNQFvlKhVQHKDRQuf7YR
F+hnTdMd7nM5VgB/qGNKSCG5WuxDF1c6AXatpywUHGBxS//FOb8lU5oR+/i9YYv2oqqmOl0TEgC/
A9T4nP+GvzgkdM+b9PPY6OV+THt27muRY3EQwtwYNhTZDW0QZMO+R7+oKh+C8upRMvv424bNHUgm
MQJkkam0iYfRU4o8mP5mkcU30RhJUpsVX/s23n18nqSJOzDZbpkr8WTqSInQjDP+Q3d4J0IXMlaO
ZtFuA5w+JZ9tKbQ57fBGuRqXpasDUFJ+/2UGfPyDFFJ2bP253aVyFlRfyIMMbfvDGEKC2kk+n0Ej
OOIWHOfRvfhKWLtgFrCl0bWPDe5k1moIy9SyWrH9BmKb5k26mIqWJXnyWJ73EQmBsgC2IhmA4Ki+
UPnh5AlaCODWJKiGWLbLyIgF4zT8Tje7L7W978eNcnqy+iW8+n1K5pL5irmyiaFRoLIrZES0H5K5
yxsGjvc3MPjGsEEVSwpJFFjkIt6hXgMiXOCKHzeJkzNZuZylQU/0b7Y0f46d1ZZ3TgjT05QyvcQA
GoU0NWhJY88x+61oaPuvdKjriaPOnvxLO8y3w45mKBIYNOUubywcKXB+jimC7+JJw8EbwkBWEdTj
cRgYhGxO78tRGYIZp8UBO/sirwTB9g9JIauiBrZfKfBGnAxIlpcwL653C6P0SeEZC99DG01WKeWv
/K8rJxeJGRyWD8DinhQ9EJYDnZsvVsLaZ+0uV4I/G1vVDrYY45oQ6wukivjiLNlYX/iOEpkVry6J
v0MYxpDLUsDc1/9+ArPDKl/O1lHlNLyIlN+QSKvycj4uFqiDLJUhBeGNqqWEJ4icNxiR9ZfZJ6sR
GG0Pqtudj909M218pDUD47WrGOEET5VK7MwDD8vPqG9M+jmzOwLafJz9NmRzyeCtC67z76oiJN9Y
QC9dOGzFERWzz1AX6MPPy5fAUjbuHcz5UPemyk0/Zk4ldOgM5XkJvTrmfeaDxKq0OdTE/YKQLfRM
HjW9CAX664uh+P/MGL0BQ5EXd2iQjPFAECvVp9KwpyxpSxlsU7HTQ5NXL1xIDeMkkxb42ZrzjQIp
hUMDBXcm3mz+0XMeIRVUb1jy4lXN0Yh7ZfnbWhN53PAh1X02+ERFs+EZF215yxI/P/Aar7EpDI7c
jk/frEiV+7M2UTjuuqNPKmEoxBXuu2R1E6/BNmUb2frSmnn6yDhlRl/cXhlOzeZljr1UuDNgePCo
SjXm27EBjYp3YaPBIgmR19YKN8j+WqedvEnc+oySqFiTorT+QhGOg8p7sdQBXG+1kjsFiUHOcFX+
r2+GeBizd30y1niFht/YTCci6Ce0gPALollyQir8RG52Xv80uxuNlGEBrHZTexRGgjQqudT2+CSa
I60JRWp6yB/dEpYUZLU+H5MwKXtWnp9SRYMYXOuahZv4FmuA3WTRuTa/2R8WOlYGAVuSiHMgF50d
Q5es41SLN16JBfmj6MfwYmM+FhdNbc4y10n37kZTOQGNg74rtyIeePpqGqrzI6+x9p59VRsVp+eo
bQ9140P7IxvxzDEQBz4qMjc1hr1WPxZcQamtsoXBfvqSJNLepVmUUH9vo9m4nfWwzIarJnFNnn3Y
YyAQ6Q0VqPmmELakvJNxVZx2lL/qxQp0Qw/ZYSQGipqycLp5RDH7f1rWXuqingUx1TFTkBWYR5R/
PaKIF0fq9/stiRCIyVmpO5ZrGGd8reNRnoVXjPAWXAwVu6PMM39xmOdpLAguDHskq4aPwP3qm62L
BQrxNWCZBRoM4qYRY/YJGfi4IUlC7+icbv9ke7IsEKxVsnJJynvkN1wbxZ7GJ+J160BvDZaL01vF
nbgWrvh8ijyJIxrGMSinUmRVwVuB7VAx9szofi60h0LP3ImTtaXZPPEn8eeiazBWz4RVq6qSeq3v
HSt3/FUCtZCY4DctsysY8yVzh1E0RHW4o3GzJjOnGCe/d4N0gb9pqA4kuLfMPecTDZdk8X7MYd6i
C5J/YI/fTo/dpLjqrBd88vO53rke0+a7jopnlDNTGTsvlush/dppnBFKEb39whW/USuzFTbewT+c
56motm3nsmoFev3dvu9c/2emiRgLKZKuM0GdtsXVoauD2gLrA2P6L092MKCzKvam79TTYDXblS+E
rhhKELQhjFy5eK/t/C5SXvcP2VCepxhPzLtZhFGU9T+sVqtrlqajdRiFuyTnLDuH6dL8L5Rrmyjo
MBkF58ZDzlbv/K0HXwfs6h1MxGuxDopu00ZsHyOqC/kvW3dCh2bRxiNguZVp9rmEjF19aojbWC9B
WiO5UnnCKe+XT1QqZpL23jCdvzPRumdsVNvu8nIKBKJ0ibxvGBafylJ1hzgU3Ofep+zTaIKYUHh7
IryFYU7aHXDeZhQ1fT4FYOKj52A4PlNIk8wiSpwnp43bc3rehaHHOw7DbfiU9uJUJdaT5w++ZgVz
9ZaxJ2oWCzhQjm+/oyVtDPY52v6OmdumpBxjmkg6FpNhbruZjcQDMvCWLRX71fRmgsxjCunCMQJs
XjMTtFEjGOGW/kmDrIfE0Y+Qo066GnGsTx7u8lm8KRiNoNvlC1IU+uFbWnjxOzTZhX3oaEs0konJ
4BZVBuwrTexobd8IhwminJZMVIgX2o5HlDbnDKAvqAu8EgkrxzLlQiu+/RN0lrWAcDW8h6vZwoNx
Pd+ymT8mHtKm9OxWbcfXh5ylObjUtYMGwhUn9bcL9xjFpw1sELFw8MNvFFi0QOtVbjrR74bXJ+Vw
7n2l7DnFuzYP7JNE5pa0bt1zNHG+XnbxHcY/tr13XT8BUEUM1F1jDjX5GGfNFoAHTpwvvI/i+ab3
S+yS/bhCzBy8P5g1Z25/fv+iogAgWfuB8SXmuIfMI22WDChs3EzV3c2N0b/MHQNIzmxCl9H8+BPW
TF18HJ6RDrc9V0+3Xr/RLIh60AvmQl2zyhYT23jcXxU18u2vj8hJDOsQoPQB+Ok9LKni5NCVyacC
yw7eGNjhsuPqcQE7hI0dcP5uDrVj/NTJ55XPXQkjyy9NP8aWec1zayCAkJtv4gUY9kUZn6jR5emH
Dga+HN6n7HdtjlJIJmBNuPN2OsE+egR0jylzQPdaq2QIieG0gpyhjyyncI7Qx5/Kz4Gk5+l01O8J
EmqZNvTzRPbYjotYHriq9H6ImLZ8wFouYWVpkwfBkYMxWhMLUMfYEO8eae8PW9dfzCAXMpua58P1
PfmbCn9Q6f8KLCHiseEeGkufdC3DhwRdUB8+zUXYBDBKoCEX2AUilhuwXe19b2BMgfhn1RlcOVmM
SbXK9UNFZch80VYRcWP5jARQkmNZQomHAqkwe5K37gRiA5Umac1N3TNaqYM65fAcofic/NLW6Ej3
nxixRB5/uuFYw0bFDvb41dq1ayfqLmCimvZn2t0TGcSr76Q2cqWo72ks9Yz/nNJ7KdZENddOiHoS
KCmGyswZLXE6EstW1CsYep4K0go3Vpz8oFu6ANnaq1XybSwbsPy5u37ioMWM9YyBi16Aib6pPjX1
gJheuBZ424ywEr2in2ESHqXY2lJC6SoSSbRXgNdsb78oFrnMUSaQf6KfTIzmkjQ9DLDtPyWvdUlv
IsHBVh827KUWEx8jYkaBh25kyI8ohAZZJ1IZjWh0iep/rtzRHpspqUQy9JtVXWYHeUEbL/xfPGdS
R8eSbjkw7HFeRX+8dwZJOLC45HnjifCF6VDag2iK46nhQj+t6Eh3Sv89C6NGKKoOhamgcrgPizOb
9PojtG+/qmBPaw1hVYmTpoH1nH9yaQOjr10h0T7zWjyRlAwn89ccUgvEo3+FgRghzTAuiClADWnX
VMcrDyaztnYEGxMYZF2JWsJpc7qHeUxLMdXGyrVQosAdPTj5sZ8T2RZThFDUVTNoFk93WwPJz/xS
HCg7WdmnhnEIJHvOe8Tq3hBd9qJdoJwJIpr4+gY6Tm3k+yl6FTfAy06reY1PT5ijZEAP5zCFaG6B
Zd1QmQtz+vg7oKUE8d+P6tMa0kt8cc4/GtuUmG6I6Vtec9FgfwlbLdZxGl+wzwLsHe2sSDs5YOzg
qRrEg/4bVEVz6tTFkfsvt6ogXDZxI17gzBmLYwav6WLxa88W32V31NSioHL7/q+I/7jHt/fb3BYR
SsjbigbT6GdNPv4qAV6XrHVzmKq6kAM5TA0NBeAkqe5ylaAMRKaXlCETS6ZknJIjIzf8ANs51oFT
vfYehiOI4nlXhR4pWatYg/7Kaa7sypzEIqJWu3c9AepZest2ilt/nnvs/l0FYHT60l45yH8Sgii2
Ql7m7SWyhNfpbbWeznjLFLzpLthmKUdM++8HK+Y2tZ5qaxUx3CnFgTm7126LxtnMnHPiXLCcDRH5
U2B+ObQGYG+A3bh82kjwPywPE8LEOHOy7+r/Gdwe9XP5kxtiuztnlWbMUYb21lFtIwarYMSwq0AQ
qDbvfyiyXGD/RwoqyLpdH/PSq346z11n7gdLtu/iSRiqPZL0FnFowgBsMR/BuDE+PgiTwT9DiJL3
MlsGzQTPHlVOb+qgVaERerVkQwgu9g1UmGN8W/SynKFWAIMiVgr4+ULhF9uhOEEp35uKOWckscs3
IA2ImwAc0qmNCe5M5Hj/6wFYzirBiYwas5nKhdTCKpSJkZAmdit+1NShe5tTmBo/S557Qe+qqN6Z
lLYswvv2XCJhYcDYOYzUuzc5dfmJ0DH8Klel5UIzAcAOzcgX8aoS9o95u98f0Q5fjjVB8/taKuT2
Ydan86uHskx0jwPJbX3xgkM84E9msWIaMulrfuHJRncg19ZF58PjtV6h7FXLcJE9Ve1lsbKDfEwr
o8cRd9WoM9/41edOIwGYz4aTKSKbRdvpeUh9wiTSriQ4zhga0xkoCnG68KcJUSe+1uIPi4rIL7g5
0aHbmahm+1qrnatvWp5C3PjcqR5XZRvsjzz4Nu020ta3GIJNIQCP/GaeDL7Pxnr6jsXBS3dJqUzu
FTWv4o0LxwTate0h1pgNifjmszKSImUGOdl9Zy3G+jaqeZKQbfMvODz/nQePJJeF4Xk6cVefd1Mh
rxTwnXY4YWWt1wkyfJSZA0/ym8gmSZuItLXXoAsEKnpO22svGw+ZS1Qss4+Dh2PRQUNg5NoGZwJo
7bWh1RzGbShYHLgsJxEuzqgzv2gIVn9wPbwuWlox8ImyKD5s9Y9AUEVlZeLeAYYLUcv+8321pqNE
ib4QmiVAI+bh/rq049prIejm7JL7uKOCl4XefjRvvss2Mwyr7Nmbbusti58JUgVcraAR2GaRVPDC
cs9oTXfyMOK9isuiFi7Vpq5WFTEldiO8NtHBkQw2H1n3RJNFD+uu8r7ewBo0IAwmsGuwJR6svcIH
X64467gCG3vtbcwK6YkT9VGAkPJzy+4KEKzCLDZBnlDScSN+U+IFGlfQxJNKF/3yHA7H9AQbkka2
xLTDToMPW3EgmiOTap3pT+qpcGdzfxTVcybZ/Yzj+Hayy/Gvw9HalATjvTMN/xBf9J98PzM0AzC0
63tvX+wFv2Ca8Yn8cs9xaPsrfmsURJ8t0Pdal3xwWQD8rU3mC+SNVxHPqsI6pnHproZkHn0+QyM+
hqudS5OtG5HAPSQti2beFJivV7QlpRe6TEaJOYdAIt4ZSDToKBpIiu8rvZ3XUxcH2x4zYeeelf5m
OFt2jqVr9uLzX44JxKJy+N3/warU4HDJNIzyzhe2jO1PZHFyJNsoYCyMJnVrBf5siSAJk2um4oh0
SK2FN4C95067Vq6NhWmDiYF1WW10LXl5vrC2ug8CoSQVC/atwH439z2rUcw1DtgDu4ZA/gkC1gOG
qIbVG0cYpWsYwDYIrLMOdjmUh9hKbzLCmNVuQ+XjDgJkalpZbuo52TRMUK0flDTr12DmzkNfmRwH
yYVqMWIXKtTipgVgGsRQtbyOcnsa6ZrLNVl5RpHPfSprgw8Bxk4zVZl/CuIGZ3mJ3APKANu91l46
vHPW8nJBAY/x/Vc2n2Io51aFDbJ9DoUALz0A4F4MSIuudHSNo2XuMqgCGZjwQ1uRnWSlJCupK7SD
ATD9qHbUpwWbnF/B/gJ8VYKU0o9LWbBMPoVdfh3SyTnxwhoiI3qv1ZHwX+SaVs7+5UG/sR2XY/al
cwHMCz+L7vLEMUMqpnAGLHKLHhZ/5i02gLpp81ALkboshRnJ9ZipIq3d2vxl2X4yJW1Bm/lrGKhi
IkUkRueAE7j5T0mofLW4Trd470QK22GTnMln4offGzI8i20FoLc4hT0DpVFpc93quClulPA9KbNJ
dWZJE1E3gHJ698DGwyarxqyVVjwyx2sKDf7+0uG2QPZNneMbXxm6TPVwfTBMoakFFE/Y9wmFlz+B
7h9nt9+eZWsozz30PVqE0yxw7c8TQBUxRyEPPw/rRu6P3pABmLNwfPWO/KWb/DbQ3dROOhhQIP3Q
YDje1+/e9J2hQSRiQfrYRy9wWJpTP+0FBYcGoYDfPBVq53Z5X2G+/sn62Dpwiz3nYIaoWk3Jmksk
ekBOtZujzQcitayZdzOdoxVJy+JizlMVTyRnOxzh51U5owLf4/ijRzYqiDq/y/SNQrNndvEXQ50f
byG2r3Y+W1eOFW3lIyZoX7q+wNSdmAR81Z74aLiV6mBzy3k3lam+8GqMCCwDykmSX5i1F5cJ04LU
5c9xGtlLYqEWyu1RjtPYxA6X8ZIRS5zrIs7PqNopk3cLxWqM8GaKE0WO+Xusy5S15Jg/YamkKOH9
P6Oz2IXZpqHhmfzxgkMiTnewES2pxrib3+jAsAagzF4wKIQ9RTEbUgrhliFlPLeCiE3SBsjf2qO+
4sLPmv1c5O6vzfLKd4XIO6IOumkqK/8S2hWcSuj3kvk9clNpdzki5M5de+lZyKyvDBKRr1iRrk7D
s2QXxrOlyRVc0Qe5e0ORFu/wjkCQ+9l0lOwUH9ZX0QkHWsB5LEdzOd+n0n1Ci+2uJF9hkwsL0zZ/
IIQfw6ltIAst2hpTRvysORjGUI+ypXYilVuGRzbTzTXhwKsqQGOWnHg5wVfsUmYV+KK8XeCBhlCW
XM2SCpCVESt5E+cRodgFvs/45Ydyg3e5UFwwKZxke1cS3Mf/2dWySOzBp7TiWH9yNt6bYFr9v223
Iqj31+/t6Hi4L69FOaIQjmW96BCv0+CD+hmXYTYbB86cTe4sRMYCq0bZhaVgnZ3cAsV7oqfpwgyo
ECJbtjZ7J5hEyuya2RC47s2D02bkpf7djxGw3aYjwjGeKgrIDWsTSjwJQygRudYPWk2w6RMrWRBz
7kkKtXRFzlCT4Ayr6EsOJMHWAMvgJjcnSnjAaNwShCA3Ix7Aku3OeWh7rPh+Eo5ui3/2/kCMnDvq
VwHQRWGpcS+9Sq5BF33mLBnaxaGjO6ZwMA4HLBgBrQWWGKnkj9l1+G2kyL2Au7hq+AyAVIkPz3DN
2glOsoJRJDnY2QwHfkcLZp71mxvCLr2KZLIYJnHDOWUcteh8qKujxn+h8GSTgTBkHOp8t7pG5Tt6
QREzaHCBFT6fIUSxioFAMhknSjlSNVnj93ZSCgCVEIUPRq1VQ9Fjj2z1CSbMw1AWv9ckwn+5I5/v
Td/13/Uo/JqsW9D7btzpgwd9Ej+KjNKwNJcr4eHW+ubyyb/Gc+8JYxriCLNlGFVLHs5dNeL0qC9K
qoI3HN7h3ZSyZPY/i26GbKwkJWEBAOstajOmwrXVoTmeXdp4M4R8NEfYEzBaWa3PwLFXVRDwwQpi
qt1p98BqUMc4zqryvfDIqBiyISkhwKF2ZcgnpU6RbXJlYsPk/HwK3Khbn5MB8fdRAQWeDiexGBz8
GwBYSEeezrPO/Aug/OyshaWdrYb+JeFwngb0g+7k+VxcQhcpRL3t6DSio+Lah/TsrDwGQjv/kMY+
nwZnq3L8cm/GvOGIM0aoilMKEhDuxKcXCZG8luqM7cSe67Gzn6fzb2vOemMReCUdRr95nEhFxXAc
9qn9aao0tZqTK8MzRhUf77YR8E7YwVL+kzXyubUldhdtnEDCB5gCt40X0Aywo5S/Art2Bpz0Xsi3
3YdyKL4bj9p42f3Iddlt4ZR50bzYIgA3msT78dUQN9UYsukSoU+fDHieeK8rcCR+4mKW6eKGgZFX
ot2Hjmdm64x6PbCyQYUKZwKuRpV0xCeufAC7zcOmQgnJDWivcovljJvalDDZwuwiHxjep0Q2f/O0
wMRarqS5qeT3nWXQElDBVhIwa6m0QCVOcIFknKjP/3yJj2DU5v0NsvyjZGaO0JaJGws1dZtnPPoM
LrdpFM6sjwkHaSaj5J3bONWtfQJGbszAih0pqGS/iEYzNV0+VqDRASeK1kzw4ISHho+aLYxg7xe7
uHSGkUxt9vhsTlGhkXdD0Iy+ltGnUapqA4nUlbr57bmKQmMot55b4cVY0ZNbbXC0df64J9BlbAq8
GeE1CmLxNJ2GmTmER3D/sGMAzr2k36Yo8+3m5w6IM/nR6oSgyaUGAOyYRJt0BLPLXj0iZdatnYWA
INu5+9vSZXIjwiq0uRlKTaKZikuURBlbDsDef//puSD1WMk/zVDqhxfl6PHrjrrXOpLPfQS/9fI7
4WYnvD6nUyeUSabVyQB0gIQ36/rR06kMGJSgIff4VMtDXuM0NsUKQxvU+vFNDANkj1Th7sZqHaaa
W/xr/z9wBc6jaX+Udn7qAk59lz4/jJntOJISarLZQIWxMmCKljs5ybF1TBGLfKRYQDGARey0+G/N
SzuxrTDEf10R1zW7CJ06rVcWJ4u//tMyMazpp91o8tMX7a/Cgo92IEM/YAbNqiojlUHJZkZKPk9C
+Td93yRkezrVwbllvxOL+COxBgh1LJd+LJV0Cl1LiZMAF96IjF2+euDqf59EEAp7q3OEEGqAYCN9
iPaJp9J7Yj5DAgpGLJtAnC72rwuf7BTEAz4p/qsdH5kz6shEsyNaTqnSOoEH0BvymFdMJIOrElyh
HqEFhOblUGytnxnlaMObycgt2Weio+khb5ZY9EFwmFb7P5LXCbalnzUehC4hOQYmlqznRFD8ZB+p
8qcQxPStfJLB6eZ8lU16cCq963tomgdMAZoN9nvWoQNf7788Ezcd81X+lSQ1WhrVasNlSaJEiTOR
f6summbriwpI5/d6Ec/L5/kp5RjG9B9U9edy54ayyMTmjNRgos+LlylUUAijkN2bY5K8dM2FUE1I
IUt6EVTDAGhY5/JAuvlwiUFJ9IYVuSv99PvywNQOjidMTven3yAS38fVTH+EPzpKAW7DECSfTX6+
yBub765EkPJNGQgaEnnMfTG8jTM2Qf2hr4jCbfLgl+GNBBewK/79YoHW7NIIYQ6AKPDYu0p2Eq56
1pXLws9weyZ5IYsheOZhw66Gpd/yrpVc9Xda7qwatRvpNFFT5fdZXV2geDzM16sGaeE7a82A5Drm
kKfooBw/nipE6MdArpT0tclcGI5A7VDfi6WSQyZQJzXUaAojPw2tEt87riY7Hj+Uk/35bdkn2kgQ
/ZciedJvPDL9Hk1VOL43daSvnOWchHycNx3WWBWABMOq5xKRtl5sNwLOvwjD2WFNmcYCju/8kUyi
lyjOWuwwuSvzTcZhvHJOq+v9Gwp422nNPGBGNonbdUbupH5aMb0IjG9kue1ASh4r9/t49QYmTUOK
m0PhEHZbu7bgihfD2eBSgKPVKMeoGpX5qBx6Dlk1Sorx1Gd65miKfknWHlLS3IDLOeVygE0dVyFe
iNqIGfa3Zoh5aqgI9qOZgzWhvvd2TmBzpAnLAWYosfT1C/QjaL5FLM5ijqxD8AC1ymINFcImOW5b
Klkp/R4w28T+x3ylS/b0McZkBaTY2g0lMZxkWADsEWpGc209jTSFsCIfrpAy/bxdWuPyTf5queKp
mb5v36iwgRauoQL66oOKbWDnE3OOg2JvWN1Th/KZ5EQ0awYYKe86WifokQeD7pBsPO8ZPqPyQIRN
Ncmj7m0S23bCgjRttl4vRRgSmJlQsSpiFZ732egZv5t/59yGDmWEAs/ITNAV5SlinJxmeG+BrK1c
2unxiFWkaMqWBfpPg0NMx11ggj127OCLcLdLrGb53PfRh53DUxPWFmK3YXMzIegZKHYBp/DuohdN
cefJ8CaXmAV1dNcfEehlPOPVw5uw41JKtKh+TCsVlhsV9fgGPKMkQPAe2bqzRxNxpHTvTXgdL3Bq
1mIRWz618mtW3JVJHboLhpRFPLr4On0NlvpNZvV4Y/jzuCR/2NqosDANOn5Dcbc8ItJHgKuJWacX
e3VhIYCgelQ3I4WZd61aEM5lH2Vbw5g9a67rxfbWKmfAswrhq7Vs1A2aQpFMMq84fCbAwwSoHzIN
IE8LAxmaySbwIMd8Vo8ZSdSBmjLqN/gcR3ikjfNWgcwqotZP5kC2SQpUNnK0bqJiRgceRlmLjZFV
luxBYqz/x2FRW71LfjbZESVXSj8ad0bPRMO8w93Zp0vybyZXnGtOy14vN9UNx0gOnwBNq6nlQAnq
sfw2iEe3napnPx8xPPRgiQZA0tC/Jcv+n05ZgvjxvnyCFbYakHq2tVyqVGRuwP/QDXEiAemYqs8W
Uar1FA27W+L44n2jEUvKVDpqDg+wgIDVZsE2cOxq+w1QMm4IjPUhIn1Fi9PyI3TBQ+OJX+ZZ/hlx
Y5O3Cz0vttkxsyl0Js3OANa+Cbmb55I8IhGKRnz/TNICNLznBZdSuzAyHePeYXErATj3SSWdCA3x
V2XtptbU5RREWXVxN4tp40nS+HUBzpijGMKyCZMOBaHdDCV1NSO1ZEt/lPZI59nH4i17v4kGoQBC
spVLhVLUB1s817aQk4NxeSwDyGGHf0bn59qL34bufXgAUL4BOiAngWQlEYfzE6r1DumMEPMAnH7r
kvcKHvozcHjFhDZydUCQZF3ZjQslE2E85vQPgk+7XecHAq97kVadId+FH34hCcx3Uanv1AYJzLa5
hMhYhVArXsyGtSoch8f5rsrZq2Q+H09cU63N+rhhrhYZauq+0F+NFJmLnhnyHGG7vYKVOhF0mMsm
zgkYGKEUnjuzxOjollVelpngmnJDcwvx6M0MTEgs2efKZJyCkQaFdw+T7Oys/bwyShipzlIFo/4q
tIR4LUfXUpRRS+27x5YGFQeNiCWiZ0Rr3KRRLBxXlyn9FbsROlYEoxudmiZY8cE8cfHUv4DNZoKB
/vUoL6zHx0t7iUWH11XAYDiQq+8sHNPYnRSqRoz5bexf5UGLisPVgfY9TTpO6eLx6myqDqh7Nadj
5rAjo2YGUmbpr8DsHcvsHNdMFl54sGQL5L1xj5MZdh5x4lEajO3Pt930VesqQdurCXcL7Bk2oLpz
Wg8X7Z/luuU6shw0DDP2PS8zwWQ1qN3oL7jKGCUJzFS+7afbCargdyi+UvajDaogwz3yaMc+MHfs
+gJzUImFeuStuh/wFsEUjaIsdLs0g8xXkjGf2DmqGNd3y1tbvWt4q7GtC76mjrVL5YIdIKCcqGlq
pCEZkXzjZ9o2oc4N5aBVjWbsYBgjNS4RMDP/ocA6trmRUa7ssmIOq1MBtJf37jEYGdjwlPfP6BnN
yoycxy5efisxU1v1+EXNdVpq6xegCIkXS3GAqPSAx3ZIXnfOvxCK2fyaGVPorSpsVE2dNwcDULtI
omCJ5ZTJIS/wzs5yaEhbZ1bcEVvZiEF19qIZi8sCwxSfXvLxCLNBQajnUqkFkzjPIwCf/x/QmwWy
IyzkEJIwQ0gUFEj+LIIRXCmwCOu0bn3SW7NsF5vvAKC+xDUdK7+fsr9ckX5yII5xljg19zywo/4g
v+L/9oQ6vr9vjY2J5e2Oq7ECS4QPmfT6njHj9IN80HeANyy0o8olTXu/1/xV7BEfnKGYP3UYbGZX
NM5fRFoQZn/kDXcSeZD3vztzqskLaM/hxXmEm4sQkF2Y34tilyiiSBkh2SwG+4dPbpo084aFZvij
+W/kc3RE+vjLravcFfo3s0a6qGepjvBizZkBpcG4LTWdLS03f5VOXNXDYOdsKUqoalhpSe8HufvB
WW550A/ZmZQwGHDeeCesgStl+PiJWHTc+HMfOv7tFxlnCGp3OibRV/Uj6FMXCO6q4km/8jrwx5P0
i5qv8j86mf38y0NKxqJlj1krUA4TF5OWf9U/hRey6zs7+iQbh//DAAUGB+JKN0vkfT0VKgh2lYRR
jHxb6xg728X56DZpd5YsFGveighl84i6SLEXrPVGC2QbZml9WaBZztoFkuXoVx+EmVkoOdz1o5zg
vraTLUrMHi2aT/1902TDWzPpQDf6UA+YSE7yYT8Tc85NgFnW0UKQ820yJCEzVuOeozgdaAvRdvxN
piWwjS3zU+O2k6leimZ8bavT+C60AYRYyQVCjY9birsVKreoJ2FsTLCLmqGui3fTPs2kEONr99Uf
dRFSyMdf03ek2TyyDTrBZ4DPD6v1j7n0fdR+5jqnqn6NT86wUQ+tpnetZBwprGOwSRczHf+xQQhq
j9Yfx5+zB6WjwMb7Lb8pFVSH46pks5YvMF4p2NhoUsmhyZTEcQDm/9srSh1RmpVSe5/Ju/ELB2qp
HZOzQVProUu7Xv9iAbW4li8D/gpGWlQCU9Y+YDLmkugv4RbrEt8fzj1wUnN7R5gXlEaGlJPu3tOb
/gP8vYpec2FCe7inhX3S+rOFvdBybjv2QSZmEOgodkx4iiBboCaEMOZch/sKUAN2T4H5NdpIFQqD
a8VM4POwG/abiKDa8T+rZm71H3TP3vCpFspvtHf1sx6sIvzDkyf5+Ab8oEeY2uyaJHpowIpPYCEM
H08YLiy7JqEyA/lDGq+zClybHuK7FNPadrmoHPrRYrcjRoJGc3dUasTkcB6g1kt4e3liX3RcRET3
WmJ4M2JFDh3nksuhl2mI/+/LOeQxHkeu7l4LHvzsrrq01msO341PN1OypHRFDTtGEKAbMr0ZKMCn
2UpJ+luI9qs8qk6YF1qSFxGZz3vFlqRaQBeJpG/e+2SImzkNodRWcfxe8iY1x9CCy9iCrDiFlO0g
YSEo2slTvITrhrR+xmcaW/5es27cFckt8Yxf3xerf1RrDLsGJa69RyPdfdmK032x0WftBrhHChOv
Aq4hdSPc/p9aWUcVUk9NspGEkbYVYPA4t7bAlWACq/HSagWqUD/C8h/5XA5RyeErrFmztuM1mX8h
eoNNBHK4PqEI23NYLz9Oz7dgLnvvyqgnT+IUcHfzjaWLdV0iJw2uuk2+WcoZmZKTeuUeHU53LiK2
sU1rsvG6LIsbWqRBoXKUyOQZijctvR5HlKuQPIseemG3BY1eRk9AcJs0KVDTa/gk91RaR72AxqV3
E8x/AlaIcsl/0NOkJXmzxluTmEffLCmQNUWgC6Z5/N/zYnu2Ez1gSJmKsTWY5ylHisi0bQ+p92fV
TpIeVisT6+1pAxw4r0Ihzch6MWiaRlEktZ/kOLDtlfN8oknsCRnUS9hBI0RJUMZsKPgkbPkyb0Wd
m7jsE8O0MjUHBuaxMzoybf7oYv/T4U5gP+IkgVjUKJDVzchYqREwwSpCmz3yD1/abtlSW7vxemSi
Ar5n7vbKiFsSEZccbSRPEcHzB/hrL+bkXB4VkaxttVnfbUJS5BTRUTvmVNvNOX69hwmb0QmCGggd
lCzlYYX8jR6cnwFhvbWeOVqPiPQxEjY21OPWkwAvqQvXuHpZnhXiiU0St12onB5F0tOlW7g+1P9U
smK3AEr+anRJZwhSaRhZ9OtnBoT8PD0GjAXM+stVLZwIFmw4RW7rApNF7y0F3NE0jlQlSCoUJvGd
raPISfPm52j5j3qhJ5pTGmLwQHzYLCUWV2I34VIdvfo3X61wqieTkrC9C4/UOzGCL82xtFHejtga
lkC0Tgy8+BHSCUV9M03XAXfH0S25cLVt1yC5TKhJVJLh2n56u/bjoVFJamDgSfBXF9XfI5G6fWXb
sgszl8+Ki393jxyACy9fS3Rx4nf3GVvrIyKubvH/gpWspJpTGCyGuODC/vopLkOxyGlAdD0u4/TB
sWxG7zyKtM2xDv/z7G7cgzhskEjXWlmhLMhEkbtpil2x3YR+wGrYJ8Ybbq9Oruo3IaufBhXWTKYD
hUOQyLlSkfcVlW4b0qhVx7YtdCDFmSXFHP750U1d60wZB7UiEaKsyuVq4T5G2uepggetKlNWz8lF
3wE0wCXLvBDVI9jEsibsj/BU/Y1tjyL9ISloEJoPfe177luWDwLsnV33PhUED3sHs6AMg13D939j
zZNegAsrcdYtgw2gbi4Agde3c8t6Swp3C83FKEn6/fy1FLO2CHBHt9/UlagMA/lt94kxfVDYFB6V
y6CpSCyQmQ1x1xEM0ABgcQk7UElp+LiznakTZ693ybfUYIW/HeiIZEkuu6xG3HLGP0yrBcgb+fei
RcHhfiZYDSk85ic1Vt31CKNRwZrPApShHquPBocmVTD/lfSRYRDj5jMoTnFXC+kp39ALNstjZyfm
sk7jCRKlFjM4+uPYggQTWprMyTboJNR6H2wlmXothIcih50zifyolW61H30zyMG1rGKDnOth2aW2
64wXJyAfZWCsFnbcKrPActl/pebpXAV7uw85RTXTEoejxmaowfv83/o+WjMcbmTT4EERM5D6VgOS
Y4l1NLHQ09GkRmL8e9VPrTbn7bXSJfotPq0Eb3dJbVZNacfa2Qx2nDalGZShoC5wPmhlYQFIfR89
rG99o3/G+RyOWqpQirkCybAHJfYvdMutKO4ysWbeixMPIn9J4iHP2TSm/CpOMDtNBbfpiJJcYFx0
8u1g2zGlhZOqXXWYBQcBMYIAyQqpCrCyv6IP5RwdPb6tCB9yJpz/gRI2ne6JOL8t+50RVqOQoruJ
ODz3lrfAezgM/MTjM00qTPA2Em2M2qyGC0BcVQ9j7L7hDS3PS7fhaXqCmz05sHrZ9Pghr+hC01A8
F7M+dEeWlsl1otMoPExGf7csY+nsKOhZp3Ua0TjW54VPOw7+9hQkGzxJZWgg3xDk1EAOOk1SJFLI
Zosfa2XltXuIi064EFi/RDnrbjBNKRCvQifI8oqDZyMUAtDR3/wu6ewrdTSyegAA43Yy967VxCYa
HO7p4xMlTebQ5CgmXt1G6M3UJNP6jhIbwwlczOeC4HsuuEMCayIWyRCnPIgT87Jq+Y6QcEQy5a6s
1OifgpfChJAFyMLbCKOu7qDT6unoYn1RuatqYMa4bv6nHiY6lxD55DHfGuWIXGyEoDfrkXsp78X2
jw0p2mY20jiD+ZVRFFKWBazihv1qJsvGzdPu/0OAskWKurpLbEpMyuL/cAt8NxK4/NCWbQARd2Eu
lBk5iTc4Ne2n8WL0nRla07T40UjdJz9RmIhH8byfwyJ3DnFlUckCTkWFjvG0llxv5XyZ94q279nq
LzRX5pc9vM3h8FchktzMwN2kOQSYXQdu4i12WE7pfVzV/CPDQ3BTdIUMWoQ1bLNlEyyjIW7itDoL
x5tmBPK28l3nUK+Dteeem2z6I2onkAQHWG62oDJbXEown1ei9FgbA5A3Hv3fgw2Ar8PCl00Ha4h3
DVUG5XRb4MsC+ZzBK/jsjvPryGPQBXezBz/yZx9c6XnIkf7ooYtzTT4mdkaiXALda4T6RPcDuAWG
LQFq218sj7Y5QMg5GvWtCn0ehO19YkAlarDt0hj/5tBvyoFbpNyqbAe7li8ifumY3QYO61auB33G
vW5pSTSkkhg09ksb2yMCH73O/C52PRrWt3PHkrI+072GxZifwOmZfISUtadIJO0Xd6jm+jJA56h/
D3/+TabgfAm0gnKCKS+WD4N0zzOnJJ0c9/Qxq/9+5TwCJyTymZ01n0uTEO8CF8YhqT9gReTSvV7k
fgimtS5w2IZAclX35MslGQx8hZ2WQHDAX9AJBsvU9eE0dRvlinP54djUkDWzTOHozmgnDUmRVLSZ
ExHL6zpxrdtq5O6oKnf3WwwUGwTLBitMIYYGomKQ1nTfKd8Xf/K4Trhg3ehlKqDH3yrYKBNNDRdf
MsuK8RYQ1FEIE+jfbF4f0NggsbayPx3ksmq97x9Afp7bMuP6Xj/LJQNZb2BWZUTlFwmIEEZvdoAj
8tbJfKRkRSI+C/ErVMZ4+jyMh9JvMXNxtKSi2WR0vNxOU1c6ozOynrHTiB+yzv3tr12diPYGgwsr
XRtUILGU6a9yfVe12RRVzC9U88VVNmvzZlK4c65ufrJd1yBT0O1ABCm8ZhPY8N8En8Ls5hLeN8II
q0YV31gfRJavh13+o4xUNfCbBb3dwfAGGeP1E4kGru5S7y/d7pbCa54NS6GQT5TyB9bAsS1Cv5Mf
3D+jt/6KBbxVSJOLxTfBp+rLmJ3w8+Tr/vKrfmDt9v8XyGCZgKzdRj5iCbnzigaPhXarQRx9NN7X
JTE3CNCr8Mf84mRkqtmdmTYhotnQuCd9mbUjI2abctXB9HwsmmMxoSSbLQ2aG1PZpsZ/gt+rIhaD
t8+Km6uY2Hwqi7zE8BIR9hsLh/C5dx8Cbjyn+q+4XKiyzuh+6OFu1mq+gF7H97ApFOqxfpK/rpca
xZaxDFwuSmBuYm3TELIX5d4sq5wqpzzl9/HVkuPBDEgfmc9KO4W7DsdVRaTWcvxvFbxvsnhB+BDF
SDdeLC660L5mRjajzkJRUba6UhsAZPKOWdheATgRuEHteqP8qp5j12Y9++Gi07g2cBP1gctwjRMk
5IVJFIMPZ8ANRqYxPBkouHG0W7CObNQXDzl4ObV3zEV7VfMSjDlyrXwq3de2R7UPg2cM+G1ttCVv
lVp5nquUilhJ+r3xKvxkXcn1APFDwk6AmG/3G+mlYlARiyjMzqZc1NJ/fwQwN/gz9YEyJ9vMGL8I
/WZYcCokv3hgFBwxy+TeHHGYpxHpMV2pgNO+oyYs4FcSbeK1zaeOAJKkWNiDIS3sRdQCVnOXnCi2
COIh8uHqVovskW5Vz5O/mNwpuV75PiAXkdBwAO0qGxATxaUbfA+8KdL8R4Rt4FtdUZ0bh/3iRjuH
20lcNe3SZV4Cs51jCOPlm7L/QB91Fki2//i8DbbtkuFZeTeW9nsRJQ13rnhQRBPQwvUKe9qmA3Kn
bB6dM5KbVlc4CM53DSoTOm63M0LSbl/AevgzhE9ea7CWBrWQck6LA6Tt5d/7OUkcGjz6Phr91wIT
VgFeXt7Cq/kgvRvvv6kRQCIYZAvP/VcmA1lzUx1SmaFkb1BrTDK/9xL0XJ2sszaNWz0B5a3uLP5D
c5J/IwaO0Id57YtX9yM1ZKi0yMzf0QDL/VGd3nOvTtRrqmMSMDlgT29O+f9xMbWQWp7tOM91a6m0
guKwsPpq43R9ZWxOUJshGAML05yPAm8UtxvwtGv+d2574BfEyXFafB/bMbu4mi3wxFL4bPSfcmzS
S+tmYePjj4cIAilwLeJA4rWYUKEpnXm7X9SxGZeL/HZp3kf0ywW1Vyk2MM7RvqTowXxrFZjm2BoH
L3v9xMseOv0oK0Ok+ZmKKyiVrjty0U0VsfvmLxqWB+SLFapDkUJqIuocHiCYh1lNO7Nv/kN3FMop
ckNWcZH0HZ2bqrt0GKWluznPG8tarsodZgj/PMs+EWgJPh2JIU794rDhLxnSMdNUIiPv90fX+x8i
rFhhUW/yTSk0IHouZAIyqYOnhKW/L8IUpwFgvajJsVETCJnRR6Qys7XmRZUhWxz54XPOBCWiV5dr
B4wSYNLIa7+EkIMAlZ5NxJ5e6XSFnnqhT3rQPSFi2++cQ+AM82KuHbFEEDoaCmFYcAB6LwoD2w24
WbYyQE3FeJpjsqOZp/jpO+rrPMbbsCZ1OXHPhcCJyYOwTEbpU/Ab1N+LM0kgBTn9V0MPWPhmsHEv
InzCuZhedovnlJ+EyBgzVgU4DBxj/kpW8C6/AfzyDPsofAOKJBlMIJt+OKZq9LJwiH603GitoSzq
/LTOy1JiarGQgBiNd0sQIsdAuAGPTaQdZ/ZtJCoSgxtK2N5Hxg4Ci6bJklDQnGVrxKPCMbT2Omp1
cd0o9gQMYtcc3B9sesluG9I+2rATP2uiZ/VqXqfuaQyrmGWqyPXSCAEePUeG54zKUmyb+6TZyvKq
m5nwlWXOsjSKV8Fchici9cQkk3OaiJQzO/xITZF6IqahfhX4h2lGpacF9HRw2nf6eapTHSqWBjX/
s00gC0eMO0TjPNG6BPGBOtK0PM7HfEvLzpgZz7njy6YnKv31s9A0SyIJC0q0d6PLnZ+/E7s1BUsb
SG/KUp5GoVnPIKe4Me5pAwlH5+CGi4GPV+wkl3aXvxTPX0erwM4wjjWH0pWBJBihU9+wP6scU0rX
q6Gs0NAZ7HT6zQZEGu93xvcUqfGNpmYq9uNVP7Jmy/cqN6oonmClimMVdVvbEAIrCrGMNmPrFN+m
IObTdJmGJNNEkWG0ENhpicm6MGKP4HEPJ3Jlkf0BEj7qeZRujgBX8o5YR1/UXmnn5B0hqsYPHxUd
BaSrjTpre5z2BeqsI7HOmLHNf3dNB47+RlH4wiB+0W9Ah/0CGfkWK2ax6JjJYJXcCYcl0tP7Mflk
mYXXP1WuoDF7ps/u2Z3ym8ztD2iYkzSmdnXlsBTD1r5nFPgSdvizXTprlxLA0WtpRDe7fjqbxn5a
3VlBP+h/0wXp7x+9u7OkA6I6hJ8mBZiZkx2BgShhnwKjmFjVQSa5hcFkh/06Gw23Qb+KuQdXDNVm
ac4LWt5KLQ0/N0yxsyoiwP3Vug+KnZ8fcFR0lZtNvb7zNIUa0a6RDyBN+MjkJRkqtmC8fOpmLqqS
7ZZQubFJXhTeQUDruuy+MCuJhQy/KSk2hITItzlMm7IdWf8RGaxW2KBmP5sMB1aCnFow2ss5Z1Ai
mxDcVLLaTKoUh7KB2ng2RpelZQngJ3oOT2d6iA9fEx2OJcPojFwum/NkqnMOW+S4KASoYTEytnJZ
xM8TgpJ3NWaYTyFQ0HOnequYNMQgHELZhnUywwxOlpHCRFDgfAfZ1YXsVKB3IdLvaJ2Kk9VLGR/7
mlyNA5tg9GLkOOavYmOxyulOFMUv8waJpeD3XqSz6wFv3+rcX9ZAs3Gu9GSC8kkTPrgzxXHHVYAG
p+bMe0sqHMtsx5Rz1QG93G+loxTmen0gKO7kqFKSp3zHg/drmuWdUHodPWXfg1T7kq6NFmtwnVoZ
k81EcyfQtXfb76VkBMQqygoYu18Ohk0AxQJCKpvrReGHupNP/8qhpXYwC8EXvEmvkod3VC8kMy9a
kydP4bJRLx7NurjaEvKEWHAZqIrxM8lyji9uE42TYtP9umpCkQgIYJW5h6+c0S+75QNRb+M5Q66n
xe/TyT3xN1WplLtrvshD+cItxr9q6pR4H0lRPVkhiQrsqxT0+APpEFPYBuhdu9zgi3pq3QctCI+2
WgtUG1vxqBGateQM6SbYiZhu1kQj+UpNTwJhnZXK94qBFg9+tlXxZLY+5/NmjS3xHmEHAgVoLK3v
V0ik8DwCyMw1oODpAmUh/Nr1saWiWnkE877wlxi2mKtaIAmgge4n+8WT7H0gOrE44AT+RkXhuk5z
Z7Nl0OmNiCjSuQCF+NtSkgEqFnTGZjQK4OD/eoxWqGPf9AIpNkqEF7/1WQvJi1ne22WTkpKUqn2Z
/kuQWvNJA7TSE/g4pRJiMbWyU6qEYf7EPG1dQkPPXzyKoEEb2bkp36+bYDhZ+DjVn23669rmvF2s
OXQ+5LpNQDE34QPkRLiUk+pAzGW7nmv3dcsDrnDcz+hFJwuUOT5l97WXGKG8r8rvfGws1hRRPuP4
B2NwKHnAc5Zt632aI6OKtAqm+X6Uw43OvS5hDX91cgmuaQKUWS4wriWw5pXFDflnKopGqE61BWpT
QPoZTlej29dpOzS65n8jhtySVRbs1TMLWOQvEPL/mAcgwQu93qV5i7jjgD1AqC+P4OCcgQ48Q1LB
0Q2BP3BLiUvJe7QGp2z6af9U4EjrZZM2M9tjBIxMedci9894hfqj5rHPKVF0FsO0uuyOCQg7KiwJ
qCwg6d9gyStVwqxr/xnnviLVm9TxmOoyYxcqSwNLQhZwLKzX4hcvf+CAR/4C9MlVOMzb4/ZkZmon
wkqv4rUMm4g7bdz6cSZfEp91dK+8LA7o9CQC0Td2LsI0Gd/oAjhyw7FyZIYcsuJY65Ogxq6L7/Qo
QBXYakPME1sKagjm6r5VLitKh0RLBC+YLvv5enaAKi4yjrEPQxQBCdibCFWBEV/xG1/PG2rlfrB6
QmIcSQ7nifb5VwZTRTJwtw14m8j70k7wYOXbTASnw35u7d4wuSQVPGm9vOQ91tSV9WuKJ6gM4clv
7GuMAdLCd35gStTraKsWA4PZqcheSSZdEh3/8vLLtZR2b40V+i2G1Je64dvmSbff7oj0UAy0p00V
xrfTDiyEh8lDdgUBYNRTL8LoFtq5IHuQet65P3a/+BdMNfIksL53PKuDpJuXXX4QCuRFqPgp9vhy
BANQk997UqR885HH/otUnOwsUSEpN0+2xXibNKh+r7eszuLaZmNehIsRK9pXwu8QtAMioJI/g0Y+
HM35RSH+biqNLvzjGK56ruR3nWc+tOYu6OluuLEPOSm30BcCeK/T5Dz+VNDNmVNFxjNdW3cG1IA5
f+KYPQ8f2uaXQTmwYf5u1Ast/vLUvUfII6m9D6cUygdGBIuqrKN37/KMud8eL+BSxfX8dZkgUkx+
c4NSmM+UTwsxZEvbrPw9I6oc0u/Zv08yT5ZAoBQWz9N7mQPrm2FqHx6f1LdvWr/D3p1uW5LhCcBF
gE057K2fClA1H3sTUtRotVu+KCqGMS4iRAUy3nQtgBFAczUGtU28hok2yph4o7V0F5aXPL6kMWju
AeTvzf1xzzY9qZK+CYmOtQVgkdGzpcHJfGrqHsjqdwgJ2UobrVJxTx85wm5kf/Dlguj99bAhnwD1
PLvNB2wDRRi07XRJ3ds71qCUZpVeWqCFFK14JxS/cziLTfwh5Tjq6QoMC4o7TKd6j9yTDZqdDuA9
aouz9eU/vGrBvuzvWPFpLNQVTt5z1EbO346iWZvz+Tig3WGdAmoq0fyLMvkyGEseFYfe8pGbKR2g
E264j6M+eG0uXTny6ZfwgTtJNUhIeuoDR4oQnv54EKOCSDyYA4C4VFjb4gNlMQ0BNo3aBaqJjL/7
hkdndC0UnlVS8hre5HlNcEy+VgtO3nR6IZG2tX00Ce19C9M5RJjnWTCgSmKUXr1xHa8Ro08Sk8Zz
VNeVUiLol3lseyWx1NJcSoET90Pi6UILgfxRLCr/rB9UDujP0zL+o0czu2k4Bbyi/4Vfl603vFR2
d+pDeQusjhP3oyu48cqhJhRAk+8hI+BBHvmxgevrXD/Zph3TuFZ7XbZHpE73jy91tsCY6u46MKvy
uRomXMQ90kTlRPF87YOqS1xn5dO3oX8ho0A8NSP/Jxcy1KKOhb29GkqVtfi6KxQoecc4tSFJmFLz
XNsHaHRn8meBxM4RPoZmje454LHxQ55TQQNcuJ9xmB1gX6zjFElf9dQSV1hbXbqtmsTsIKIJCzCq
6v6WXSYfcE/z4kb7DNDnyiVQhhyNwJ7U82caZzzEKE6MFO9O3apusUCbsy6QclnB3mCmJ30L/2jm
4uym1V+BoMpAeI41oGZWXkhCcCt4opIhCK6yjJm/c39rjl9vhsvamadW2HQLgYP7Z74rawS2uzYq
q8o4xypYaLcQJUyfkB09Y68y/jpjh3OD0+NUBL+iCsDGVIIVaw6C+wTuc6fp0AIUWJIjnfEJ3Y+C
iYH6fqHohrNDw+toHWWY5vYhuItcRBO2/ebaADv8ElJdMTvTsze6gqkVzLurBbjz8I1QTBQc/eqQ
67JAErJrc85k8cTLNGg+hX/toHJaAmxcYkue6IOuFsti0ffvrO0eiX1rFtB8iNxgs5to21gqTqej
s2W44sCzQq3pCLa4hO2kZdlOTs8AvWl6AzwqMJ0nLMpski6KA3Tn/Jd5mbiGC1asO0vEcIoTpMf6
7p4V0Eh4y9aYKGlMtrMFNJte077ut01UffXm1hIQ4RKTnWS9JJgFn7GKM19eMEWaiOMVvqV6+3Hk
G+/Ys0iq5KdpoIJymdmZZ3kymJXSAJO24VGPLSp1M22Hyr9SNUsa3iY8bu8rdfVqZlK61Z7095Ni
adfDWBMrfJq5uaBUrjP2hS7giZfUQUVReGvUPubpWgUcWuK5NALPU3c9J2e+pPa2m2TfZkemf0J8
inlnNqQJWg9tMBTC1y8Zt1ebpyK6GFx/A1Xojepwmhk0BG2Mu/ut6O9UDH2FIQPbVqDRrzhoOdfq
/23O/iI2GqT5VgcSzZBfGP1EULaI7cGzfYSorYVanePm6TtJa9tg8r9FGqPGZooaupiEN0pyLRgU
mouctm/o0/PD3CZQBF6Zf405Y7DECJ0Xt2qnAsoS4Aju9J6dmuXCF7T8iBA1GwENgdM+zUhqIMKk
mSjrJyvadDqCbhum8zpIk/WCdL8Lt28O5RzHztXm4F31FB2GPkM1Lb1NLJXM76ye0w04hsDoMX6e
s7qw0Wre4K0Qfdsy4hqyTAPQ90L/7kWuuJeg2zhsGAIajsrfhn4dy3s5CbbpvfSsyRkcIexc0CmI
08FbFckQAcum0l4R6tQcFG2+rGFjVM6ir/XLpnZ3VdjyjYy9/cQ/p8ph9mu0/Tp0O+/+6kPlaTYA
JN0EPXsiz9soqs9oJwGIjDPz0BZqP6uOg2OauCP120V74rwvqB0AM2qi5knHteyGTuMe9660IkSr
rlF7glr11oZcUxZev8pt6YYD85wziHv1mNRtgD6ygAu/TodLxbxfKu3pnkOyF1Bt62mOO4XVQHbU
OuqvL28YjgAIHGoRSzzHJhfa8SLA3swbYOE6rLs2FVGDzEy0FTFsNAtscRYUqYM7EHmcRPyrj8wd
j0sn/0sVj17RPZdCxy88BZKC9//hsczIiOI+sGvzBKvBFpcaNg5fp92/0IV7/OLbC1wIr6Fr9gPh
VNEVxuNznRtORVwXfOVbdfmjnpKmbsAoZlxPEnaUMp7zhbzS9d+pY96FRDzfunToOROLZN3pxdeX
6nd9u3mzKJ6bc9ekUw1BLM6xV+fQm6R6j78Ag5BMNWhT+PTp+5UMgkN4U8D6HOdKJLVDEtH41zkq
Owpo1tzFEY205ky9p/87I3BgTAJ8g6VJBHJLYlKijyOEU6NK5iaQB6sXZl/eFwPwyVQLBvyu+hR1
HiQoP49JdaaU2xmpzCpf5xHpkEiiUd1B3k+/2XVnE5smky/cSwyE/l9wkRHkoPNhsDZ7zgSc4ccY
+tfprMVixORJzOMpNneMToPYWWiJaf/k+UQMZvahELi8QS7x8EDJzfPshiZWh3Wnwn0n9JmSXlry
TEGCX/T4MKvVGOS1r0yEBy7dMQJ7uliuaKw2SFhQJlsXTUu2gmOZJ4wWPYZe4Td/QFO2oFnzr6mM
I483SHFn/imWEB7LrJvd4tUgrmaKwLRunhEe7SWa+RDhw8/3djHWa22u79mj8vKpzPdbFLFRIMxP
J96QUgmBYC8etEWFakCIyKZClidRPhU2dLfiBM+Wh6XJn3F+p+2zM4s+b0r6cVlJlDDfTvI7LH0Z
bRyLGTQtaF904/syQSrdfhG1hPkgtxlgzIUcz0m0SM5NlUjANHEJmDBydAcPCn3pMWbzs61Q6jEE
Z/PCbyUbj8+hy4qqk7MOjMMO9UuOvVmmvWUes777M9TtJX0+oJUC61sd6TlYglU52mSd39LBUs8S
edofLSF9lry4kBww0E2DiM49R/KS1Dl1Ydgm8kpRhRBnd6GjiZJ+O5WTk8Wsklq0fczMQX94bnil
M9EvWKD1Bkaq1IvEiNcxkLi1ADaoGB9Jbt0yn5qtKKdNGcCqCDoHIxKr3s7tG8TJmi7JVt1gIf5o
GK2IoLSpwuZiYUn6et6omObHgoqRtzxOw8gd/OeCIsIZ2nW4PzZiXq5ka7OGFiV6+xRxU+4g+HHT
M7/bJmY/rCREk4gQvMlCoW366xciWtzKU+kdjvCe4kIEhDjQBrcZ0ryVu5nPWmHMzfc8OQWs5KtB
SSaaSoCtQPLhhUw3v/fM1M4h71SgktKHJYoacO+feSk23CjYrXz0hqyS5wsa8CaxrRd3iHMs+MkY
oLrQU/aUdWAvo7MpwBRdVFVtLM8x5AOi1X3dIjRDA6QmS/ckAwxXqu3aWFvYD5qsnfVMZY6YlUmn
/u44m9f5skQEkt7pwnZkye96ymszJgXPkiDaP7di5CUH/u7s0uHymQ/wRsuwRfupd5gwDdkEJVOk
JZ6+PHUFthJrCVYC7heau4ftQvusjzS2zOZLxLuaKkqFpvzlhxlZ+THgZa1tuRWHtCuvUU7LXFSl
nbDiLYG0r6c5/nedLVnjZjv/ZVvHh7CBSNPRfYA7FTS5dkpFaZ4RMjUaNpKXIDZu2Lndtx83hmCp
bvKlATX7QpW7MGiM+5N63sKYHGIjxiECPZ+2NKo3Cpxre2Ams+ynuAlQifRtocdgzDB1jzMJ/DKa
x2KzxBBxc83mocv29EC+PUrWjXnZvn0RtNyI2lsFipWQ6etQjUgzBYsfSUcRAYvLHjau0x/acLp5
c09kuTy+z9CU3oCLiA106dxAbWgFcer/VGKWAxehVr66GOS1JxdkJsvlsowKUzut3RaB4X10T4uD
W/vVfZ+owRFrjJbGCFIwU51zYiturFgIj8OpFTinc4OaOrtJfKoSJ6cR3fqFOb7d1wx8NrP0ws2w
Tb3+8Fv5O8S3ves+qq7Jz5vcR2qjUwh/5VIpJ8N+UFKJbrFmIcPh7xH6esXGZaiMU46Z9PiUP/At
VVLPZEVXfhifUftEToTMbsy0nmpFzf9iq4nKxTUgpAsF2rEV+2ssA2KtW4I+SJtyjE0ZwbcYn44a
GR/mqjeTPR/Z2eOsqU9VWaJHE53IxGoGiullk050o/iduU2V/ndW23+NYiesKSEqYgFvxSYTWETp
2h/5A0jHhjWIZfpoRCkuPtDCrI5SXmnOCs3K1YXkcCEEEyDJsOyYIpZyAMoJoXbw3nDQzaVx+f4L
DgAkKa4w8pjmQna/uCutNgAvuECLUM7uE7aVpFtW82DshBYqhDR6gGJms/jgEMNu1p3Vp34iy8M3
PG+XLJO+fvIpXgqN3abFZAlXXC5XBQWELIoMTzR9tIstkv2YtsJ84iZpE0vfKO7ayfj4OzaPoyjw
aViuGt3ha8fZS/UEbGLZpmsZ/mqO1Njmz2T2IdbrSnvs3YNM1egdzS3HVIbQ89aen4NEaE/oJCre
+U+zPi1gzlYkdBKvg1cEG0dWZjABgdqLzv02SrR6u5Zdkw/dLovcMYA9Pm9dLqhQIfE+MCVSs8HS
Xu3gVY8YDS4h08KpuYnRMdG3HJzf7Aa7e8h+Ba4mPYoTKuEnmzsHHhPsSHnfFZtuw3vM6sCTFpWE
Y+lz9/RFy8zMarLfPe74EDpV9WQEjji4nHxfKczIuCLMoAvrrXBiiaeN6eD8q8dMlfvtiDsoWiV4
R6ATyrsPQaCwF7agKa6QcfnPfT6hXWI1X+K5IWCz+imUcsimKFZGYg0I31p39hlzSLuHnn/O+Pto
N4i2W1s8woFtaJgrzX8l6f51G7/DLqZRMCC8DqEOhwht0vwN6RGBamU7qFyQH990NtyI1GZ9bmfD
qD5n4FnasjwR0NXD9OhQus5oAga/ggMb61iWw8nCTMs0ABzFn46nWzYG7h0v82NRrFBXCGDlX07l
jVYK+okE8881glog6/40yq+EoNcFgy5O2k4zVyWTz3uLGlAmMHaHqqU/09URscdGXUL24E0PsA+9
YAVBjvL2TSxE6Aakd4sKluv8uhue5SdBs5DzKZV0rB6VC5LTi2edmqcEoNafI/bkizjZTfZojdIz
PAoqWkftx7nCirwjhPJkIO+wyLe53TjNaA5USC3CIttogVHVLxP2vcdBozBn4PA/UebYf/LmRRxF
Xi0ieuH5L5aWveUL5b67QxVUuMU1GDqUMYXnyLz53jaxfJw9fhpr+YiuJPggv+1Ijyes9kzjmQDz
z5jZLM2GfUTmHroDlq+zbdnM3w+XOioKJ41jgwONBYkihhzX7DCjW+CUv8cAPEVnBpim/E7+1iQo
0hXRa7EbjMWMRTrPpC5hSXM9AKU6x8qPgasukuf9WBapVZ+9OoKf/abrgM5hExWGzIbKQS1FpPMw
AHh1gmuVaSM4q1I/C3xawBycEotCDjP/r53RbLJOuHkesgi0sjpIDauXO46KBwWoQUB9YlWZ1w08
92ZgA7fzP8j9ZPrC2Jp7AQwoSFzuq6eMO8N6oth0BwEZHXFA55l5kIpAZY6gqzbxZaYZl/IR5aeS
9PLZPnNCMNFwAqcLUjesOybtYwkPPsAKFeW3YrGGMBxBw68pkYzoOwTPOnsUEnspiFTMFF43YZUc
4FS0NB7Wfc+R7IAYxvxqxFbgnZ/S6Cj0RD+os2Xr9wSVlAgm1ARlrvHRDuxXf9XirUiuUVBl1Dsw
wilC0yP9W0V0x8oG3LA3SaJVkJLrPcpJDXEQYnfozWbhdmnT7DRvvC9yVOZb1GGIybU2KKCvk+SG
S64sQoqmofdeVbnOmQfWDGcmlCXD4bK27HbCNLcguTFpO4qd+SSzAOEmajiAkrifo/IGYbe1/v0A
d96YDOKKg020yFv9R4VOw6RqoDNRUaC7qwBxgS4QfGihSrCdGRDXQZeI9ZHmDEplf9STD/1RlcKN
zECiVIAS2LRw838nj3krr3uRldq+0TVqYgtoPY4kFfgmtdfr6q+NVBttSQvI0kEWL7dDRHS28Sow
OvloaRjvM508vrgpCcRPzeMMnnuz6vXp+Upcjyyo5Ep6RrD5XGB+NdxDsEKmxwsi0ndfYyppWc2r
75Q5IexlSgXG97ZNiOhDQO1rKXbW5QyS5zDVF8jMwXvoTTGrKdhqp8x8XihQ0H1Stv1A+VBrAKcv
An8eAdvRRj9oNLigyEjx2ZYuv+SBvMBGRfw+zpQ5YjOZArPApZcOzhr8BmMSVGbQZaj+eJkfk5LJ
gvWIwBy6SlvgB3z+P0EJ9dGrNjkXtENDWgCE6n3f++pUYaKRpG+klORRqOWwC8jGYZhEf3mnLCsk
vr7aclDunmsZSWPy1XpN8sSW0T0pTq+ZrxR7u62NZI+PvHgQenPmsaAKk/BU4TvZvu7Z11NXOnxq
04hyryfS849J7mZu0796RKqVdH91tYQx2lFZTPBLIydyhVKN465t47Aqhpq74sg1mEy6n4f5sxxW
4UFkseCvocXSYIvWSTUo+tM4Ft4ykgYKI9ohYr7XIaXPHKqgVt2r+f7arepQZQRToaLuCTLpos0o
b4Ui5B9RH1smMhX5EeynmhFn/vdpunwNjvMn3Ue5dFUafXweu0+rh8KbGDILXTL78g2dPkeFJWFB
Pxv4KFDdwWL1Y+fZDKjqKr8htUn/tFIxEqoGWFDZlVajAO+gAgGylhNveIqTwxnYQK2aI5lIU0+G
mXjLA9CZLKeTCRfnplmRN3+vrXZ65mBX2+uCAzxqQe9jPPJoXqG2y5yO5PRpQvD948okVMhXhoCl
KjCRQbJcqxdXBb4cW4p7GaVcc5J2l/ffd0qNpvVU1TjIfm8MUStaVLtx0MKOUoGzuSZAZXh8ZmYJ
340lS7+3hqjIR8As7zK6sbip2flu33sCjJiI7msDh8QYww5j2hXdwrK44lVuBSBw4VzTUxPqFiUk
ZxDezvwC/IWU6OMf2iMmuVFUBBOEaTpy8e4VFwYFiIUmq9CYF8fp8gcbfFo+yvEBKzkVIDYaBeuY
jU50ArY+WbK7Fu6jC6YMyq00jl8imoqCqcwVdGEYl82+6XYHAH6GNnfd3A7UG6YdaUFVm927uvX3
R/u59LpeTHyjyL5l41YnE/HsW/eqt1WuCbbRqkeqvS9XLSHRTaV0RABUjLlV+DtxNCvBfmV2XXRV
NMKDMroRyXipDRs+uJQoWI9YkU1x1oSsB4zRwti1/Vym75C6xWlNmh7FRWjzOwAQ1ag5El4GXLq/
DdxiQv1hsElmfDVjgaPgaThgm6gSXguNMgvYPDA9BVGDMyACiRBj9iqBfCtfrbUJRy+rA55HYELG
YF1SH7yG8HSf+XmHB0vbtEMXSR1glFvObyDN/bk4l17Xl3Iba99jHE2OxK3/Bt+93E1nqXYYhnv6
gQMNQg6MkZUWhy+2/1gJ+vRoGRVt9/VkhvhPubt2KtXws76X2sLP8cSIF39r7OZN7cW/nC5uTmun
pfnULex8uE6bglyTVsCZ8MmSBSRvPtR0RDyTutiC0lv8H1IFwcnbu24gpLBL++tIGcT/oR229wtj
a1njUsIEbY3FIR0th5LMpDxrLSg2y/ACb3I2w9ZJ+MYuAwGaPO59JSjA6HUsi5bSYQkTVf+mcxFq
lJkHaqR5jq9oPevMqsnhOWSqRoeY4l5rbmEK+/E0anQj9oDw8QZ6HI7alOLlTAAb6ytl4p57XDlf
t8d+xComXJRr5Uce3+ML/7IRCKV0P2dGxpLw+kx7Nqs6xQ1moLu0lGVn1czN2A74nNj96rJyhEsl
7AGCZlfJZ/NGdqMthlSnDh2uGaQHfWEI5Ps8TTyOlN8CD4dbT2aNjJXxQwQCKXT/jqXhxB4F6BpQ
flqrFMDRzcT5V/rwEK9H3KgXYXD9Wlktgelw0VnWfCcV9ytIze3vj1irzgT0/anxdRAzHBxcHUJq
K4IPEzrGppj02rNT3KLZooTN1k2PB73wqsOJ1vlRx9d/b6/F/Ma0NB3kd8IciQyBOjSiskX1irOD
dtS7NKosiMqKWzm3F5h9Jlej7hddsk2Um1MlN2jOfCetxnF9BE2dXFnTQGig+Sp7Di8okCxvS8/L
lc+qsMUj2bdMqbIQ0azyed+hdVlt2oksTU6EH3X/MfbST80WE5Nj2jdxRdMckpYGI/QrGMUm7WC7
uhoNHgOhB5uZjfySyUaVB7k4k3hr7nBn4a5C+p24ash1d+43ROcZkN+wzkdFLYRDaHZ4nujcew0l
e2p36/kADee9XkEUKsypcG9NzWKLsWQdDULeD22cVCPTqrKLrORtP2fTK7Ulm0Vw4jn45lUm/LoW
YY5XpxoWV6TyjDXKMJ49Hu0gWjVlJVfegsNMtu8IXErSDm03ukEj+ID9z7k1mm7w4hacVsm8NPUk
/Gv6tXdFDaDUn/1Yoy/EZrpECpuzFZ0t82aQvposQCSF+80WwjwOp8/t6D4wIqscAhJi/Ii1j3nL
8VNRM4rH5d62Yfdq7kfdahBv5zPgxgC2Ak99QR5R6eLAyqDD1BShG9ETDs9c1NHgZ7ac0R31mKUU
cyTa07gEnzlOoCHagtjGRrsqmcfJv1S9SOxYYxDFSn0RMgbYQ9SZU35Pb1nxpOlEEFY0dI5oWOFr
9w0Zmu8gmvepm9MZGfH1r1N/RlwWGIrwouk2LmOSwrYYqkY0FwkUciyF2iiA/k7YLilJ3ctug9CE
ExBcl0Jwfp0ybhjIt7s77W3TW8IyL3aoGVSYXNU73ceV10H4E/VDn0I3h+2SSsxz0/VQLQ4ehtJ3
JrBwJGMOsTZIQiBjkg5eMs8WQ708qUuaZ5SaqrKYbVOvmONPlC+ClIa6SPmmFmtDQHBJPWQQTwWL
vHTc/oObquCXewaSBgmiXAuuwad72dRsk2wRwkKV3NNE53tBdIDf45KHzWdGWdhAthXTOePZG2uX
8WHe9wz3bhaj9UxCWdRbmKfkUlfxpKGQlgVBN4zqcoqq7zpyHflx0UQRR0axb86VNrPlWvX9GVUB
QExAP2V1eGFbsjhnYpwak8VWDqnj0h1zxzXmpPFA4TYK87g7OUZzzN9LQY5FjNHEtIThibh/ehH1
pKHERfC4Nj5fiakCUy9KGaOCyzuEuw1B0Pcrtdnd5QSwqpvl1cwaaGqDlqXUkntEYuSL0RFAFo+D
cJi1ifHrpu0YpimrPf24rRQAzwSc45yqQleEJrtQYsvdvulnbF/MKY/5gRHHwo8af1zTjY+dFfVL
4O8v0U6OkD8uJK5C47p964nhZLtmMHhw3yhdgIQkvKz1/yybvWpV2yK+1SnZpxRuYunS7nuzt5c6
ItP6z0zBlu053S0PJPE+Kc0IDxQWK6RRdFiCzNY0oP2UemxsL3Xo2xdBzNFh2JhWyBd8S8f+uVVm
Y/ZZVr+9Ih2QwHo4SyfbWrNXVKzI/kUHHlV2Ba0YmfNK+ngj2wVI3HjVgf5LYvWTerxO24GPUz9b
w0fiTOsZDT/xKmJOetGT9HA/TF6SXsGPABZ/RO65rxwRNcg1mzus0TuImhxEqdMpUQXWE1Y6qV/l
rZ/DznT+HLchvXKMZUNs3zGpjeEbS8id+eRa+bzdYuRnXlRRou+Cxvl0azwcC2ox+ZcuCxAmYSW3
d4hWhrIha/9D1UBqKfSPQ3IPh8Kx7mK9rF5ZS4Jbny9toiL8vXA4MDu6faPuc68lxhrn7k9FOjiJ
E9s/yCDcjwlath/Hp0IQAT2pyYedy56WF8evLijdQhdGPpT4a1OLkDSmyEeMq7glbmoLamnaeeHs
fH1eyytcjl3+QewoEznsFEg6l5raYKvGE9OUprXBlXHexaq8Mf868bfwC82pH/hr9AL41DXntQFA
gnyq1RVdJmTG4xRV06EF0r+cpzGxqwwdUY0mztxw49wXtj7tYE/+1lTB/a+jf2LZKHeHAKgVjMGl
sWao5Q4VzPEMt19D6bGjqPXshkGezYnfV/h8pUNY/OwMy7fBDGeCq8A1KDTnExb4AEX0ImsnBUwq
mgzdgvNIQM8JKrCUata3EGjkPiPp9zi9OZupUjwpHJXUeD0lIfeW0tpmmJIHp382Pj5fMFVlgBS6
i69eug9RNvYScD3jE0K+kBV1i+o/tjjntLzP2o06Mk01hhHx/fQMNQb6rN6TAQUsuVVz9gssj3pf
soBg85wwY36TzPHsweNuzF7i/p/nFBFRBORbtBn1pcF/yD6Mfcv10ci++CqBr5D8zXh8ENoTdmR6
Koc5Zjnj8j3AKcz02MpTeJnl6o7Gl7DUux7UgC4tS/IX7bz6NC+cJzMy4Rh1Q8t7h7kuY0ULf693
EfqdPMo+yFqDkyutO2DvG2x5GQDBBve4HX5E0aUW5N+i5swLmo3dt2xE2DUlup8+DEqHZFPJCgy5
KOXmUNNpfVkYjrVkHKu1oxPJ0ADFLvF8/DpDDHbOAvu4RMDlVvY9cG3Ln8e30mx9K5zPN5fRDnAq
u4RVmFVnoadQyyiRITTebFSLXDQYu7FuzrkXmM9PQEDXoRw40TjIwj6Z7Ov9MG0BUUEN6BOcHaAF
NHOMCWjvrGc60aYeq5BHG9MXRmBAILfvRZ397t/uOJYBtkhuaV7BfLxDtJFvTU9dtNs+1zd2Bi6P
gIt3dXVrqcLvy5onK+mlaNzKcdYKwKa1QtV4nc0zwj+zLqCdgDmPjSumJ1cHXMR6bqRdjC42pHha
PHTsUWoJTvi086GBd4MnQ/6FKckO3t3f8S4S9eLZyG2WWhqvTKvO/nKqCuhPSClCDP7b2Kc5CC4/
gPeqeulCxZ2vj/VzNIsWt43llT9fv1EHyiMpKJ2ADbyxOLAJGhF7HDxgwMFo59H4aSTitXHsSSar
0BUOJaocP6miE0A3Fek2LnEJiq9M3ii/5PFejwk0/a0TpTufHeU9qEqLVlPyGN+D+KKfB8/6y5W/
3e2SNa2TTINNyGXfPHJOcphL+Nc/AAkJ5paZk9t6+qzrYqH/18OKywTPysjWIRLGNnsWJiegKgNL
EIsKWlhr7sr23uZjakOuVUVOepg9CJtubiC/+Jhs9WBLSf+7+xGgI/UIuzvEIOTkXWTTmFIqWAUX
GcbXa6Mzrtheyh6iLk5Kvo6+ZF7hpdo9s3RHbq07aGW945BgBmrQCPwRpk+cStSkdxSldbxHhtW3
w3fCMlIZ0EMKVNJ1WmEtQkRViH0JJyGTHdhluIkaxuhpZV+MydVwHB1802+wtipJJEH942xjnexG
3M3qoU9hMp90hBfx1Zpj+dFidcPl7Th1IxkCsJ1AB9rERuvxAGq+ULO8Hx0bH8XhoN4n/GSn9h+8
5oPwgkTLyymCiqsrcwudjGzajFInR/WwMksiNr9lKCvcfchWh03ov/4HGIKf7Xl3FyGXnWnfdYxM
Hmy//1YSVO6LO2j9kt1yovsei2ckFlR9R5V0tF1fqJAOE4oOVINo50Z8ImireGIlAFCfiigfJVHZ
oYyWjtOrq86QWNqkaEVS9IX3QmfDXSChw7ktkhkRxivEoPPJYC/n+f/ntahHBLNTA7qz3YxQHKat
DKcEulAGzc7nI4NttMlyH1ZsTtpqj5JN1yUYXO02Mu9Wx05K8sDh/XR63Fp1uw9b3WXLTncfAuqt
fV7FyGtQpekWC/B5RElNd4ilPk8JY4Y1dMEhPbaUoaQut3aDm+Bgik3gToG8I/fltgrV7Fd9myoH
d4QoU4grgPUrM89tvCciQrV8lfJqBgOHqdtc5P+cBKk/eIucYwDjIufmytD4ZcPtMGjDDuMqzRfT
RyZpNhryvH3Sk9Jlen7zNM28AoPML4NyylBPUoIvZrILOHtSEt4oVlACuzjxzp7YCHmek/XcC+RY
PsxgOrQHWIDP+DNsfTmk8XEWXfOjgBtR1nnuJXG4nEOZH9TdX9rKwK+SYkvsI6vsehnHHanL7tsk
kLgMgZvlcOXolv80+qO0adNPirEU//hYgH7beJYeBDMh6CK9uPEwTMWVVtb0WeE474o/eYcPAtEf
d6p79RYPdGJSNEj8Tmbj4DDtqevQUjiVJ7VMctU8D5LCRi+0yQfmXkD4oTl37Y7vyjlKvKiWIGqd
kAAxLMFAQVmdTKGIZb8wDxpUkc9fBsyp/Ujn8FLqDzh/uHmbLHCkGe6Lwp7yCgEhQyZ4PWgvxCXL
zp8aCp0F9//JoOCBiVxuC7J7b1/jR4+eqlA7IaFtVPLwz5gP502hjkk8yWg28JIR7PYGSRAre/eq
LnXEhnaXxh51QNqpsydoki7QTC5+GcAihFsIGHBhFaNmjEnWF//N2gG3Dj8mhWuNgzj+kRk9Y3ph
gVynfm70R6Z6+QHen7MQVOOf9BQjmYzq65yNeZmadEEhxKPfPx87tGF0tNnFWjzxJmCJPHQ4ypF3
36vhuiS7tuGdkff3KtSDGfOZoz6/SMta5mZrpSk/0mnB/BWl5vX5dVPUve9DDOttp0qUk403/4HA
TSF3ya3smLGVGtjsnU3KbX5cCe35cMWv1kn19Oeg7qQVv+cVRQtFdRXpUnwVqkIwQG9paxh0IkUU
Co7ebV5jE1GKoGojOCcRDkRJH0sCfh3I6RMZKl6CTjgdYWHPuDfrYSnnsGLuRvMbZqXvsUQnZzzG
aUrSK0FrXqEXtcxh7xtzrYjdC3No7dM78nRtGPpns5+nY0gJnaAbQC4U39UyYUB/fUiPnUTMCp1t
6EiVGjfxVVqysk+YzB0A0CF9THr8YqRwH9hXuqDrOr/+a9PxZG8W2Q622ntnrmOYGkxn1USerHcY
k/OgHJ+iibGidBW1wap2792h7OYp/cxbLbUg10q6Aol3Zvt7NcJrh/RL3QC3bCEYGSnYKfoJwios
rBG7T7vnJ8Jqx3VoHwzcG/DCcanimNOtlbwECzjkAGZovcefn+V/+z/rdP35vbcRn3t+561wbkjj
3reA5w5sjA77N2vQTT5z8wcTzgXd9Z4oOhLIlypx5NhyhhAfTeIcKQUcjXJbUCCUtfe2Beyf/P4+
LNRd2XQhzm2s4CwjlfKdtgnsRsOJJTHS9Y2CHs8Q3EXVQ+dbUNzy2Wo9EAoZHt3U0ivApxlvHN8t
N0/fGtv7qbEdC8hQJq73d5uqTvkNruAptUTg2diZ848M2iBo2oltccWnj4KYdHmeMT+/rDqXnbRF
4seexu4HKuhGjNaZgiSJqjp5o0s/qN401ajUPKrSX+BxdIza1TTNEqIrCbQFHAtupVNmglWc1dL9
YpbiNK9tT3VPoDhnEimszQBE22I14rMHp3holSdDsoLT26mBDtMChPl+xgVxioJ6MFZ5p4GiiYGp
rftiOkBkiYf4GYVkjfRCdzferd/IC76pEL+1/ijUEDmF0e8GaNT9yQA3qpbavKx1TYjPwwrmyo6u
n4Kp414mZHfH1OUF4pAN0Ci+37yxgYkHQfhiEJHlo35APtkggdil1LPOlwLmeOBp0fPZTA2Fcg9f
skOG8MxBzxWGUqKybiIUHC6GP1/ElnJa/KJ4+zp/D9id0PH4E+6GXkMdENoK3PugQFqtR7OBlXLB
o4Ckllz8r3mEXJgDmVIsduEMAXPnYahBPw03SPFB/T1b9bYjVnfChcP1P4xkXylBKRVYyA4JlxPG
Dn7B/Nckj8fjRyJlIWssTR5V9cVXJHNp3+pF530bIn3QsJqsNCXVJWE18gBtDze+O2ZEzYGKe/pP
W0F0Gx5glJWLViKzNJebwz7hXyS+LdmquiXT0sdsAcjnAS86SBhEDW5Kb7ZUnNcF85mDy7EJRfKN
Ynp1uYzygUAl2FiXZA8UX/TJWEYvFGvsIdWwcGwPKLUzZJt12UglQRFK8ZtmSKlHAiNxskWxe4EP
Od0bDvcfcU3xtjQYttGIlxt5Ml6jiHClhZBL6HutEocA5n90t/DqLVNieQfeRAnvWzYvAv592ZDT
CkBNCJi1sTjmwjWlKMN9y9hx/wyFiqY/F8h/68Mi9kNNY8M7A95i/97WTBBB1Vg4QAVAdE3QxJVO
9jsxfBw0Gus1PbBVl8zgTxNI1+DkiKCrx43euo4ymUyNuEUgggHfo18E8yOaSQAURdClLFsb64iU
SVZ6iRMH0sR5edcgP3FPMewgVhWOlwWWomyFe5ElWiiLjjMOJPzDKsXecRkL8iR/wgxqDCF8MKct
rP5KWc8AnLF6nNKv3ft1cLYto8chP2n22nYGHVPMnoc1HPKn+MVLItqNAqx/UAcGV6/b+Mo20GCF
16kqI+cfdb4oyjn95XnYHt0mjC4341T85ecB5fTREk7s0+V8KwK+LEVKpByBDDQtDtdgqvOTcdYQ
McAU2zNtECU0fOHXTaBg6u2JuFlejhiBZCtMUDOZwpjdofDylsh/91Uq1+SVY6h3Lhb2cyBJD1UT
nT4yKE9qVCEayae5MoupG3x+KSkbUAEdFA6Hn3O/CqK8QkDa4TWqB/zVjj2GZCNnOeNBiQRnT3t9
eypLJ0k8I11jnonG74vSYLSWv2j/Z2/apLiCOPOGL8YllKAXOGthBQfdofuJwgN6vSXHmlQnGemy
On7fVVXQLQySTIqJaCEZMr6MmcvDw8766o5YN9RasGMTwD1cuUnTBim1wWmxJXiTP+42ca5cw04U
+NWB3jStTib1mmfSDqREGkZdL3cuDSX/N74OpFAEHDGhmKU8HGbJX2D5MArQzxermSLuw2SlNxat
1oJqQ1kfQkFJeN0SqbHR+6Lln24glUbudJCcMgp0lLxBDLcxB796JIWlCp0LJeDPXG/GXqU9YCQG
wPHcDPOkxZySndjGdEFsZ/a5KaWorn1MEln1LBxqBsEYqawyPxdK8GEORWLmxYKSYCe0KfhSucr7
gjk10uSOZ/4ZnY8P6jG5Ux6Ycz+WfpFSFFuQ5a9i4xHiwZsno97f2SZObqq6/q2r4vt3RZfd0EgW
W+wOrjpyrgaXrjrlJYiOiAXhZBSOV3lzJbl246GpwBGPDQfzEMudwC7u6EK91Q6QfMmthzPXXooN
xxwX6Ljs0h+RAVpKJa4X71yNNt58uYJ+7g90St18r5XMVjPPhVkf/1EdDwV+gA3jRDKSIrvWcxk/
yfu5fHUqD4RObrFIEN48ioCITIosqQ2fA7A9IJY7T+yHBI7RirIdm/fyrI3eBBfnCFsBdXoF+h4z
oDbIPHWhr2Ir5fZVc6bXQSCS629zvG31bqcob6NBbRXpO6JBwsSPAJ5zFqrWglBXWhBGtncE369q
2uqd6tuUHz+6KJEyNKctHbOyF+CW7T+0A5NpmPQLkSpQuB9pWVfbkzfMFnTyqIHK+dj3hnY4aY9p
eA/2pts6T2aDXhqicNXiiHG9st/N4Sk4Hkxa8pZMN45YN4CYg1CclelwVQKD670dVJUXXwdujlLc
nffDTxANxdswuuKDggYLfJcm+cF69v2W3Wd5qYjHNElCfQtlzrQzqSUjpGRib4QbFjU1I0teO0LB
rQab/dIiR69D2jcEfGkbV8mlJ3q6X5Wxq8YQXEWV00ZvreOfVccYt4ScOZczVl/oRDMU/GZs52or
e2T90MgKnS7UHX39YH0eVPGyuFW7ASTNwH9jU3J2VMe7r0UCMFI/ATlppSb/Js3yyGVsnqVGJWS+
QKsYGzoHmEHb9KBKQO1lhjNIajp3dG5jVlVHNpSWXyBJ1Ya/dM6kMk8kdzcvoQgLy6MFfKLaLXiT
Gvb/It7uYkUzZWWREy6iHvwHvk5ix97A7LefjlpAZSwjPKHUcNRAA1n8zfbbNjaqXxO40nrZE/wN
7qSvlmlnXBtZ75mrSnVVL/OLzW1VxGhf0WF5n3Hk6qEp0+wh31cbiM88CZ3P8DliTcHlFkOTYW+E
9rkQmWAcee8lyfA4j9JlNO/XL57gQUF5ghbe138COWMjNND7ctFyR0W++gnIWvqVCtxjWSEcvZ+o
3sSyGjpnmv/GiIVrjbd04AzVH5n8UgwSWHC7uUNGfAPYOrkboe4+evCOoohPLWnmmgOCVyOG7/dy
ApACLd1KbCmOvToJSc+0wcq2cbCg5iBOTN0wTjOnG/Odvdfe0SsO2eJKxdvoV9fMSuRIvPrFNEEu
1JbiSF+YRbzu0EJeM6cc3Kx3jTVgXZMLu++1TpSo2p7z7l4U9tANYaqB8mJ7k8Glwhlc47JJi/ys
/dl9eDs2s/H+kps7IlEF2DT3ScseADHyyzBXJuB66O8ITV1zAgVZEfAfUdnRG/mFG/irsEt+VTue
FrutufdsgFjkiQSGun4GH9XBYLtWGRFC/SQdjOQunXYBKs0zuZNwEIyloeOEwAOkmOV/6LQWjyDl
5kQBZiyhK1MAWlWsWg7f93sB+IoExKhBb6eDJ3t0495B180FMUBkpzzegXLe2PzEJjpoCr7nDrxl
Y39gHLQN8HoYJSmow0msT0IG6Vs+2NihX9bz/P7QKuSZ7zGuWOQNn0ZV4MJFNE/wDPezAupjgfCF
QlJG9zfiwPUPLQZQhOx4F5B6CyH5+mJ9SUUYtYjDVgu506El3fNyJzGrfz6LmuZR5ULFi9EKIZu6
UF6gqcA2ahlSg06vhqO+ouFFWNysNRv3dsUyga6lq7dwhVitURGRcn+DElErp9ftaAAPaWaL0bXy
PFNE/ucbcCS6D9CdmM56wLGGgw5B+OsAkB4CfqIg4P3VosU0act8iMJCVzWfFeR3t8eKS21Ksj0R
jcfqsZtgG4sMt76Mw3NILrN74WzRawYwP2qeabPVFbh66/nohmP5nBNgw9TAaAQVQeEryB9nxACt
JDkq0xRCiGXC7K2ULVd8I0XuxgEbLCwhc2k77Kdp+Dh7vInwNI2sJE9/Zy5WMBrVifDkUSfgL9X4
hayrQXfGfi6fUjlS7DuA0WYGUUR0Fx1jgx14fcrumTdCeZN2lat9JFLlusLRVe3XeNBc/jmwYnAa
ihqaHZiFQgAoWgV7b2Z9xOyAbbTHsUw7Mr917Q79IkUXRviFVBSVuPWsagg81MJgt9GTrHrkrL4Q
nTom397y2ZVY9okNCmmdskUAthx2N/fLuTd3WR2rMmyNF5BdnPHFH32bF5oW1+701EjcBliY/eIz
XNR+TNL8cVlyJ6N2RQjeW1E1wt/LPKLd2bWxx83O4txLh+gamarFwiR2+f8L2JOB2Kg5z/3B5Oke
I9A5G3fo3X8DGwL4ur0lyJT4xXyvrvS9cmuiTkZNKyJWPOzvTBPhNRThdKfj9j0mLao367O5IiJu
g992ZkiOS25n8qzYnmbXLxl7TwUZXWFngN12BKfprh5w3PR5VQEJCHLJBj8wsZcXLcY5Tv74Mcbu
2Oi6f7RGvql5p8CPm/lIYr1HZwkutjRj8de+dzpmMPs3DXUoKax+uQif0KdlnmxmrYa3gCOvyzci
MmYNIMNVnS3M9kFFbJS5D1RWkgW5ZeIspgQzA3pSHSUprEVufNpQc5IN0FC+GmXqzMdlW/vnhlkT
/iSxE00eW9uYyQM4J0xrELsRKm7UiPGULi5oJm4l1SiiQdPaBqZmrg831ET6xrTKUz58tYTp8tby
4Cm9zcs5AF3/R96Ei05A/zDgWWMf6OosEigpS2KBorUVNE4ODpYluNCKXKBwiYLH/O5rGLXCFcV5
k4AG13nppL4aAudiDsO8YG989EZsSuqY8UeosSyHPLVFQIYc5cp264sGNranwPiRrOKWiOq+1RIr
RC6i7kPwAOb2J7lyCyKgA3IEMrVPTlX6AF//6slpcsAhHmK5EXHKzJd2z3+lAfOWzpJo7G71/siA
Uv9oI5BAirVN2pAR2QUln/uk0bJMWL4Cyg1OtbcZX7Nhw0+cGble6Rb6epFg531vq4cUTsQVZa34
h63bRbM/dCjdq9hKnJhdK4f5jys8UBTSR32fkLdTuJkKdz1hQhhUgkYFZpxfycQ5ZEomO3CREF9Z
+C67RJjQSLqEL7wrTZTXDBxynj1D0IqARKTgHk39z33vss8jDehmOfSPMgQ/6qAog0CI63OGU04K
EZo/M+PVDUEaKnclPDQ7AZR0DtBcpMJqtmRBYwc5GCiIehenWHSWTQDG22+VbytfVcFgiLb23FUX
w5SJ9R86OWUAIOi9P6nuEI+lVLfnLX7nPkXgZvNpguKVqi7pdiVA/fc6iGQdJ7IguKlXbMYzsjAj
55ze0Xwx1Zg4+4RP3vsiuqTD4c9GubVqBVzwTWlCNaLsOrUQYU4YWaIn7KWt+cRXtkl/We54330m
WCqWKMdoLoFCiCDek4m6XCMEmQPj0mVO5fbivL2RB5T8ZZXKV4TDG4L6/J4dAYp5AS2PM/N220tB
dJFRTENNPw2nKSapWY581un72Wr/RT3QN3LvEuv5Ozb2NmTZyy+hhxwQDLbMx19XuQ3tSvBt/4Re
rDhItsNmOtKV4AFUJCp7Om0QSG3DBtf/EyuIo5FALuzOxkLOS0kMFcrGLtbW3da1xNqPJrNufoOA
5oSWfYoAuOXAE5rxsHqKCOYVKsjS1rTlzs3OFqD8sfNxwqvnr9iI++OgCJ+dlSm0DlrZirU5j9u1
iaJhrDA/uRee6cZ34xRVrlUC/lcvh3vP5tpQu/QJB8RBzhDGdEofmfPFdX2Zo2Rrq+/2LceVJ6xr
VwRueM6w+Ob+zrVvscx6EwiZ0dduVfPX2PWOnJHPl0YVheFdgWWm6zcqCrZU9U2HgjKxwuxMG+Oh
XH+XRp7Vy1FWEqZ5N7V8wcd/bpLDy/0p63JRI9hRXKxtE4Qs0BOu2s3/Z5F9b2XvK0yrnv9w9rtV
tLp672zqiuGTxCiNWL5+C8Eu3IKBtwuG6ez+SFc7htoG7liLG0JAJLn49Kd8dZER41fR2Pw42kJ/
wrY92Tb4dogDmIPi4Pg5SbOOJw4sy2zHjw+i6R8PnP9LTUxeWPCJ2EvmD4RhS8Aoaz6Ict+dk7lw
ERvVRMif/+O5y4/5r3OSIX8WoxdsFN+ax3kDvl2azo3GA0Gddfu5VwB00bpCQ5ZdbHu71O17oaW7
u5wIlwfjfpNz6YT37YcvlnDTenDm/jr7QlVwSgk2J0Y6oTmB0d2/c9nl3zpWAOg4hTTktXBbHYb3
r/Yv72jR+HNTkntPU7nRUwB6HZGU9ONucBp813dUOTm5/W36LXp0nyFg4DPosh7oMocGmqdPTLeq
oQJJXHArfAoNoCFF4zbnCM6qfkEW2MmueyHU6iW9DpbSsAq5aL6F0vTkKuVKYuHWFjBSzj5S8WVb
KXLtFii36r5iC5q/hYuwy6aHCzNMLzV+CngdbBalDc2bo55YyykQoFMsi/uDRu9+OgHETb/CIe0/
0WBQPhIKbNJGc3IFCWf5cqSLzZ4S6+Fb9M1suEpNX2Ro8Rjj8WQbsN10Zk2MdmuHwYcEhfwaZB4E
60LXMYMEDFtlyjeH2SX6jKlwiX7zD24mr0t17RB8AesmscBot6uH4t8muBikSvbyPulDULy32gSO
MkuwZNQ36lmZt7BgeYiLZP0sd7VXUE/V2m+be8eqpmK4wVaklGrNTS58HOI9W80GiHW9RaK8nuNH
FZTXY6UUWWlA1s1VyB2ug3i7w939DB5n7+JGFd8X1LtzW9DZ151fg+b7ykR4Hb5g2U7noj6KaI5e
oVnzGzojBg7EK2d2U3qzF4skiuFM6sIfr2Tkk4GwkcSFtkVJ9kacKyoCHBQb0R0cjTlymsHsnONJ
4PcXBkfwWLRB8kHjCSJzg8cZxWzbVAGCijBNfLRA+FhOr9B8EVuL8s+EuaKNyTtlBxYBcVYSJ+1B
HO8c622fJFJQgHVLpuWuDZfInHk84KYAJAwMToVxninJamweDa80aVn2A7IPrYRk8cdVzQqxmu5y
hgFYp2KtBGt2cHidHMOmtjCGkZr1/RMxN9hNDPT+10ZWquWBdMhDJXpC833PjGDdjaWwENSWqNyC
1PiPiwgWquCqQT9VvgqPTUCZHjSS6GLH2TKB/a5Q68fII9/kG0aVPLTmWDVeH8cJezP7D/YkFXsG
159Jdxu0LrFVeB7GOq4LyOTjPQFBEs3Cgaq9bR8gSjVAObp/q6UBROi1az9KrBxCmJzIPG1+aiW7
NN6VVALZyzWTZfhmw+OfJW0u2Twq0O1gDeEUJyNRP/56EHZge3GD/atj7c20bk6KiIWqYXv3ecNj
d3AI3+er7d+KFpQy6yF5nM4/3Mro6UQT0rdpfYKZ5wPiNb3nYv08Yd4VGok0Zs3VAt/MlLyykNLI
CCDugvRyMs6YZdTbnH9kQJ+fl093oXyfsaljl+qVvBIfEeCIXiVYrkZYnkzySO+5DklmfULArJ6k
FohPCvbl6ZojtMqHhtbFjraKLm2hkDz0n1HL06k/9rJL4AHBd3iF1TaXxO+HQG6scuNXRJtKU/KQ
D7JCZy0Azqh3igAP4ycmjHn/T10rEEhhABvaW/V0yCY29VFiK8oush3Y5cRQ23sxkYYTPBmd8RLU
zxDyn9FmqqUioSrNBRCqVJ5SYG4LdmLeHiUpfKQfVbPHcsWUsWIbaG25x81Jm8+bsTgI2KH+6qVg
YlC/4CgsZmpY25d/clyzbUm++tgcdYeC1bLToK48x0StwzvxqNs903PDWQUeMABk965W6mSbDnpv
awZQTEfgYDvdpR4m2ICe49NUvxRxfqEZg12ecwXiimpPNwh7jSReP894neUDgxCZ4bX656KLdQhj
RNHt7Hn5TgplRmfRFndnn3HX2cCa9BvOuA5XomLdiBcgkvuYQtEYnjYooZSa9qmVA9F/aIVNf35B
3J6MU+WPrn1H3BDsRMBDunm1drnojmki7+UEkw+K+xdXoXOCR39QSdc39uL+6eEIWCagCUFHhj6a
8gxMqGvFRNHsGuY9zyo4I8Zb02XZyct3HwgigQJkRYvlRYsMrErCwliwmzdoKlvea100yGAKjEmC
2BHNFYm8fJXQKZ4NWO87oZp27ayTjwJw4Y2FtjlBf/nb8uy5rVwPd7G8987f7F0wWUb6yopyP7wh
jgsBcocld7WAy+BvUzWEfOveTHmuShDGHJJcq6k+C8v7lqs5Jd10S23OwQf0SKH0NSZxyvm3xHyl
8FyC6opvDdxk1sgq6OE7VvXYWNR1vTBFqr3LQqOhD+nKuIeqz74VimG5jOyEboCZcllzmzdabiRx
f63I9MRzVVMDufgyZC/9RnbQWRzP++3n1o5szoyoKVs7FrocgojTuVn/XcT2LrYXACQTGMKP3Gks
z0f4NHV1or9gV+zMIemHoyn6PBNRfrqtRD5fjJMkCxT+t73Vy11315wpe9a96jS0+FtZDHzaZutG
HPtCV961Hps9V8DbXVUWSYd+yYS9nQIS8A2q0AbJsntjMQ8RJk1IvOCXUDnqTy236hveINQ5BPvC
dX6pGetv2KsBGYq72YUF5IkXiEDvSADMJVWBb910/UENaY09FwdZpsfgQ3EaaF43IUmfXUIvSxUr
HGImXt5CncOqxjD160CwGhRQNfjcdLAmIQqli99UHZH3Yb8QBSduWwqWQrmU3qPr401ZzjHvXmXP
kx9221LpZsI+jSkz7Unc61Cy1fj0H5O4kBDDKP2K2ov4mlge5YuJx3rmt/RJhQJzTCLEDCjRteSg
lncVqssi/i2D5+TLF8haVEIj4exCN51c5NlX3fIO4yeyTf+OhU/GZnSosHvU1mCG0ZiIvmr9dDTd
VQTFLNTui+1jzi7Ip4ILu1B/BZLpMTC66r4fU+VcS1WWG+idmfnY07KSEWsptLZaUe4sO1gGMNZB
COe7WqSpIAyKwaYPh5I+oHPqhGfBuY4NzgmJ0Yt/QyrGsGwAuCLFZrG1FfIoRDNIRKn0506Z6VPz
2EZAJRBZV/JoJwnf7SaJJRIYBuYIgvWsi6dy07kjBL/5XC9IPdoamCwW4indOnFwEn9JdGgjZYFn
83M/3QYH5xNQ/jL76Z+9B5ak/FoDuiU+2/wBo/Pm4vkpazyGOKhiuzvfFTwpbNfUBIWjsyVG2EzF
68oBeFzwh3PgV2phZk30Jofjl05bRIMxuYxlQeJY9q8F4hlhujbblu626PvRBMfoVClz1l4nBUNA
BVHip2I2cY3S1uZBWM43dniOhp5ZvSr3sSgAYovjywlvN4D4tMLhgn7mbwgr4vW/rt4mV4OU9Iiq
3/4VDqlgb1kGJRT1rIx+9oXyuQvoAIehoteJIW9v4BoIX2Yb1e8uB0+FPdM2D1vsMdFwGyT70/mQ
uC1R6gEa8UP3rYFsSc+4Km7LkW8ze3VyP0Ysqz2JXCB7VX1OBT/t8zSg3ciRLeigtDKOUnyV90wo
HM4WVrc44QdWEBXT5B7Bj3k3HgLxWGFi0d0lF6g6JskUUg7D3URy/TDGkMjyZLGTwhuHJcnEzF0V
vLXyPkF9SYUB9cuk8qYwtsQEJt8NCzhmD68ThXNjRjEgwiN/MM8IkN3CBpYG30HXqP4eeADaJdCd
ZDzXnCtYbc70Z7dgsTsO+0DwTxi5Qp8i5oKY1p0LrAD41ofSl+87G8yY1rvQ+KBS9iztpBp+LqHG
r17j/+aC+auxFrd6uP3T2pFxeJnCd/cN3vMG3aH+/O//7YjMx6miiM0wHiZ61j8GAt87wPwTeDxt
3i/P8d5wSYcY6C0EKTgEDe2MPKskc/WunFevpjiy6BYAkhyXSrwnN0KycrXOMIKKDeF8XvB7u4ZA
H7agyLsYJV7lWNH3XAyBCgw3EjJZXR30zcHEWPw/s4Xd6ondge+zH3jHIRbdOORiiWK2v7GmYhp7
gT2YSDMcBaTXwm3rA5qEVt6K8GZ9gpFUYSle+zzZXuQsMw0BUB7gjGbEoNCvOekFWK0p3bFb+Bc9
0G5J8XU1sJE9YEAP2UMOcA7pwl80Zd/iX4vSh3M90rL1q2yikb6oLkJvxMzWMxkH8/lzKfDsB+pb
Rx8kWMJ3z7+P8QdU3fcI3OXyL+MkCeoQhW1xp9OULAzwU1cH21ZC8iKQdD+5yMEusyKg8wNoOzrB
yrmNNRdLUAHy3z2OHJ59YpmAa8B/xd8PRiosc2YEhl70UCijbkAy/0jAa2Q3o919RiwlVhZaR2b/
gKptO7IJjyq3bJanMoaL9NluI3GfPY2/fNgvqJ3XtrHgXzcmKSvFDdneyCqkgU0ay84ynB/ECK9J
4eBwxHfGwifLRVb/GCBvAp27NtXAgvLaXJRZd5AWyAG41M+3AeTooBrI1/FEiejjYRx+fh8qWZzT
OBDIRloZ6Ql19iGnu1X7mzF+7Rbz4tAUZzvFnLCR/8ufn7AbJyuRtZgZlAsY+ziZ2X+X+5pbW1s2
SyK7z0oNHYG5j8I3+48xqeiUaPYfanlCx7Tib9k97MxNbgx/D3bvn4LCYIOJiZPWLa22cFESl8Nm
uPdJHEOVuTXCiCfPdoJva+owRahQ7WEIQjAUhZxij0DgouCxfYUsxlIutl4UauEh+t+LXMf/Zn8v
RrlUAgOGUY+Z62TcdoD+TwJoCdPrtnDQX+McrdC/GDdamr8uERSYfiK0zLAOB48wOQAE7uAA+IPn
YqZWKZ0Zgn14hUmRZbp7O1bRbosCDyF96HRDxZQwEcq4A/G0tjDpca/P2btUeti3ZwCxcToUXpWQ
76QJbO6D05p2S6MwIkCO7skPvbbEQVPxKSprCn3VgbxcftxoGHsQafEF2BP60X/k+k8tDNWTJ+cF
rGCD/ue9WF0LdXg3uvX6dyGrLYYOQygp2kCNbaSjKC8TuFa6EXGcL7bfK33WlLACPgvF9dUwH0Ej
d78cPVd8t6gK3ct0ZvaMj7SeaSIRj9Rt5zcOvsxEbtMAdK3fAuHTjMLet4HGEFI863DFc5HESMs8
XxF6FyNws4bFEj06dOG/iVatLDT3iES/A8P53pGuttO6sfHRBqKbCwMo3EyDfpSlQv0K50aB1TTd
bfSVNcnqnos2rwOzVIT4INSh11iO0TzDX7hHblGoo1zXcqpwldQ6TxTL6/cHTAiRJCSxWn2RC2nN
U043zQTf6o0RbNrDyUNh7pzuUCWOx74EC1dNWS1zMT2Kkvz5wj/x5QrovqttuGJeF0tHT7yO4zgp
g81JQzKQs8dqE8KOVssWcg2H2356Kcu8EE3KI2QbqoU5s+ntDqIG/eXzAT0BH+i2AbAZyqhiCQED
JPjvxwYvNJTbnc7l4/l76hUnLlvFenGNf0NhPA==
`protect end_protected
