`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
TorW/AXU6/wm/SUJXLZEd40KkEvka8gW2pygLKFhNRqansr+9rb3s8nNqJi4pu4h+GC568H/hDW5
rNLurdXPYg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
lQ7ilJ7E6OA/M+IzYr/DuD6WjLuxukISczm5g4x46Sr8WW85CuQfj1+zvki/PMY+HGMH9JAtSKCV
Cp7096Fy2xPJjxDfgrjyKBvmiAA9GKh4sSAynHZK2zGcTORi49ZHtPkeeoz5VLOgZnSnMFB38+u7
C38nVk2AX/pdXVIBQH4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
paQL0AiQJAezFh3gBESrp3wF9lVFRuhxQZYirMxU4H851Ll4jBO3JWI6CpOU2VraLSeEE3s3vVRv
YDQB4jAakRoIVQ8PVMo+eVGkg3cAb3rWmUfXrHmNU3nPKGMnWowaWkihGl7oWFyPK3eDH7W0n2M7
nmp1ba/C/gfyFP1m2H1f5sQHCmTPdyhiUSBS8wcpgHVytyEJmnWIx4ak+QhpGJi7bBkGhSMiQOZP
Lboar+n/6WJgbVXdde91VZ9CbWWKqmWBQIYpvJAZkB3F5s/g4bFhc4fyUcQKqo2xe4kKVSgd51aD
f969lpaPRRSHu6OgcEVopl3QQLu3o6VaatufJQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OI6lGAzJzR2sY3RqzFVslaY+R/mE4FUA5fTWt4alX+srRiDurgL8W+5L1NjbYkj8iscBXodvp6kr
LP7VGJwXjz42dHYI1WC0zktqS0OAKEAmrs72opfueiFOWghPyadGUmDPL/l3XnYLgAr++rXXqEve
KWt8QsAlZ1PRvZs0LfF/l9nRCuEdzbuNF7C56ZTZanh6nPRHR25FbxBXo1G3FUziPeCLutH+ozIX
iyLU5aKxe+fjd4C9eBg+1PZ9kVnqRgUHS5uBAh4Yvz+xkxxVOzCdpcjkgIAD5Z66BqWKM9mA4KX3
8QotwK3M+PU4lDfgnqq99QM2XJ7j/4xd/Fr6mw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eE6W8ibR/0hWbHMVXu/v6taCP8gIESr7bpnSbXMPwzsbHwS+YgrKfK+P8lTKgAel7ucodBSLfTRj
s2CX5tq0NZzM3EPm4I6IU7rA/uX51FII9xH+C0wjKJz8NJAYO90KtpzJz8ypjBUHaRlNk0fH9pSB
Mvf4wmyiVvPY31eS2k8nCGuB3XhOQY0lzFabZBJCRo1kr1L7XUTw9//cMg/bq+oSfJEst0+YKMNs
XRSrQsnmQvVXdPJzI0SYKL14xeGbb7z6LuPlOmBQAxWRZAqjW1tSYqVCnohIMKCVxO2cakl5MBH2
J16HQK0bfAl14anILJIQaLiO00cKlnhjepWZtA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qUwn8dQIFPfDwI6HY1YGWiIPJWqQpoYKDzHcZyh1zaIYg+sJ34RLEVf5c0XkL17oM+t3DgYq2sCF
HYqsiUn3c4F3Scp4jp5Gsl2rF9VCOkIhUfSA1URkiLFY50Poys9L7otSR/f1pzwyy1n2oU1xIvT5
2jGGBpogmreBirgmfNo=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QU6xSOTTqIAoG7iy7Fw8B7BxIq5jd3eo7XrYP/j+h0dKAgrwZYtZBCMJaw4KXwoIL/vvA0yZudGe
Usn1UEZ6YgblwdrdaAFUHOBF706mtSRiswpXWw/nZrkAXr5GFVDzf1VsTzTuKdnrLckIwgsUGTSy
mfVqdF/B/zziKhzx5/UZvPtpaShEtpA/isGusTjL7ew36ShTf4j1eVu7AQZm7GX2PrxI5Y3d2DRS
PFqwKeah+DZVpIbzt6hMdSO0aMbZsFoBIk6xpy+vUxmwfgCh1ya2fbqvE1wyMO0qhyGvLUvTJR/R
EPS0/fk8heAws1e/dcRxaokCqZaRgLiEjh+ecg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 214096)
`protect data_block
X0ENe4qQUd3xqJ1qCm83K6vdc2tQ5ra7CoEDYoxg2vmK3MLJNxN+Ux2z+mpvVI0/QKdzsxSFNJqx
x4hf953PQ/r97YkdfhmhvGor5szjzslemEJTPh4ZlbGEkAC4Hj9mpAiw++rP9HEHb05I9hArlQ4Q
5oo1w6oVkILvCCtlNpJ//0bSUQzb3oHZvRujNZx9ZfxZYyioccSwIqeD2tWnmuovarc77AKP7S4O
UXfu8lSheBrb5sP39H4qoXUQsfEyL6kQRIaRu3uPpdqJ2eYH80ZO1+1NKz2zl4XVWArw9MiwR0g4
wPqZxjMS50VtwWc/H6clwq2/SCSsyFFjvjBA/o+WqFwcXOCAMUo9FD9fWfGH3dODn5tW0K25Wc3D
9tEV2GXXLvyLDQ+rdOA/GCvPEqgcW+fNEjyeIkOrD6OMiOMpKA+pOLN4s/r6DOYyxXhQh5p7xQ/G
sHVn0LtPStQo50ZopSzQ5IPyNHUeshUGNvC+NyNSlW/fMPSMVBOMSrO0SdCeZ32S7t2OIV+sXqXr
A3bXJmQtC0dNlAE2055aOW8scuEdYjaqKIhMzaRPKz3z6JeB9rNDVRhVrlfScM29lA5XBKY7tzyA
jG+Ay9g3f+z2V8W3bkWr4f1KxAftnA0NL0SlMVG3urQsmMX9DvjtmYm/EoDhy0rTdAhx8WOyQMtQ
AZk/rSjfi+AKevcym0B89iMDl4rqkJrAbImDIXQ/F/PzW7XjK7gb5HaQ78QkBnSD6Dj/iOpgeMIU
ZgAEP6DVubuh6hYBC4CmDbM5SAsETX5Laic6oexa9Ur/aNr7/jJZVDyDP/yu9f1NkxzmofOpf0dg
xDOfn+N09HYIO4q7OjCTxNdVWDbeL/EErKK+am7vjbjlaGs4D8PpmJ4YixWtLnRrHwhkCr0SHliv
QffajpzlYle5DGEn1o8cFuAefAKQcQNPTjE/KRAuYde0Tx6jrp05kQmpyQG+XiyZiWyU+Khsnp6Z
k1q87d/6R03nX769ETBQDi52NnTD9WQ8601D4jJOvHxTLEqMthAe1JNkvSxm2hcBcih5/ElKmQ2Z
lDmW+DFnjhTqCqRwsKQMC1knIJNbcv3O7Wz0zS/KSKErdcOAE8gvU1wYxjehw5JnPIonevRgyaNd
QUSESLncYbJfcrUtAhYEdOYmPekpgeTbX3sFxQGys1wlKWilcSXLPAUVGBN9ZM6ibZf2hppKuoup
IA3eIPLSdwEBxqZhNTupg8AeHUgZQou21gGu4Knbx3BBP1B7FgpvzvtCZGpwTOdbs3QeiwoBrAfh
pjGgaZ8p04kp5wekBXX3kKx2KueVX7scSX2HY2IfMNLBTSGeeIjRyjdrUcVEu8M79t3H5oOaPJDw
DGVfC69HfSzsnBh7Qcjqzk5FMWXee5atu3VSJeA979/lHyiaitRIbbGC+FRPrNtyM83EUFSH9bLP
R4qYww8+c0i6x0dSxu9bgSPVBfPrsVRRPPi/t5RvZS2RPe3vUVvc8f92eregkE2QqtjCQ5VMqQbe
D1QUa7jwyi+sh7LuHbrT5mb10ntLXZMj53yxYFEyhXioo9viKLZreG/UrBumlBVAwLylU7mkUS2W
NMUZ5MtgLZ6Qi8sfDtfb/ytLMuVyw96u5fyrrlc+161FbDk04NpLJVJpORr7T1P+UlSeKPWB7v7M
SlHP75zXKRMHZLkZyolU3b72N9xXgGjUK+nWJu7ZFRav1cxW2tWwJvuAjtmvlg1/mHLfax7KNQLv
F2tAMHrZQ2qHl+o7aVs9MByt5OnagiK/wtL6Yq+qbHzmFK7ZE94rg9ECmDM4K4LOHZtA6vCCG+DA
qm16uggJUZqb1o+VQoiVhjZ90mF02QQB+eGmMcHkOxB6cIugqpf+rG8ug9Y/jjgs2VD9HbNqdHLb
Q4hTdRKJuHBtcqnbbVlQ832ofp3jhkoQhCX1NoANrMs1TJU30tVj8Q/pf8ZjYFMZm9wuD+M9qmLA
JX+BFfAFWIUbaqWvpTI3yJNCU49Mh6DAyeHK+9Gbl+pRAMn4eRZ/ZHhN4gOch1XTVQs6K03CHude
twX7mPbzl5PF5xmFQFVEBTzYnzAlXAWbMCziKXbIR/jN6FlosZNcw/ybhmARaNq5W7q8aejHd4nG
VjqmOKePjNXbQVCzoFMYh3QuXHO8BvVq+h7alcByYlz+Z/1F+tpeccbFP4asFxIX9yaF6qGHoSSb
Lw3Wzmc2YArcXh7qhlw0IRqbmyqtIS0iGeZG9rc2dUOMf8E04b+9EhQykaIT3e9HxuZj+e0NqSw7
bQpA0YZPJPmvqFu53UUMhdqONglYgLaZkvahDCHT55x8YkyCoirEFp58JJ6ks8ifc+PmgGnRvMCD
qmhZjhHJayxMcDnXMvbwC4ngcwhSG79pCjlAYg9EhI/gf+o8FIEtW8NPAqIvSA/98JNOa84CnXop
Q/WBz2yHjcUngN3leUVowAHqnYgDFP8fr7YvxCXYRhhDsBdAXU3Du7e3goIOD0vV/OXqkgVMORzg
ofwa3l7w01HeNg9Yg7ABd18ediqJlp58mgWCsD660wKoezHAE43vQhN2FXWoOW5BZApPmV338JBa
0ElaAhPDIyqbozajq0zzLLVrpr9lKSEZUQ8EaMKq5wPmUL8Wy2y7CtVI8kcTYfWupYpZ8uXmI9Hp
U2dhR2bBypHorn6HwLO4Suva1jPx8vCgFqfipg37C4c54jabSJzTq36w0sPgVIcIPuNFeiW1Pijf
w3HU6T0NYhZnjo/pFQ9Rd3oMaNpnTXjX9lquSdahdjPjcwBmfGF30zkPDJt94gK2s/cuVUevEFBS
qTzGcUW6ZmfCDn0fMnl+vxK9W1QA3yma2A56t2nC+ivachAQUkKTTd80kCoCap7KA4aoh3/x5VNR
cdjOG9PiCHZGWvTNjL7uedSy806/TM1552Hl35VvjgSMNYBF6Wwpk2PxPJ5iL64iuVfLQLVirS81
enUQgj+PgdCncheFKG7tHSFKdWkwvUtuYA56tehZ5/3l7cTBC7Oykt6nRrwuGK+WJY9yRTcnQ665
1pIjHBLXdqMwB4SF9aKB7gyrjQhZY9Z3a08FlSUYfD32lqtvnaLYwxe4JW9VXoLanMKfqlrtxzr8
yU3diNxVX/cnSGPSTM12PfY0BEc4gA542KoAjYWeCd7/eSqTH9v3Q31LbsZ667L60UjBCCjxd7mk
WoQqzHf4Nm3kNFZhj4AYRUspDRaQg3DMUwGp4uKAqArjzfUr+/jzrtzpcajuX+ibrlzJEBRneZ4V
WlZKWtFv2DrtPW2jNK/wUZi3UM2ZZnopFUaeQhCtldu7fvWEkl13H1kHPrTYcqB7eRLJPqQ4AfLA
ZSwj4choenGFu228j1iAPGSMgRf1JWvONQGn+WpvLW27UnruL+9PLbz6jKvsRztfc/6p6IkBE7oc
CNKRYCGkX+Po29tjlWAJoerUE/x25z8IRB9dsfiK1UoX9hED2tspOi0IeLGZ/83KOx7qyNnXClI4
ioFwDsiJSW2eh78muT6iM7GFQqy/YJeaUdG7EBJXSJeDlcyXLw7k47679s5WjoZJbJGbqZHSd8xO
qXLUXvyCrqJ85E1EoCwpPnpU2TwZ3dDipFJEMvqFuRTXVFADnaFxeDq/5Ev9GWRhCGWDQ0Lns0dy
z4vQlogqg5F7zjDkw0FhECJeMvYamKRQXIuFigBqeFKzMkwoMnVHw8nj7zyDFlO85KBh0+Vrf9DM
e8GaDJgweFzpmwiOzTuBIi7OCJ7/BKnC1meCqG8tZ9HVM6ku6TYljCFUe83cesYftbt7iivDtcrY
d9EZakOmlDK2/XayLOlDUWjKnQHA0vKo4s0WFLbzCtZwcH/LknRHQYySKhjWwjSlRwjNzMbQeuJK
xqUIBazkoUKB5gOiRdZycS/R+TatKYlWKkMgglMjkAiE30SIns+Hnzbi73Y/PuUGCMVv6GI9m9lq
cRsozi0U+BWjONuqDmS6osb1wZWsoOy/9UtuexFz5kxh5IeeZRLpWQGgd2h9JfC9Fgo1B56kh41G
gLT2Zh5XiGiLYGTq2F750DS1JvTwcf65Zlbryxn5OwdoirsgiChGDRbmZnrixqR5z2R6HIergxb6
SFdlNIs0xv2eIRm3JdwyM99jS2C15fBwxnPcz1W24kYsNY09JmaLITWg/Vw5s43gsKxXzsppNMvl
wK0XebGn1qnzGY85eBL9+XSvoA0gWTKziTZFlStP1Yb+EnDl/ujqs0eUyqzgAwqy4zoG14TQSNdg
HdppwXje+Yh0jNPnxZ9A6tU0lVHUtlaCLY+/lBEm/0sHhLjetu2odsgc/zkKfz3F+cJ2aOr+/1O9
4EpqPAAeXpRCk+G8vTaFHP1EvO+sK9VhK3eipvbE+oXx3Yulwk6v5uQkEP6EYjM+7wq9dOR6vP+W
Sax/uFJc3tb+z8jZ6N2nPnDZEjqBbl8kYWdc1yHKjg4+WDJGzxkkai9P6cKHMTP6gxN6T4ZSlc1T
tpN6Z9Ubh+H0ABbTtpi6Yk/VtpVIYDDbhNxCO6I+RHsYxYgSnmxBgebL7WAw4UNZaszaDYlvN7aN
ycQAvwU2E2/SPsC+C+jGCY/TieNzHWlLczXtlQk1pyB62a99RomFRKqKYtR5lqmS2DqW5yfDKED6
b/jzJ0v82NC0K6LWuO9z9DG29CdoX+i44z/w4voKPQqu3ugxAwQYWPWaZQF4yeeM5HUG1WIqfQZi
KpXc2nnjl8fVAna1grG392tkHMT9iQNcmywDm/Zfdw9OFmvoOxQOFcC9GJaoSZA0cPaVH3769p3r
ukOxv41y/e5GUcq6VUVyraeWPq7HzWmfZNk77Gei6BNonTEKyPAtj6KIi6ce0cjoHkSO4BDphW73
xnPgVSJCoqcLGIqbuN6YrV8cce8BEXn8KdqXpxnkJVe9kByTX5g0DDOJrumOCmcWeEUdbR7fAnqB
NI9Inj6fMIMO+6E0bjuOGinVYiZJGZDty7Z5kVfVpjomCQUX32KyBNgRgq/Kp5n0Girl/PyJQ7+8
QZIhY2dFxDZMdSbu0uzifHUZ4mRLIZgv5Q+j20tjnZy8TFP795n+w83KTbhR4sR8toYK5am+mcJl
Q04efpDEE4K9qyNHoDsQ7D0nTAnMZzvV+nY6DvqYfYtdcBvG1J+/fjrdWEC1Ias4RkctWq65nol5
jmgZCPBXwbCrl7clkY5kvxKZKURu2e32sLVXzdGnlITYJKXspjuErIluveTyedEVcDoswjDx16ao
+JB2eEGnXuuzMOxpxnX7EjAdTtagY0f8gxtTCF2RLaniRum1q/+86hM/31EUv1//55tFzl+UHmW7
a8cxy8kXaa3nIboVejwED3/gi/7ShKIqeQ7FVRhCOQ2ujo3jgYpUxazBx00kLVOfJHFQKUwRt527
lAXqJAYr2CKKF01Blsx+H/mY8dpcSDlMYZLZiwX6BnbAXdkRJG5NNk3t7c9fHfBIWXa7+apKSTAy
+SkpYOc98I6EmvbEWDQUj3swRrJAUWEBt39r5Y4UgcYmLQEEcboDLZNUzxrPQnkAKy6IbNVool+c
u/qaUiwMWAatmzPkVJKqdtq6noyIoZieNgZMHOtwtfyns6fYt5mYMOULJmAZpYi6fUgP6vhYTa0C
tlfndtL6hPsKyOyhYiMgWllRxC/QIy1sB2LBTF0itOzAu7PbhDnwVpGOpFTz5i6BDl6DSw4Sj/sy
/fTpNlqw1GsA4H8KjCZZJ5PQL+OxQRwmJqR/dwQNKjENFZQYp0l43Ne5NCjO3BqEu+XZJoAMESsw
pMwjGF+tYJD2NXKfAQzwc92jrbcslnVyjNkSfUxWZncUMJ/h7XV12audJ3X1u7jKkBm0PV2V0CX4
inx4dGCEv7B3hxA1RCyMHOPvhpj17pbVlY24WUuLP+ipD4XeUOWLxAXIlUUZcOLD88wlxj5w6GFJ
2JsDFkssExniAVlWeO4VmV/yRCP3DJHoErtLXO16tNOZ95irvJuKJ3bS2k5TAwcUXqcP79Kjp6JK
Tg2sBtcKKxyYPu3wx49M6jJEGf5fT1CSMsyhxArKDUKmpqVysCklGEyzVYSXM7AvIYbpqYn1cm7s
yz08Bn4DzqhYLKpPW+Pqd/qSQQqmt7j8IkOJlytVxG2q+w336649ig7ZW4l7LxeeRBjAxBpJ2ZK2
pv10fhUF4p7yfZ/PJ+Hkugk8NXOt1Lzy89GQfHFIr/Ie4TU8q143n3cNIHr9NN6x5H7WUMF/YUM6
ylfatJdIFqb/9SgyZa+UfaWkgjhGusnl7AbqvhBbE/dcm+vxZIOG3TDwkTPpEqnCdM2z7sg/gTbG
UbeBGQZeboXSBpxQOIeB1hzU+TrW169tw4nxzAn1ETUbr2BRT771Exu9AS/CDByEoP8ryA0Pssh8
wm7sXu7ssmoW1/VFXEvFqd2CrIljmoQI3Ea5JciEvONq45IhdWG0TDdZCAWZc4bSm2iUfk72mysL
F34jJsBSCaDECMCeni1KypDuJwiV81fg+2+txnE++6YyWIzzvSA6LmMXOvAyRP0ZYkgaDj6ZBQdf
RvJCvV5RkRVT5RnjdPRT5EZ8hve3Ixb+/8fSqY3xxghVvxW+UjE1zZt6Oo8OoQAV7CNsODqNNzC6
yV1wgKUDnxABMMrt9+TqyFnoKao9wtbANgxMiRogH1PkPTKMHzsQKrN71mAL8rACkeLPom1ONXHZ
rYfWUPA5zojiScU7lhPZa7Rw3s6dZTOQQq01PvroqbaDUQ1rr8djC9dnX7VCeiIF2AWFPZdv0HVa
+tuDylppIPfNW4qDIV73PSwpBhj7WyuyphPiiFETe9ScjCJA0ZIVObI1fqbGr4sHYZhNlS/k0n1s
UFYZyW63d+EnQuOXoq5eriZUGrJy7tPj9XR/VEymiTlG0t4aFV257o3JXO0zmDtk7MbqvDV8mum2
J5BJf6uZe3sjwFNo0jKlUGzRHRmxTteLAv3tQ43dIeqFe1kNJxHC8bDKdPxnJMGcp2yMakXFD7cb
W58crqaNG8JgxIQn4zqvVIj5eB+fn8Fqaa+9yBIEBkdphLwHIp+DBOeRTjF3KqaEr3w/rjChse9+
GtOVz/EARK2+RjeEn/I9CxKbhrW/UFRF0Hrw6LAF6tDpBXNpVxMvm/xWBq7fsVxOOhWC4mDBTdlx
roqpGefiOmukwU4WE6Ih5GYTUkCYE0VQLmwK8YXAWc7s2Dbw3NX95Ui7o9kwF1iak1sOCDOEPUGq
kgNbpYzX0LzhJmBrCJ2LVX3HYsmAxoQu479An9CnDcrx0kL9IhlIOOhfxk4I9i6nVeu3mQa/pEb/
+eV9k0FCXUFkghgfFJlNN5UZEOQK8KlLrkcc1lrwwZzsZoNEIsPuxBHfJuO8mXk0m6Td4CdN8or8
WirzrHcSylOENzorxHvHAhunjoRmkWYN3y+HhwYTcTMjWg8AFH7SeM6+iKm2PR/OOXUisyAG7bHr
9kKzrth1OxxgX63JywtO5NY+21QXW7b8PTH1M9Ke+IYXO9IAc3cDZrjqVn12P9al0z1p2CAKY14v
udU/0V0am1xVSERDFCZECflBS4wReG671ZV25dQ10Md5lshDFtMouysWVjgiijNb9NIFke+0gr7m
zuK0pY5oCn/fZB5Cdfc9s6pnVzAJUw458eLTpqOfjO317T8KfzdA0fOPME634aH+wdQL8y8ZAgBG
a0YAa7yaCMcZS8FqtipGtdkd6DrmiPhsbu1av/7nGmKKHJbP3Prv66BMDqZtvjbveKN7BP1GyBvQ
i+p4l3j+o3pHVRpp7OszuDyXMx70lCAc6grT1c29qW/jQMrxzweZcIOE8uRvmiUOo9/6NNLHERQm
AYz4ekcoZxnhAE+bkSmMVLHQt70Zp0MlIZgFtm8x7r6dUVnX0FSez98T8uE8jtYogPk2rFn58zvf
xHCG+0L3XgVdACCb0nXKQ0+P9ZrMTVbGG9xgfMfABBo81XQUFQUl7jF2xmoQz5nSDZk9Fr/Lmbhw
Gy9xZDVQwXjbNrkv1oiTsLRPSoGZOEBiyGWaKGwbAiT2Pdrl7XluP8cd7Qmxk+alaLkOCFSqVp8p
qT32IlmEWmbOHiU8zSdsCe7EgDI5uFnyCg+mdQExNLn4FitxAwx5MDDjFRhd+QwAsGERVkk3GPzl
q33S3998i2jMhPUfUrdxtj9QnVxzm9emgkTj6yQxVwL5AD8XknC0t3LTzsMigMib7yJoWiHRCxgD
ZKmFve3rSHEFCyWYb3fjurnigvlfnCAHjsqmMsCPAp2xVK/sr4sK5a3xXa54xk8G/aXQtO1haCiE
e7z7QqzVCp7VhEOVL9Qr45y0HCrMhL0kEAs3RUj94tVxCT8fTDsJBObdU9EL8mljCv427uqEOjNH
4aTVMj6rgyNJSkvooroyKVHemPacnPZrW+7pN0lEAn3CZX42ou+3gB2+r1zyinE7Lz1JWXo5Ot8Y
hEsPXsPkmDoZN8NApfZqsEv+VwOJ0J/HTLxgpsWjvfe4xlESSXEK8T6ii0fdXqfqsE8iRjrTWezG
Kgqb71jekb6grarbUuVVCqQkmZJVSIOS6fnKzA3R+57LfTmSO7tbZjszuywuIR3YkNqBUdYerRo+
UO8dd3s3MKgoJqLEIYLPtNfr1rfza+3zi+rUPNtTGr9V/LXuQpaAKSULojlUrVMvc+4O4wndj09n
4C7rHSK1LDeW//AA2zmmkP6dJGEzipvmwH0F648jPo+QPWs080pYtTT9gR8FZBBqQcFJUcdsJPs+
JefFbv0greOV8Un19O4htYuNblMXuE5chjj3covPJuQY3MtEKztXWL2wB2c0C/4ACgsnrpoVNi4S
cdCuPamtw0YW+FQn1Bi2WzP8D69NPNyYfc6TQtGZTKqWEVnE9UpiuSScjL1bGSa4fSsoHWn+tDLk
x0OSG7NDgpfglbeBZ6KpavRiF61RLZU0QsSv/Fd565Cta+uDGqQ6zxYQpozIQ+djZT6fUiPmz/91
xWrKtpS5q7f/VaAJYRwzRZD4yY/NHRgXgPmGCk1q5TPZMthmqxS26IzH72LR4W18bC/sP++8878u
UMLad8M8SK28a3HWBJa9hweGugEFAXgt+Qq64R2RKAMrvHC2EDAoaOTDyxjTW16aO12pxCaN8cZm
qmspCvCXhW/smeXIVLNE4QmCiuSNSxiOotp724e2zo5Fi2sG8XGKyfIjPjPQ/wVna11zU10Inqh7
D/KmW41eeR71avpzNHF6e6hBJMT7DDV1PpVp3aZEn9fxsWx4BbD6MEW18x93TMSX8Qimlt65c4ac
GtMBwpnThPcspCRi5UmYeFjZDINU18BjFh424qjKiSBCOfBXYTq5SV3jrUp1IoLbjf5Alvjlj0AI
/r3ggguw4/JMRLC1ooruZvFmQIF0OFOU+7hWJKOkQ7wu5RAcGmUAbsuwziQ0xXugbNDbPt1+KUrJ
geTgJ05/kbBegEubmG9RbEznl4dafuMklg3zarAXlmZtDyeW2ljXOwObdWoltB/owUKztJeOP9Qp
fGhy6esCghHS9dvQnQSvQrxm1j00aiKGSI047a65PLm3SXNZNlc4sVF+jJkOSF/YDtPupRVjG3/Z
n0kYkRYUbkaBt+N+MMEPSNMAI/04v6vlvm5unbXXFhZzO3g5zXNrn8Du9DBb8Mboe9uaDxYCtoQw
ZqRoyrxCT39Zau3omDnIKFT0YKYzQ5CxXFroT5bJ4S8c3F5PGVzwFCs2oOtvV/h/9wUA6993x6Dj
4TyW8hEIQCO4vpYwKVJGYQu7rgWk1fWk3bxfWiJEeYyBqdP1IFIGPxK4WNlqZWtOxuHiWO5hwpvl
7Whogko8B4ZcJiJBDJRSESHfP6+g4Uk2YTnjX3vvxiHyiOXh5GAWo6mz2DJrmScMoU+wa15RyGeI
9gMSJQszlA6p/8GyPEQ3/dQJFv5ThwuEBvGnIBq67pVKpx+mrBsjssFYDMa25y2deNrHt9gtgx6S
19mMpNSsbS5zQ1rfbFvefEm6Z7Vh7kunzpDSQ9h/KZXekZwF8jg32W9clHxCMvn1OpSGnbVP7ZXn
JCkmkkH00g+hWb9TxyZ/TFl1u0Xk8xyfYENv9OOQ184TpM36+KheXlygagAqcaS6r4gs2hBEZRla
TQ6re3UnYveaVSFjcYf+HCDhg1HnUrxD1rA/vfKvfNuKIqfE0rW1ZXlYxeLgh2jGfDfLraD/yCTx
KPwcuzEYZ4WU0vgGKCYdGSxA6ckst4W9thp8J2cfUpTtrCcXHW42m5Oha95xRL7QwGNDsIN0+i38
S7djjaHPzA4aNpfd9y9GxuDjTT3/MCGpWPuzWkKtjQOOhft5ugY3Jz+SvlLyYObXaZ0C8e2WsNhT
xo2ZPnF215+81S5rUVFOv+4n9DWh0gJMlVV7rjg5WK1uOVrwV/ET1Q6xhiQUdW6h8welji4zFZQJ
OdJTIMlJg0zrsvsvSqal0UJqf8p/nWQGoBPE1K0iRAoo2l2Eno7OSERDGv0yc6c7f7JibytsGB1J
dYAFyi/yLd8OIcqUNxIuaDEmciN1DAX5TRuZTn2zfEXITxg+bYfYKGOvitI5SDCeeesdo+obV28r
NlObwVr+zIC5JH4jLef8SIhhGlOMUe7vMyc7RsT83Ms7VYRoSxRtPb7F1q9pE35HhPYG4GPg7UgF
ICNIfHbBdWtrO2lnRRrj9m6IO1Owa7St8YAVJx4uu4+zgCBqHk/C27BU6NKKGyVL+YPJjUzG+voQ
EUHyi8g/rGso/vwQF87Gf9FSw0/JgTy9kWpzsPD4jrwrsMu5VNlgATAZ3A47T56sfqznDG5sgLkF
nlf+2WgfZ7l/mKlIoO20Uu82TAUqx0J0pYNL+d94IbXDOUrBphGllrD3dQDV+aeXZPwAtSAZCH6k
DBay+h2TbTlhkbSvi/GRTCPnKlL5pf2iQFMGS1ZXbn7iYtvf8V35UasQmoU+BIGKqMfLWEM3Ti1l
r+RVES1lmFx3mPxsSPXgLp/+0f0oDNSz5FqueoqHElzbeohFF1Qu7LEoALy2wLytjEKMUDJLGSXP
wyqIALRd/VXfbQiI/Rwy3F8b/1AbCbZ/a2oR2FQXqbp1FBTaVf4BADAShKGpo1AtcZsB0YHiaIxZ
2Kt0tMk2BdedGva+1/uXzmPmosbAgORH+7T0cN8Dke4M3THpo3u8Lf+gN5kjCvP6K9X/u8MrF9hb
GtElPIqLu7wWQHbXecZ9RM3O5gMlzfhjfoBT4FQaScLiO6331bV4dAuNNXXIybqccFgJ4wD2NZWV
o93jBZqdZoCSASFra8uBOZEWX/KEoZms60azFxWmALT7bBsrVSHE6IZqApQzcIJGRHV/U9DqhjH2
2ZSSTEOn1Cvcyp0cx/u2xZaF4iLyqWot54BLerI/aKH4u+df01b/qew4Im6JW7nj6BalUJNB71tE
jge8LfxqPeopR2WOacF59RzCuw1Mf8ijaTb/iHZ5wrTjAmQn66uDfJM47y40C7CrGt7n0hoaOdjH
6TiyIdKDI3YMabtEMShJ7j6ycco1Z73RelWpRq5/kGziozCyqFM6OuhdRM1Xh5HVhz54AR/d+bDn
YXLk7D/WRJsz+CPjcIvKog+wPvFnhcuLw34+QNByYvzVU0mglrPg/5gP4FEBv8ZK/5TNrt6Oxoi1
lYP8cg6heufg51geo0RknyZCKhMPluT0M586LUOsioctfZJjCyArpdqtT8yFw4Qv4RPqZ2H7KYd5
mmtA2Z6wZhxydcZO06Fbqo50ZbXKWri24z31wx8kDlaQAX0tMzCp2Gq6w6EBtSMUi0aWoD1DOYN5
78S6Q9S+B8GrmztXzgPXzxE/qJ9p7xvS6YGw9dnCoAHO4TqlDew4m9uTtQzd7ltVb+Xhypuhb4oJ
KR9vRIVtiz7jdcTER4EyEgusJqSdPbBWabVBdlDpJZ2i57GlkMHqSsJEXrhJZY1bE7Abe40VSH4s
jWpA2MU7XZpg5x7w2QM7AU2O+7pwbT3q57rEiCR/7sFTdV8THb8tgfZ1uxKJibJHJ+fN+n6xBr/H
HcOZS/piiyI4QKhZT7sy9J9Sh4j+I9C254vTT8cEEWdN7+3HLIRycDaAJqUUoZFfevSEgJOI7Kc2
pzJWHbjpvSFDMbQEcLnZXo9zDnVQw0wHOsYxBLAAGeB9p5Hs4oXdi1rN2srZC5uxu94MFaP4T+Iu
ZkOpFoAWbZ8nb5jXwE9nAJFBwg7G4knL6J2vlTNTrRAh2PfQOzE1T49VllGMaos8DnXhIRxTYGlf
uhiRYMLOTeAyentQiOrs59Tdsmhu9KSPmpmDTUwTKDJQ9IdK9lGNqBc+uz98C3vgmuf7TvO6Zz/m
JqNZGxNz/baA6TDTzbPBexY82KXoLbq5c7XruEZJ5dNBy81eqxKvMdgDUi91ISnusMpMaqTVAu7n
LaxekwAbQZsD3YStwW3va3NgU3aaXYZ3N31ww9XX+vj05neBpbVLPSOlANK76IEqlVSk/mSDhlKm
184FewdDPMREvlKRtwhU9A6CkrVVxC+Lw4ufGy18VvL/RAnVv5kIzj7YAKHfsr9vxBtLB3qgr/EP
LYwQ3550I64XoGQXEpTmot2S6kQ5EA5W/mWTnircaudJvV0EMO7Y5Xd/VJNGmGzahFE9pD7NYueI
6S82/FuLZ3RYpbdsU2bFvo8mgZ3MxPv68XEaTpXUskAEJuCtjBs4af30cGTkQc4/2tk29v42Uyki
6fAmMS+2qbvAKE3C7gzw1IHbnETD/wnobJhmGagGzg2rivKEcBXEM3HSlTC5QPGIxdfyTx4DSIlF
CWzckqKHTtsWnhp2h++JIIyxGiRNkbeVKFcPbcky4NlsRvg9W+DgUV4c7yjuYEf2Fis4Wk03oNxG
XwvhvuIwLgsfn20hfaA/5uZ2HdoDAQxLQneH+UibGbJ/RM5Yma+j1AJbYNkQNTo063WRPFiNclk1
ewFN2tE+CKFWqH1+1H2MOcSm4GBwUOvFzLvdR+YaSpa+RR3Apj9rYhMmvUiaTGPbBml5q9KGfwTd
8ETFi15rIH0Lihe2Np9monJXhPXV1Gz9FVQnj2owdFf9PUlqRWpnjC0Ggc+UqOZk9cL4AIe1j9SB
XAfs4GpaB21/RyTFFRQ9WrGQXAUopmjCcfOGfActhV5G396ScD11H6tDBkcmY5uGntm4Bfr+hBHD
T0j36XyyVuViXD1yImToE+jKumu6BMsfwlvQAJraPqSoIPD6T8+rgvLxB+BJZbXRxne5dvIDgisF
WEmQZLvQoQJL0LxAKH+oRZ8kfr4lUa7HPe5EUrcGg3Wm0WLljpUNDdjJN2mcMJr1tpc46MTqEEoS
d8f1DwPuG5semKk90U0NQNceWKk3O09nrEQVZOHs0kXjwgZ5AJO/b4vD/D7og90J1OH02ygU8bG0
z3Rno+H0BdSeVne+0WL+EtmO6pDSTP0b2tbI9H5CnKxqGQr5vErxBDW8CUyLbr4E/VGTvHJJYe16
wmXacYdc5c6kv2RICZZdbaomOvIQtpfDnnK9tD0Aj6jxsTo1DtMWyN+NzeU0KZ6TRrqg7aJyiclx
hbS6uvnv8h7MpCfnRL/XkrzQ8i3M0flQGHG5CmPY68VbO0y9rCDqOP1EO343iJOXXrSscfdF1kQj
Z9+ylo8e4Oy6ZShq4/hCrcmdlojMS8vfM1+dSjqvqTv8aQb0crEKppwwoIUz4EXjIpDhztV/edyS
f5WrN/DwBtJO9MppHNITr3DVff5SXeX4G0Bdg115Cs8mnK8Ek/itCouJJGJ/oxmfOnBusb/0tM5x
2vS2eZSFH7J1lwKt6A1IuYwoypySd0KhheqooaDZIMz9ZH7Li0NYf1JoR8mEszr2+Vp7O3IYwxRK
CBqf/H8kdmYKRSZaKb17os0r+j08OiinWukH3kcZ0fw+6DDh6D08HRTfECfZHr5NAKeatEmdqrlQ
qK06Z0dM3a7SoX20Ajci9CMKllS+vocUfFWuVASvJ4npJZh026ZOr7FBfMjQuMzbUODIO6E+GSxY
WhzUPjM5QZil4WlbLFmuBFquRP3KokClQNalee0BNm9vbVN+S0OLymq0g9vPiQeyJSI62zupu87n
gyUhrMuAM7ruJStDQNO+W7lvhQBa98zSqfJPFKWLskbNPNTA0Pv/cLgUgyKZLNwFjWS8Ce9ixx/Q
y1dj/fpBxS9LkOhIIcnRnV9tEiJiWfBMWD9dA0x6yaQFwaX52xVm7bYLKl2GcGR/bCNzxsVy7MS5
PjruKD9qsa3eH4hEdrthTHYdJeHQljXYgT4zODLJpMDVxUwUwoZQ5911UA7+VZ5QrXROUCmQ3ARV
1VKDSzNeTCTAUGr61Jlsd+5cszNRCiIRzgYw0HJf6YJ102JegGWm3e7c9jTH8fOKIc0wAVPp62K3
PnsOL/eYw5NRmsxo0f6mwRO8IBB5/zH3JB5HQoTrAjjyqwfs3Y7a7wIjs2HUvtHId4MNKUch2Byo
0JjEm9oPkWtvdlCUyQSZjCyodKc0BYBNX/HBvDgHiCs0EYD98pz61bwh4G1KsATstzU33Cg4SiCD
k6UurgE+cQ1Z5yk/raNcoaGOYhsNc0hFl1k1UvMzOgxka9v1KgpWwonj/RYSQy6jwJ1YyR1VON+1
a8WoxKfn72TKrmVSSbbndjEo2TZJieWQmdEmBbkXYAjNURLiPEtpzLIqO5rqLAiaeoGa/5tuUxDx
r4ADyTS5+CBg/X1HpJVLFk+OBjhwC/Py3oB1tmj6YjzzrrFxv705lxE/pnlvCHVkSPXkH0fcpOf2
QaWKtd1OrktDLOzYlKmG721rNwZhasLYgu7qcUF0aMy21Fflu15JnxA4m85TPBx8vGgVjPSF/m1O
WnqY3RW7oZZrCLAXFI52d5nzll28kJ3xMnqFRra0CBYTcPx1nf4RIr/aHwi3l+6MPxbrrHM8V8LN
ZvqtgUwkh0BAJ1MyS+5aA0WMNluu5YlBZZ1IdgfQAt4oUQspOdra2iDfXZ9xXs5Cp2RUEF919+/+
jbP4bFDchTe7kij++gfiUXhQ4J+PL0ZOWw0q7NrbpwvzPVhq4eUuLRF/XfYzVWF8A6kUInRzajwv
AiCqervK9TWIjeyIwB4DTvB/0GeHQAkj9KY/Lq+/S+4klwUubvyvxAO4Jmr5rQsmgq6CDzHcY5YM
nhTIU+JembG7+Rw6TdII/ztgrazJ9DDLWBCWtJbiyIWS5RrL0r9CSAYVeDESn34k5+yqQwJRckTu
i0+Dfcq+XFe7bbbLtsJRUAmVxh8n3ADTjsFdQW1sPpU639tzDmUvObzZ+a0KrsIJ0qJBueENbLuz
4uoHV/gGPxNm/jDU3hY+6+hwasreOkhQFRpGPPVqLfzga+zYOnzN0FajrIodh6ooFmYQzGB5AVaP
Zp/OCM/+wCkIgawVvtHj2coG/alYiiV0fB3FTiwSsmQ70Y/0ia/jkZyhIpq2/1EnZPL7W2/oPa7+
wzUAOL7t+1eV+9KRcFqCS878DApJRk5wY4NOh2tumQf9SSmsBDDdv6TVZCsfG2TffpeoPRFGZkm4
88egZBOF00y6HMM5FN/T0dsO6T6OYzHPaJfJRrD5bS13wAdnggKH895JAXn1rmT/dPvZyqs/vIue
JWQEDyQ8oQJZJecJD7L4XGwtGatdkGLDom3diJ8eyYCO3+mhzs0kd9gFVdkslvRHIc6Ikdv5A9Fe
TubaFf5HIxKa9fid+PiVUJIQfH5XkEXBY579Au/NMcGnFyqlXyiScy/xVAOTxIoc4+a+Q+sXfUPg
l6AnvVPR7C6ctfcycE5T3mIHYFDWQakjSrmqROTACWjjBAyylKsgDpA25tdizHpVlAHvpyHlqMp7
iL9QyaE3t/tWjtSUMlFlREe/0yQKEQs2r1HWBaQvQfqae9oo+uoLHewybmi681jUkxo/lH0zwO4g
oyDj3/wpDPE3HpdrisonifsgGjHOZBG++5hpLNRGBH+5vlLcLH0A7x+ngH480zZ2W0gDtKooOwXu
6zbHKhBLB8BdwMoFNDLJ+DC8vnMFEjIHDdmVwcQZO+PL1Hh5LmHtezfgwcGI3N9T8gN7vLe35E2m
m7wasv5wQrT0DPtfPmXvo0iunqOFHk72lw9eOQy2ujgwHI+lpHXdz60xXEhWGVIeogZUJF6Tc9Ty
W7gpJPk/S182k0mvC29VnXM7OZ6CSUHtCHfyDm7y2BrWcv3Dso+3qlM3P9Oesw1VCWTZSyhkqLN1
JgOEkPHbNw9osR18EiGu4+Y87/W+IXUgvm7zI/TcVTIKTe8nI2jritQ44pheSu/BjbXEH4sIhSgF
Lol835HioclFDaxtpgEftel+5ZNuVSva/lI8wc4LXrG23MIlmryOuW41J7m7SV5EKQG1LkA8b5jC
TyoxTgMwiZh4nz35J9AllnIJgVnRhJhs3BFk/E0+9D4IDuFwmxktKU5wul3EctAgT65kAMy/SB5z
5gvbWf7DrxB5KZTMxKVXX/9228lc6kS05/QGtl7T0ZQHIJjsz2UqBiE78ZVjyY0/5CH3f5YmzTpd
qJYOcC0qawok27wPQu3hBIxNSM5rw2P1/Q+QGHXnnSXh75dREQtQtEDD+MqU7gmXQ37CYudK4Dm9
f3A8cM54WTzLEfux/fiarRFN3Y50K0FBAZV1hA3uqc+OuKzIYbAW5rtC/H4WGvswJKAr6+KyfR9t
pdl8x180mdylxv2bJbjUZJ5/49gxqX5jdj6NFBlfY5Amtbp/lp4EZsscQe0biaXJq0OtxNmdWRKp
zhpSH28Fh2AadYqbRcDCPQbAZZ8YmN1HXuI4ZmqrCCZs1ffcVW2qg9co1vl2ui+G6uk88MJ/aEpf
6/6C0YExhEg1IWmFJ5NDkRfMqNMlz6jIQf6LlIM5y5FNgZGZeLpUi4MJFyMxa0pCaCFG0+HgSB4P
n3MXW4jGYjYNfY1LPVzzDiEqLJo3C22L7tfzZpZ/8nUIinz7rrlyfYEJ1yNj1NoC1j/YkrUnpRmp
w6ij9afCc/VmO1G3vGjsa5ctTQ2SXFGu4Iuzf+nbqPPDE5ETChI8vRkatHXdXwYndpOyL2O8sZQt
2+HszV1pqpGf7Q6CnrsxJkVLj1rtoZEUdLyhjggHIpVD/3rH7vrSQ4t1RpEKCK3N+Not308mXIR/
+9UKayUnbdePWnZhpShZSySQJkFYZWFuPfNqlkzMm0nJWgbKZu61M7K37KlLNAo7cZagP+pBha2P
3XOkd4p6FG9jUjw/gUG/9RDrInIipAO+RvSrXBBhhfyo4ZnvFYgx8Rb2wo0Ope8AmeLTveHuAO8j
yZsEV/XoPmSDJx7Lw+p5qr1zXCKOwcG8JMZ9P9U6satFxeV4gi8oOQjuIjaJngxup7ds3JKOVs2d
YzkrvWEVn5JxIXaw+malJKYjPTZs68j+leOyq/mzz4nZ8a7zGFkatHL4eRnzWO4arJ9wt+n+9kM6
ackmz0F1ibbyKM9eJMwho35t8zKwWgmVd/+Y5hgVi3QV4seUjELI7CbaKylV4D9etcTBzAjhpgr7
O+1LXaXopJtSeTcTSaREwQ7OiU2L7mNFfJuDdmCVjMH+ktmkYwcjGFzftqnZC5ortZd4LUyNPB5h
Hrx26S4+ozvaZYyFFSNj3X0vFdcGf8JkLvHTAVLEeLE79ChI3qkY5zOVcdWwP19b0QtLu2gZWeKL
/sIRPhKYrbHZDN62yEEtTuK6x7Knd9NLy8wvbC2dnmQXNpouy/l7lX/qtO0axymn4Me8NDFvKtCR
vI/9XPJr9RKNXMLh27zIxnEW7JSSzG8RpsGtOf1EkkK2Wod74fiaIpknsyOT/Ece1gAJ0nNrDxUc
RWwnvK64EQeHsn2pU+pqMTUAD7ZI+ekLcICOGKflrnmk8l1UT++BC+Hhl4r3aMRqMastiHookhXJ
M94gq7unHEyX/otD2HEtajKM3qXu2HW7mBKEAeuiRsRGcPsFnk/SenQgY4AvupqKOu8xKy0QBDez
bqcKMXB83VwcPiKD/GiwowC0ZZ8sHVQ2Twivn0iWANSJkWVRF8iErBOuqY2+SRxmATBndUudZ77k
rn6kvXgsJrbRnJ5+S547TC2ML7CdOVPzmMvWdBMSodnZzquAqk06hVK/WJYeaMJCrwivXV4sBTLT
spy5sduatc27sVsnRAoROWHqS0ES7J3JcZ8k9oe1l3wasPN44SFKzNquPldMN9TXwac0Opos8mfX
khSi32VxcMpVdtORIHH08dV7V6mGZBhDAMBb/bvMZQprvXlxJQjoqKr4iNbbbhYfOxG0sumbTy6D
f7iPIsGM09xpl/wpSFrYCWDeSdIGwPaAeNz9tUbEWforVakwNXcwyyP8kibQjS9oGryJI+T/5zRe
DDVh/Gx15W+cTQ2n4cgvMoeNFkur7F5hLNxMztQwUR68Sh5BUneHXLeNgm/NwuB0ZbpQoJNIivSS
Wbm5HLHolW27ZFkv45jtPWGlV4nTVSQqd/43emfWZumioUrg1BDBe3uZgdTOxMOhXoW/OibxZ0Th
n0QsZ66ThJiySHn6PpaWFVBAizcXIVtfzlCkqFpZjxBdRejjpsgL5p22gAFpcEgftGq63BKJIQ0c
bPoOQErxKBsoIq+gtLtlZ3BXKdxctqnN8+USZx6OshD//pLQJbar6Y+39B4t5/VpX/SREMgzb1lP
+5Kaspd1axQ04cbHUrpkFtfyHJSuS1S8yVkNTdypvN09GqhJTFvFU9+Z4xmy31FlSosdgL2IGEz/
ADt8V5jppbL2EnQTTMk6YrR1KoeFezz1Q1hNJTBpuRvehZDDcOqeifh2V8RtqiHXBuAXar/3sZEo
tkftPSixr74okodmnn8rwktB/wUtEtT1XPhXGqz5VQzxxUYdJ0WK9/1Fjka5FswLDenl4129H5/J
dDt28EYWMv79/cAPKOhbGKrZAdU4LexqoGwDoh+7EJm7NF9x4U/sM+e951lLAzhuTvjRcKnXnOmb
aWcYe7Q9MbI54KZ085jBOjaRRBdgUxA5FnF+JGCINY3UgswVMQGQYijzEh6P5AQxdVjgYw2WPGoQ
w0ilJuRQ1o+mG36TokxFpqVC7E0wOsKuEKRbzaTpNHROMsaUG3Vmoc9o8uczrMkzGVrQRt5IHWy7
eih2Rkut4pldQFoQrVkoSqAcc3xhvvaQWM595bKYr1k31Tl2N6MpQgpljiiy3kR++SOHZRNp+5yg
PWR29r4AKe5cMjL+VtfFaTUmsBMQv6qmc1f9Z7jDTRxiZYRX5JWtDUfzccHf40G/pGdZj4ZgAzBJ
sXhqcUuUvcxJyQZZ0TJ0dILWL5l8TtYB7ssp3x2Tk4xkzdpQ4pFfwtywMt3q9/fXdIFVHCZzJpc/
RP/DDgy5H97vB50k9IQ0Lsuq/Z07WMplPGyTA10tsJWNzo1ndy908wOMCpXD75zBmv9O/AXDHXLl
FXqGo2RXP3e1IJtqAbZA6EGh744o85Ber6SllJie9G1ZjSqTf3yHZatgEeds5m8q34bIce62tNqY
M3or+rClKniVIbNuvHTLkZ9qOZmEIdHS4zbAqrkDBJiVsyjJaTCx+fmfjkq2/TGVC37g2Ha30stc
+Jb4m39s0NCDxCwECvEMbR+DOMFzlJPagnCN9goHJC6ca9V4nSybjqugX5wY6reBG508u/RANsgp
sy9n2wkARv4Qod+07gzAVB4AkDmPPgW+5BG/s6zBexO8jM0OtkTkWEagdsL9CuQqvhqLgv1h51ny
8GhIG0kBxVlntot9b441bjL3WX96NpQhkkVmHfiSdLYXsSCgV66+iG54/O+GGVB2CMl42dVHdJIC
ViigfDqseRSXaoRJDunVV+rnCNhotfboLQUPBjQ07Ei7bzE7NZtu5S/47wGLC7Xo0RAs6dJ8J49t
WK6A9+e6A/X26+TQKvmXMRyo5b9NxJ1dLRtS3oq2ZcH+uhTrtQALdW8OtOe6s3e/rPJsvEpslSVl
bD2rTZuG+xK49+0P9GKPlUb08H77U0XgwC1W+SbaAdCHEscHtIzQGJnnqlJsCq5HYA5sS+TUNUoZ
n44q8azK0ZMffEkEkqchSpmjW6K9mz/lL8uPc9/OEjEdRsZNFGEVxkyJCweIVW3dl0kvRapgDfM1
Svgdrj6dBrVQiKmmkgLB/Ml4TRAM2eqjC9K5Cq3B5yVXUGpA0wcA4gYO7x95yTtnqxkN4CKve2Fy
vFJHvICEFiLu6lsGt0UoGIo/lDF63r+acw/9sercKNb3nh5CyfglAms1yWGWhDmUlHvr58k/okxw
AM51SP9dktvhNxcN9AIB5XD8kZNdvUDQitEQZQgIVsJQCKf1xS8NmvnB89zuRP5WZvttUNSIUFK4
fcxf2UbE6Sp8YFIlkzn6JOZ/rW9eyoIpe+xjRxJDQCx5V7H1DxLLnHwsaSuKY6KZSk/S8yzc1UQW
3hnT+g81hdI/CPO6X8TeMNvC5ktXdB/c6yFuW5jM8yIiNwj+GSPdUYh6uv9kqPT0N4AoTZ0fSFHy
GK+ol3UluuXxxNZa2WhErhqYY4p+0mERCIIO/1y/vk2vfM0rOghIhWlD1THvr158g+NN8o+INyjN
TdrfymleUuG/7qf/qLQpehcWqA8xKmnfKZMNwAfbtSCu5MAKxKdJPrCdZfzx5ft/3y6UXlvz5gu9
O5rUzT0GxfOT5hnyVZ42An0wpJMeBCdzV253tG6G8a1cUykInzfUZrOtXxgeXYd0FgnyessnfxHu
WCTs7Ejtf6YALPPqv853G75CLtU12nrnsrhOeLR15c6IgAP5GafVZFrcChVJyKrHFx0tgXofKX6x
BIhreTpBNBg6FS2LQkjWkybpb/N0FD8V26QY0X4J+ci+y+ZiR5p6ycHfj70Cm3alnIqZFn910A+K
Dn9PEKcKPZlDtWfjd67PFopH2kFuO0d7r8pikn+9xIxSuFAIjS297itKBsuCsJSwy8MaXACj8u/4
D9jqoblzt5KdwI1HQbmBnuIgN7bvWyZ/eLOvyQFo9TG1pkGZC9Di3KIjHFgyvh+lRK0q8dbAEpfr
LcIbtpnC8nXlkH6sEOLnZLerVvk9Vc7ibUaMHPqvGyo2Fc/A/p/akENPi/eMZ6B+TGDWaZuGw7VI
4McMncJyvEr1ukhbNpHG27iS3xN0TCGBymHELjLN4Z3lMGynMZc7h9v9gSsgzegmQWTRAixJW4XJ
VBUI52NQb66sQDIDhR6nTcLrNLjWpDlTuaKq43/Euc6NNrqqhbf4WPj1mhLrr13SGFYpByLyyBbl
hG+ecrFrlkmBoW6dQXnnsdhH2sqxlQzQETA28pyiAh7yh35toQVKLlL60pUYho/KVqWBnXGXs9xT
3eP4a2VPr6hYMg0RANn98ey7m+Ho7Coyo2b8D7MBbyTBH7S33C1dJuj/nd4Q3F2gpPCJdH1rduTD
s0aLmGKe1wBl/upQsZ8bSvBcrBGofcrAJ+JjftnWzQhnckclHFMBbxV+/esqIxxpBVOMl08QWkjm
VCNy4l4QKibAH8p8zfAeKTm8uRmPZF3qXvzdo+Ns7lYap+KDfK34K8GWyI3Voa5G3cVurDZfPMxp
g6mqHEvp47SJUF1MLvoawix55c+82C7/vkeGRk1wdq+xwhuMp9XUoZarTCseFu5N4O7laUOvi8S7
FCdKGGLCOIS74o5F2jeVwEVarJuQgkjuyaZYML6bbORFS6j0jiWLO7TOpnEu5o91k2tGK3B2Rp5h
aSf+9gYJSd08+L3x0pUx7XTHlYhN1TxDglRhW9PNcWIPwu6EzDEBKdv2CXx3/aE1sZYVEgZbukbU
z0/QHuWEN1T+FIXeiFno7Bogc6Q9iEDMCVjsidQJa7nKOmfQZAWNKbLDfB+HXx8G0+HkPyphWwJ7
+zRd/Xs0ri2gK+rkHcooMFDBFmFvJcZxQf0dASIjTr+f4neQeB4MLg+TV/Y5pjuScXdhzOGNyZip
jrMsW1sOOOOocRhwOdUqS8yVF/RZLidD/IZWPOT83O25XsqjmBOFLswCWES2+9ixd83uB0veZUTW
nwUnjSlJK2oGj04ZV5rKCAEQfKw5EpvTkgo37BQU1SmAt5hBoei1K1sQSmtst3kquLf8R2YqJ0ik
S50q4jKuxeF1wKyeHBv3JJYSTbRy859vWUvSHPs9XvXs7TwHkP+lebW5d/7BBDgq94r9SXzSYJvl
vQbNxztLfu4HUI8WoaJ6wKN90GNo4KBfW/5LFcS6fLbt+h9rp1Yw72em2hwh1/O0LhAUPoY6Vr41
2HBc7+Ewk60ZA4Aff2HfP8YB0y9L6gjLr200uxe2RFTOQtgoaaYR6CUpakkqq5Uoeok5Vt4KEa/G
PHQGGOFqnTm/ZUY5u+x6K0uAZrQ8LZVEyaoxrsSRAh+4AQs3WL5SgI4VhvWKXFKlFeYdTLT/8gDW
e+OjotNgjG089UfFez+ZGmvjEoHtp/H5nbX38zQ0AMCsSSxpMoM1n3fVd1qz256D3hL8TicT4rJd
evzhAjuVkfnUOJLJh+h/CdEvcN4pYnB+HuIlJ1utz+7OA9kIgj7l2ePVv+FVpyEDlfcK1NjcMyVW
t0wbQZ0XqV1dDMS88FbzoFtMIPobhjfnUWCewXXK1ouSl87kd1weqQGkj2UNYQFuNlkDaIn1BMMI
cMNvvkhQ9f9FUzeMOe4kCPRzSwkbeL6ooS6yQIBNqpLg4noAYoAvihc1MzF8u0irOWox1fKWN2R/
qRbmKcSsbU9kldJ5QsLrTPsI3sVjbhB9eUv2Imjxa5vYMbTJ6kTvjvMS300T1+rQIX1jtTNQOOQy
POYdQDCtx169FJCs3Kf9DEaCbm5aDwycI8nqRoM3PMunXEBeFv7emzmB4RQ0xYO8aFxn2HxFubtx
JpiHiTBcJXR4llMVvgfA6UQ46sBoq/hmEiaKKUm7orIJ4SSnFjCYzHZ2EdrzyjvzX9jp8Whmm3V6
+dlEgwteqxHuri9zn8ZyYhxAXfVfaYLfwUZVngl9lUy9RTl8ThT+63FFsDBB4Hre3qASMe8b2Kqt
dLJqcvxhZgSgHA4VgppNijZtBlN70t1Dd2mJL4xUI60QW3aGfrhfNAENMxfn+p24Vu0wmW5I0ykx
iJsXJrQpQ1m9Ey2H3rV9LtrzXK2QttmrWGQ9TAuGovgsQ8IGPVzi8PR2nzpQ0DUbWa327kKRvu8o
PyrG9TcNHH7WI593JcBOITlIvJvyiqjimnkSM884P7eo92rufRuixr5t4R2QiXIi7wH1SDqX/6gq
Ez8cCy0YucpNlRNx8flIbbMWUdvumS3eqRR7iXQoF4xS0UQ2LYzUYbIKXw7znOazj9iS+acCzZFS
HnFyxOpX6YxrEZI4Xi3uDe+p1eyi7HebwtvwIyXb779uWRiIbS3mKSvq+fF7a4zu2ut1xbe5ehXX
V4v+ur0SHEGHkwTYfNtqFJ3gKwVRhVWISSpU/hQpHVAfl+XRqhp15pQC7hOEl2CoAOlS5b7hQ0+X
+RigdbpOxmQseALyVxx6ssc+5k/lFXQD4xblJ8iW+AslP2S2CPjoJ65X/6vCt+Mk5IN83sQ4RbBy
ojAu7r/oVzgtUBbq2vNQrNwwXLcXRtQnvWLVcE+zsZxG55Ck4VkTSsixqPRAHUjDCLrK1A/zMd4F
S7es6TBnGb1ZCqsxHC2BOZZ9cCk+MaeSsFkVQ1C6G9QUh3nH9K3D2fYwMrohQTsTecv7iOsJE0uT
HPHjuBI72jdFMCpsVKCXnm0hMeIfG+6T/6feBEDzvI9ImKBIRbum5tJ0e5zzHffuBqBTXhe/4k3F
YgVjvvI7x+09zz5ktyOrfWud5iyowso3/FOeVF9jF8j5AjlyJKncvshQ1OG5sy030GCSheQI24RY
WMuSG945jp+ryz2Ds4VW7+1hCe5hI7Ex64Pbh90gQDK3B3f70HdQ02R822QC0ZV5ghH4luTIxhtB
E2ZOxAwSzFDOCGdOFdY1Gx72U2duoa3aJWk5+EmMrOXXvJwXvnmu6aVO6o0DYMAFPZYaWRxp1GU9
qYS54DOA34O8wVMJ3JoTHHL+eSQk6sOIbj0DilOrKCorhFxQwGR8RyZHzsDV8WMBAs8GWEX4l27f
q5J/OB37eRI1wZJ3Tp+PWLodZ+W6PDCwucgGmEWXXakmp+XwXmbwqepKRFmH86WhCPL7zZwX3J4h
WGrbBy0a11bpyez71UvDK8tgokkE3TfjC2Fn6FUiSj2OClH1WWRHkAln9ZmhUTLloR+FGaSlq1ay
bpL2zOjLAg7mX74I9Vvmld5bmoULkXHOpcoLPAQh6oB89/WYLaryRHu7lLk3+bct9yv9SRUp6j+f
61FCE6ItiIYj1ljVWaUJv5ck5e5oIrHaB9SHNdNpZ7pXfpU/stH9y1Ns46eCoq9UFp9pEX9AScRU
xkBABDpAueGVDthO3NO4Iqn3NlnCKR7h0nIMSBy8FWZN8rq7WauZeNGyCNVBkXw4U8+mHNKzwF4u
nLkj0Uvn4J/RGRIMkDIxfX2Gbinm33KAfshJMFfRTbB6NMmKBQWzixi57hpAQBxzBseuTSF/lKOj
E51a3n5WmIyIs4qYQtWr4MGCJ95D4Sb+l0daXPeElXEQjSzOMmNkAL8EYLPxWh3uIKDpz+++/UmH
HnF6Ps9li7afjW4kQbkP9R67ugzYiljQZMkKLxE5KbcpoQUfWngikbgxGKvGW+yJAsigZWA1+ylI
ddu58nfZH0mWGE5Gbd2S7T9RrutTgAz72wBDTwaHcueAazZsxoGCOpqd/rHFwv/xdzhbpZ7G+NoZ
9AvHwbuKYdgmuMfiv98qFNlJw4TpLhQ1b2KTTD0hA9GW7kcLMTm12GbckEl3+PhM3AwTt1cTuAih
ZFGtAAjiko2AlZszGBPyZjHBdXb/4LIIsNIeYlVnNNVCAqDCKz8MDi+cBgzaykFmBNs+ErwRLLfv
iuY+6yHrPk2143EMMglXG6mIwhI9e6FGFsY2XYRqtX1dL1++M7TGssweiPvmGlZjp1AS8OdKSl1F
rbVlvR8r11jCWYJw/gXMswmYqQEOdLq9eQFAOgxqa1Kx88Eddgzj/FxXEnp4oewIJTp6c34zcpqf
6rMAKlN76YLEykbPmryft21bgLGJtLExopbPELhcZUvoWMm3sPmMs4tIuE6fWQzqT0jmfr2broMr
3imtcvyx9PTC0BAc6PbQ2XZjqDaIGK+t7YCfuNFAtBjpW32vc6awpB7R6CBwLNDHjBi3hDXfsyZR
z4h2xSJeZfHHUje7hnZ90cNgBAXRjp+EslgNx36c7akVxE/+atmj1O21jHRkPu+XU86JsoCAa5Kk
GfvYyPoU85JM/GRTyeQTZ/N4sbaFOFbpec4eXGnGU/kCRzAe7+mMDVVKiWN0vOuvdglwvbcVBI+p
An1W8AWcIzloOih3M8SPXc7wDNb2tQ+b2VVH/vHNjb4O67o89q277PKuzO4P1HhMzh17tx7CiBUM
N+wYuVwbWEI8JEy3RoljPr3pZ5bpdjAzIwL67g5PRWX/iyoDqE7hfSa9NfsBD4ehW3s99Bqmu0TM
mXmVCpYjN13lFea0yMfFtMEKro2U5cOuDbtMGIypjvy5BDZ7nAUw3fm15U9Qf3PW99NexiCGkLt3
yp1tck1LT7qPq/H4TVOToub6emmcISwCi7zRtogyBj2OZempU3xLr4RNGnCn9ldSaP/IhwhcZMz1
U+d7DwT9nfWm6geVYgiyIXf7OucmhYjzECAVAq457T/euStQC+oi1t7ih9N+7D+zVX8nAP+Uaqbh
/kSZv52Nak8zGDhLbknTQg9EB7g80R52cm3zgA9tlrx3vV25tGp1ZeVpXbj5kQYWhj9un6ivLkfs
59uO1e/B8xfRWmEdZ2eye9z09tzt+sQgSu9uW22cQOhuMayqKpnYvk3KQl7/SxzOrlOvzepy4V8d
c72HVcgPXVMI3D5CqRWeLZef7KLnJEbyb3XLvIOBoDYDtQCwLMIMaZKcX7z/1MGPOliLYQRCgdmk
Bppt3QYcouUwG3H/S1OYx1VLGFqkz3TTj7oinW4KE1J8zYQPULa5iNFfZ2YPURllQBZBRZDZ9Q5x
OyX11B8Kv0b6VeHvXFLaJFJWY441c/2wJUHimwCVUWlz6VQ1aklr43TVuI4BMq8ZAGyepXclE6Nm
ylP2ZGvbOVtbMzDillwUZ8qmm8WWR/z2IUO7IG1nF1swl7oTAIqyliM5g+TUlcf7/71UQgV37cyb
puOXUO3eGJ7SZa7t/D9JIM2cDctjdB0xukTp794DU7PvYArvwY8kkHkIOtuF8avCYqkKPdIXaz9b
p3ztI7NK8vf6ZCNEYUWhncnHJXXfuzQX8fDeWqlYzKaZ1wdqSXFQHMPBEl/LZMZz/JFkJjP2Dw7Y
PH/W8VOv4Uum4jDY6tqt0Mlpg0Lt+DH2YU52ipLit3l5ieU32Bj1XwLRDHEGipaosvM5NwKk/Tm7
C7SjxoNM7y4s89G/q13JbwKW4vasgaIeMClvZ+hoxfEhBBTVHMm6ndrVjIGDhFKc1ysQZu7Olbdi
GO9egn4tIqLmiqdt5j60e3okJnSMzxK8EU49W1wr7NqpXmSsTYGHBM9+/SbKUYP8/X7oHU4KN0KH
lM14JrEeGP4e4YM6pwf1qWDJyPR8/BLEGAvF2gdqu/HGAm6HGs+RDr1hTtnYEizytphoYXWRb9WR
8CuAjip9zpCQgfvTJPi/faNk3BVm/HRKTWv7rQkSU2yQdfd5XQzqWvnrx+uE+OFIgZWGoVaNdNWv
oUwkpdY+N07zcKNfxTz9j5lEeCB6/QI24jBdrs71oIjCqkR1ruy71hEG2AjPbVdfTTCGWfR6cfZo
CP/i9sn0bkygIxwSvj4ODcIskrpFC2somUujYVVRaA2UP/FYk3ecTui7Y7Nqj4KYrO5fV+x0KdzE
URUjybIZ0tigsfyaCtN+ZJAf8B6fQ/xEuOre7DYeN3DCvoQ+1VhST5Su9XFIe8wJF2YLB3jTMt1r
Mz+epq989iPhkFKK8J2Fx2yC1SxyS3S9oYQl6UMVhrgCpi12u8/y8fmBuwvF+sw/rgU1PplYzSA3
iCf7DnFnZozuOUypJOKk9tdyYHUOAPyVrYvxBtmi0McLJOBoxL1+ZIMu36Qi8s+TucwmT/d1cWy2
2hSTzOezj7MeCcNWsxFEEJ893G3AjQIiodCVNEHprz4bAYOaEQc+4QzwX9aO9q9ohJo0/tf5WDvU
zYZztKe8di1iLvMhT47ubOqPc//Ftejo6s/nFhYe0b2ZONxVh5qyk0KlEXI/VhlZOsiR8n0GydYk
qG3BcydLhxvjl9Zk95YcvRzcGbPBGhEchXtmCb28obfxu4QxoAiDKufN0nVYgK2kEYBnFuBKh0Lk
cRiGkoS+KvBkYggdnwxSQ+wxEcotlUwHvXIyMCCDxTJVsQYFuVOxjWESGPUPog258h1BnWKrWCmp
QnbBL4zENvZTBsV9gROesJ5Kam3fGBErVfVKQQHYljYx2GC8TpkJydWsTDFroVBo4+5+V3KhXCkF
ddCUmfZZiElHoLAhp9xiF4uXc12d0VzEYtnNI9aGCesIgMHju5rQpCVZRUURRvHZP2tj0QzF7x/I
yNvThlGTzYz0hpXLY/bme1e+tyNeIldNScNtamCHV5RS4J/DU0uzzBdr3N5byszUClabvGVubkGk
1GSfqWGzMjXiAJ2zEdM1c+sfI0PcwHSbONoOhXIUkYSdevjsskN2IhCCkRWkp3xF+EnNatXPLFel
ASWNxSL0JxUWAjccrtVfhKZDS6b5BKRp47x0Kl/g6KpnsgZBz1Ac0ce8qgfG9iesdwbKibpwV6GZ
HuqBY/tR+B0OG2FcRvkqS/3vuM5qo9LrpV38F8IIiZbQcZr9VYQ1tZbgm1QnKEqX6v0mhNWVR0C0
4OLMZSxQ1BIVOckA/JJr40yYzuRfIcX65NAW+sM2ercCM+IhbqIxltsL0z5m4AJqx3BTfRu5mjue
ULSPEcMyohZiuNsaGwv6cKuEiATNGHBslOyEs9USqZKMhW4xn+oittfsIwOVv7uqMbRAgGKO712B
GDhkHEamB4lRJcgr4B40AekjyZAEXUFU+MiOCoPMxvurA3E7oSGpgbJF9fI4gD32WQTw7UAYoqaF
a6s1Q/GsZY8OoVZTjPOZBZfr1VNOGR/67bPvEgAeO/l4bpsUvVCFaDCMD8ScwoPsSveKaeAr4Z6b
fxXUdo1qEVkRgPmUfbKyK3K+/4h0cwMiKc5TPHfu1cA9Fyw4+Ads1i+LJK8ZpZ1PBjl4ZYlxpF1V
bjCQoM17lbhIkFUzLomTdsz0xIjolDOspJIsPuXV/2k0IfyInxd0ScNEjUCn+/de2zAOruMB4+Cc
4464EsrMSzQBZ0/9X3Z921VpIl6wnMM6NzsEYxiP+lw7ZjafhnxcRXtuGBveF6caZ3dKDkpx+liX
zvULdrHr9q8+0Hq8GghQPo1ODeUDKkR1bMhCcpT91Cg5OKPvFiueW3w8inPfUZl37Ao2g0E3O6ll
tcm6dja8oN5peZuacWB1xEAWHkjcWWUvM4ddHt5JdE0ce8Rm8fiw9K5It11IvwvPESUKTW9Xa0vD
yusk8ry764JEnopKU8HTvieyfyVwru8vuK7Oizhb5gNwOVczjbsFx0LJb3sFoE0XfRKuz+vQ67yc
V0euU6qWma1Dj+I/jtCnQO2nve91FycxI/g1XOPuMdH9fG8gOXXKdt0WjPymaDDue5Dy9vKnkYNE
BitlfIMPgbTDEDgcd6y8k3ubVeJGonxSojSk5B/5b0YL9BvHG6LqLGDzuW7DKzCgp5if8hoFL4xP
Rg8K+uQpg6aT4KjIVuOGqgA6Drjn+o6PPjUChIggIvc0cO1VENdOZin2l5WIVXw6YEbJpxtyl0Ai
jUuSRhmjveFVzArgsUt1NNt0zphIrb/VDLt5eLLsOI0vtdr9IgqozHNGrhH/3vf88LeYe7itORui
Aw5PVOPeBCCXgynR+fXTZ6//aAswJWB5uk84wjpzNrfOZUG9mR8rlP05K39jR4ZMMdUpgEGikmTL
tb27/K4lI4w9/5QDoeZ/8g+6hEWdhFxsaExMtWjESSj6f84rACA8GzBANIwjscoT4hEQ5sfDSLXs
IhadmYSx2dAIn0baC7E9FNvhbVRVpDnLkizQoqMiXepDw9Ow8THccKzsSps+AxPBEhhETUY1heOq
sW7cYJkVMbVG5Cs47BgRjopeZNtHP9sxFnShifGKBeFEYNBmHFpNrQVr/MXRfk23Vx58NN8AMEGH
mJgj4WiU24HV49oFMvU0oqKf74hQAH2mP3eF7hsj0I50F0/6s33BH2O8yq5CHVeZGZI0lzBKY9Ke
kASPomwTcug4TLd0KMsZvoehF4InHfLZ4YpeOn8yAAxXy9SO1+2EisZ7vS9m1EXNp4i3M4FeQ8sj
5DyV3CRr3AE0xkrGZ5UuW+z4A8Bl4trMhkwV70p1zRYc6H2xYvD1pIlyVOuDSfi0gLWDuIZ7SYlq
NtwiTiAPIm2cZmbpf4vlVwFT//R6+wgoOJrDctGvRXYhoa26/e1wI8lFFb/QTKjZFsYbxUiZEiTZ
s/zCSST6hZ1kuRnmNgu26MhSL0mXZfB+BJXWuNItwIhVfbrAUtzJaFpz/L6RM1FcVMrJdpPX/1K7
xpWAp51YUqZ/AvbxZxbDb8W/ZRpbO3vKOOvd5P6NChXGOd+agjdH+Pe80pYMCeXNYbv082qV0aEo
Gt7BElKI7xs5N7cXq+tC/EY7hnXeMcHdF9urIkgC71nH1OabU47TkRAKkHFIs+7YrUvhtMEENjKV
iM7ltu1GrtEwjgwB+rUAcfalXVcVyByRkq8mkJFJEMqBzAElS+ObexWvWkN4QbgyCMt8MrJv5YgV
umyqWm5orU1FOVHIdIeV//G1+JIOz30ToFSqNJLhwnjU/eeOV9o5riEX+zNdBFomoZ6jp4Ot/euF
n9y/68P69ec5FCV9aFyOUL4H+KmYOcbOqJpBgTTVG9jwdTZTePwOYeWpw8CWAlMY0V0A7GYs3nHz
ff/192AGm8+Uzca4Yl7knfrMet3Q3FTIleDI7ts0JMCLzV5SvehkvfAkMhvS6P4Gm0yzvVp0FKAY
xtHySEuUIvKiZFc6MEsfhAz2bzhb1tGLM7jnRA99ryR01do2kZ41EaKUpBaJraMSLbzfkiffStYB
ACNy1Js0eLxaDg43AEcC0p8KXK3+8hXxx0pX2n0Mwgv5lBmDZHQicmfH4I8ZNo6AYulsmZtVWX6q
gVMQoyC4IjflP6QILGXhYrxHZCATmauunNtAvl+eun4iEXo05HVTcxSIC3y2VtwMWnyoxrQVtYEZ
LzwNB5GAC24KR1HVSPz+I41pl6oxwsUfcBJaQmkFlkdOKxzIYlqFXf1XownCOt1xpVZIHGeMirZr
bkiLS3GsoK5pLViCmm+48vlL+Bah5dXuusCMfZFI+4GUXKWV93c/aKkLfO3T0+ylInzCUHnDBw6W
3py7FM4oPxype7ZmXw0iH5rpcCz9wzdRaCWfAGHpq12CRHreB+LJZKwr5w4HUkWALfDrlyytMLoq
veTzcXunLhPULABhCzdhSoEiLvXRWo4lRuAjBcU2ptEvGug78oRO7mL2Qv/jOUIb7jA7sP09fSlp
Jkz2JYIzyCRdieAiHJ+sOVhUcTuji0UgbqPOpYZAWW6EV/Vc1c/uwl8wds6VzKMOl+bS3/ERlw4e
VODxv5dJQhCK0Dq773PHweM/qpQEnqqmK5AZp1VjDNooPopPVqcVEPjhNhCnJpu7L7z3zQ0OqxwH
rwdrHFJT093SE5ZUWrk/I3VCgFHd/5p0JsojXAs/1ejzYvc0FeAPLxiY6E52iE42jdPnodr4XVry
ghstJC4pz6VG3mEMPc+oZ2i+y6OsOK6K8V0X3T6qLz3svfZoWL9la7lt/1Mr1aqIT3pwO/cv3yLS
SS7wi90EE6WTGeXMaY/1Lz2H2bCgwQ0L103Jag8owOVf9chnSlx8fRb+VtkghGWuUTDcgYQE2bZC
lN9aqjHu17kBoj2exsUQowfqfVgEY6UAOTrJeMzXHSoDMcFkFWcNo3bZW0XbpEp+u7I1Lib+wk7C
orSi2FsHguadRBZXEQZBrsgJdW3Zi7Wdge355LecCgshJWpc8E0yQgZVydz61O45u8wmVMV/FPFu
fAOCjzNq0WQdxwV/guSOyaTB2w7e/s53ybvSHQ4l5TsO/A6bUg64EQCeznh06vqUzvwvk2DgrvCH
qsqCB6Ia5+885Vr3Kf1uyRs7BGW+IFazC++I6/1CljjzP5ohoiMC5nsrMPGdw65PWsLSa7krCV4J
sTffDHU3F+fqsqdMwHWw/Hnd/ndsFm99ImhKxavA/bJZY+INAKF2YMIAj2PLWfFTl+K+ONjZackU
7VLybGt1Vku5DDmFTYks5dyPbgAJr4MX+8HR4qE5zcbY0KA/spXyx9O0i8zzzdXSr4hbAs2pw+33
FZ/TkldIjFDj6U4MPvSg4BaN5Fy10pPV3iURBdqv1OxV8/yn30cnOTHEl/kNnbf0xSQO5D9u8syK
faXg4nedAddyFfpzDaSaKEllBWkFmFnEP9Jxr42iYCTEbSQRiYS+S6EU2lPT/uv6au6g6faeV2cz
k1zL8baBp7qVsUZefCoKy17yupYimurSh5SBr58SucdiPCrd2mIGXi6RFA6EMMSFKr+mY9XVAFyD
FjdvQkBu6LGSiEQ7k1ZpNZtQ8Iur+ZzJlMKXhtVqYEIMiKqGwOQUI6m/JgwZkpIXufVw50mJLhDs
Oh+34zfwWww1BBPO5oHzo6dFE67QsvQkJtJuSBtp0+C3QRh6qhaN3945ktm4EGWn1jAYpElqhTFt
xsfqcW3k6yYRB+daLIZ2lNx/j6kV+pszO01hZCHYeY8h7yITmdKfNMFsr497g/2OLcgV4yPy9smq
UTAkTiayqJt99UXVyrd12W15djrIgQdjD5P5c1NK/dxHA5zMWuHV7TaxmySmocVW6xmBwL9dGjYL
W1I/nKuKUxRbuEPQ68TXA+snuwC+5xEGt3O/7XoUT8gWI1cZDnka+XqDDTVEIfa2nMheDCQzMleg
uIQ9yBWokJyMwxYjQzapkC7yshykg20fVBqwvz6gnCY0mQhd+DN8mjyMGBoyPLhgOySgeIepK1fm
2zi8v4mW/277q72jkLxtOIuVa8gPLU2RgrBNdMR8dlSDI6zwoMLnkfvD9JAtyWYPj/aEsPnBQJ9Z
H2Uwitf4bZpJvI91gn2VeKXnL1lpcseCfcyf3TkQPS+A9M7Pj+4nHN2EPM6atWoESSGgWcERrnPF
wkXOJtDKOQ4dhLMfkdhsSQKlg4g0z8yUGqgiL6ixxq7LVyAT1Ca1VmSRHzZfHwfobDtDBNNJ8R0g
z/WY+hKKROVBnkKwCUmwTSWgoyVU8S7C7b0FC6mLGTm87j40FTnbDjz0Bq+6j3/BPY6a01IMHEzI
t3d50cJZ/hjzvcHKe74bbFG9gMkKzRNVLgm8zva1VvzE9Djeg/El1DvNu4Mvk8F0vihHtPdaA68Y
qEfQ5nt0pruJnPUdCz4HtE5bXUkIFx+MlOcbtBPX6mTqUZNJ4umHrpWmVDRPOEVurG9/i0liPurJ
ZFMAQTSz5fmMLFos+/pChR0RLIqW/hAj+PgtkF7KNxkyLjIg2u4dLsZ1L+Gild0rOP8Pzu/JoFpl
7s7ViTQmuhaESG0OC1Gyv3Dct/5psvhQjAXfmyc3GrOlY+ND6wvT0724/f/pl9Crd0F7Z/tUH7iL
wj1mjbKaMZFDbOmeWLVEWlwXyYBb53cVPDP1OI8LMlBxj5Q1lBZ/pkP/be6DXkIm0S17QVQVw4wm
A1JUElUjJ4Mty0rW7qBA7p3lSGtTx44VwoTF0ry7Eq/y3Rc5UEBjMk+2o9EjiqjiwmwUC8T/QsjO
4c2Fmr7bu3AWRmIL0oOE/X0PBox9mLuL6MAVmd0hf8/DRq6V+jwIS3sj+egkd0aMcoeIMTr16Xbb
I2a1zOTvDJbkQI2pXlqpHsm3NczDLRFLED23hdKkBVsPnkAfQarqNnC29a0NhvsRzfDi5QXGxcbK
uWBZOYmvCwccMZHg1cwV0cCi/wv3OBNcqSAsjysMub7rVmE+fHPVbyTWVrIEG3LZK76TQacx/PUW
4nToIycfEINzWPEG/DZ/paBdM2KuddbB0ewFdzyY+eGCAg2PMoAYe4DC4H7GcYzbyY3c+FvnCWEi
KkHVQlODa0RcSsnMUgiRhuiMoOhBNOzQA+bPrI9KcrLAqmIT/W9IO17n/UR85aGp9WWsbi9Ex6eB
To9SGAkPtj6A6IeCe6oSU88YRLLFjTTAPznF1ZciGHZMQBCyYlQuq3xG+h7kJqjY8xkEnhHcmYYM
kspWiUkwMpFvqoLZUHaNsGDvX+3fikh+0C3Z84VdgY8frwG/PeMSF27Tc/oOHiI2IqRGws2xswwG
MWZv9X74FyFZpyElZ/fDisGfWDUYBlcvfiEv12UclIbEayYWKPkvH1quVOr3rSLLXC1sNb9P3Xn4
y+1Tq40n2NwCksmXRJJMwfb9TNedmYmYzSk4uRij23KmQ2hOXk+j+FChEYpKQVljCqrGauDhfeS9
5oLxL6EcBUiUJvGEXwyySfKLti7ZuL83FH0cW/BlvSYp80svUrfZRFhdIxf9IZR9I+kaObxOR8Au
QqzLVzjEVsIaVEQFgJcykoKGPlX9kcYd6N+OUybhn/nCQ4UQQ0fPUlxPHiM+bPCm09VdMN3RJy5r
Zzn2Hmy+fjYA8FOXeeGmtOI5VlRNO1pE6yIYqsUhk70szreQvphsHRuGeO6n86ReS02xDUxERoph
VFnRhwFVlTfNTbwpjMYHRmYZYs0KH9lucApUHcEvhjeJFXMtgSFaU8fvU9VA5QTxG1BUJffHBQLr
ra8Q29gHQpU/pxds5rLHvCitQ4InEkJTBX9c5IF6J7eQrXJX3gECKO5894xoYbGGXXz9Jx992Eay
gypGzh0iBDxf3v6zrliJYNuipnSvH7oM2oJmoXF+ieAUoTQ2CJ40kesJXAYklYujIZzf7gUWkcmO
m7AP1AU7CvullrlQIHfv53ieNUCH3/wZW1cQGOl6JIsIfFDmb4+1nktXiNXiOIDK/L2n3vkSPL+k
Abj4ZH8vF7V4Y94MhbZqoFx5tfJ8SctfH3DjGIYp/c2hyqn3qhHAogh2/1qpcOskqWRlgETA7ind
TPnPRalR5BFkmYSYcbVBr0Emf0C0/0iY2lXOHxppbXHiSDyNBsFmlfaysoRqtNUd/sxVx6NeR5Sv
7KI+DXkxFL9MPg3PDEQei2hgc8W6Wya+t1Z8hnkpXh+fJC6PHBnSrii0+6ZC0U6XlBMDS907FwKQ
lpzQ2XOv65beYr/jPa2fqhg7xx6akzpW4bVaWZl4GiTxlzLe2Asl5x1tlP8CdvGh9HSCvX1HbyRD
2k1MSbd4sxuKpqVSXOqQqR7QCPAKOnayPXVxwpJBedcCa0ubIUN5Upla9nMZJoqSk+ciTe5Ofo8E
PdDPra0CmEAP5ERcQ8JocLbqE5JtxdIa6y5cRvLhKVB/hZq+aKTpzps7zOY8r717sL5jAaBOS73y
jnIVoBcn6pgTzSHj+Kvt315xiRJ3ub5RDG/4YFdFFUPk/zdqAqjt9vCFriFLiEShkdGpCiH1ongj
SoxfgpITLeU6g+9Mv4MpK50gKS7hGVwfRwPdwFn+gdVYVjCUQw28T4M8YksAjMkRasF2oo+E9YwW
UZh64Gg5grVtAu66Qdx2laAvt5xPuB5tcq+yTcj8Hhpz4H9L9AnuUUBabZPCOCEnadvCKV2Sdqcl
ZYDR0rxJyL9PStpuRnB6/HVFQopABuM0JWkliEfnNe1/7oPiOmDctH1H0r5Fiu9DrH9TiXVnl8Tb
oc0xKMQFpd5IAFPOfrFIxDeGW4j8+UPbMaUS7/03kGoRqbK+yqxGwKVYYOzfByu7s8UYtI47GeLc
eN7VWm3JVRTTz1P+OX0otpgwgQdJoCVQjrOZif1ZWDQ0ynkLJDQFEZDpbh8WFubVq3VID6FoCpx3
8N7GYVm4U+MtFLN01X4Y0mA93n0crR5x3ScCu3YycD4Gno++lgMVi60vfCL2bm+hJW+v8DrKNz2e
Aqg4j0CNeU6FSOkfaRnbVmDoEKlMbFzBmrtCtuPe2HD/2bLvq4toc9V7yutK8aTwAAXrzAmhqDNp
IEY7vTVQZfSFa7OhMTq+kDvTLZm98jhpsMWPT9WVOcVhtlb/T5IYuLKR9MtRoqEoQMiBfH6sn8ny
RgvPIdBtJCs6Qp4F5fGQl1iTW2TpvjCeW2gAaf3cOnYBYe0u5f59I3DDHh3D+Rzei8p8BDsYF6NJ
ZxGXhqjOCTCueAZ+pMGnhHwuYyG9AoTFmvejfx0yzT3uMFNwfoDNBeIHG2/3AI3sG6gim7KOatX6
gQmY44h5qclkpk4YQvZdF5rZLT9cxMnGQhz2bq9bRx66X+ykp5sgbh3pP0h4U+XuTvgMGdlqp1bT
0JZfEsCPkvnjDtuYqWoxmad8G1cVMWq+rZacbBW7H29Kvm6YuZ3AqtBWQdhG6x8h72GJVYyEFTNF
UFgkWDkb/bZIOnGHbGx7oYRnh92mD0ojQ6rhhq0w6/3bRhAsmg5r332Cb7BiWRBmSs3iJe2QD5Cu
UsQ1kcLnmALAhq+Vu7Iy6q5aJ/k5cwC9Gjk1CAv7lF3aUqFn5XKkKBC6dwi1aKGgR8wqNhwB+U9i
JMLTRnYXj9RvbxleQlIJErWt4R/XvogYLnsfpMkSZUbhqJm8gm6ke4Ut5FpnHr5HknQaT9MEkMF3
0dHs3DBVyoZklt178v3Wy13tVDNmJ9Z/JE/QnTlNoaZi675S/x8UQ7aXOWYJPRXjw0dNToNg2kFj
k/pdMJ15+fzZG5j757AaxuBe0D9w57QPbs847H3l9rjmjNQormyY4efRFE44l3GzriYDSPwbjPqR
WtR0CMj6zYN54GALoMEyXFvs/89Y8RVoJt39lQ9yQGthot3ABOWMgj0thxo99YRHHtf6D75+SNGY
oSAk/TqsBijPBY3B9iXSUBaJWqTq+lJ3hjdYLKCcjdDRY7ZH+w14feD/o4mu9/RcA93H8wu73EHf
B0SJS3f+Gsei+gVxSSWQKxN62cmjSUxDH4reNnPK2hZaKzWVd1snZUMrC17XSl1BuvAXTBhevsPJ
ZaoTTEZCWYVkOdY7PTsapp6okm+TnpeLGzisWWNiLOoaV6SFol4oNZ5zECCaIuiQo/7F4ucH9Gx/
6eau98CbpZYaglr3KohiOJVJnuRCXnlx6dGrzM9lD2GVjBvWqpm5wDAi3M1LpGFl5BmLFOD3rq6p
PC+EYnwQi+DweoE7e4ZXIciZQbbwMdAjSgfN56C0SKcmCUoFgETfnZQAYieMwhvFjmymMunuhsmp
PNNPQ+wwEwmi8WyjKncg/P5Fu7+nPHIQcOo5PT7W5wCpo3k+nlqbZANjKvJk57+BzuwvOw3cx2MH
aiieTTImvxLLyWUy2PtMw03xXa2XKqVkiJD4Ft8MgUBh7B0gUrBJSddfRra2QBvF/FmGWZCOhhgr
NMUFeowKoL9OsAxj8Q9wWyYN6qVgjDBaJeOY74dfYhnzJolpSJUV3eY5kZfHvYeI0GReCXGKaoS9
zMgSdUGjJRyJ/cGw8r4mN66U/TKNrLVTNxdK4kFjOAEPN0BGJkmJ3FO0mRHJdRSQfEzfneKaKMEo
6P/274zob9pAmx/MrAHvQRFptYKcVAjxYHz/ArVtR/B1mtkhGmtO1bXQNLYY3V+j+QYaSOb+2KuU
qgwekCInEKZRxUH0VKncCVkf8M/4zC6mKemmkv/H84M+6r6lsRF6n8RfJD225zBNFIVSoviYSEQs
lAyumpQk/YH7dC/IKUYBw97aID/yZ4iK+ta/05kkcJcWjAQ/X9FbSoHMp+tegY9JDuGxda6cZ6eC
YB0AoZT50Yph3eOSqGmDR8PKlhLcMqChLh6uaG24YgcC09B2axyhpSefl9GwVe3b8q6/cvEtlIme
exrA7kOCqVAlgmiMkGbmrupgZ8KKFWTd5Kyq/zsKqZAD6r2c5jc0W44/vva42jW7o33CaiCGpmb0
m6zp1eL/rhJrstNEZINhcEsk08shTSng0K1f0BXrIo39vxNXIJ/0zaU6WvcJGNxVrwq3v73770iv
lOPFPfQH0SSEqMmsLNMUPJ33ysRc5qj6yD9QNLw5+IypCy9M7Wsaom70PDufMz1fy+E7Rv8DtLHj
1fvouO5cHwmKiD+JCqyV8ZAxoKmuhMTVrso9SfKr6qRujRwmzAHSZCK6dVsZJpgDkSI4fAL4+NMb
PBKmt+ZMAEcsDx+NV/9bo6Ir03hCOEjOQPTB5serMhqjpm4x7zlSXxI8JuTBctE80W35IkpnYaws
DJLl1MPuvQRHIWslMZ0Na+QDGSetA4DcBtsD+ngIwb3CjwecalO1961niqnlxNRfm60vd6/ZPBWD
W4owwdMKPR4CJBxfwxb+Lg9S4VusyciCOu2PteveY0F0aecdBp9snjxorBi+etN78iLwqY2MWd3L
bPQjHv91/KW9gNQQi3ZwK6mjczUsOSIqCmaPrI1JtfWMWNZzYxmoXzRVcHjWaGLMSXPlJ5LJ6PME
1m5hLI3bqP9mp6XHDJkwh8z9FlX+34ATmjhf52RzMDv44j56j5l5pAelVgeFxCZGfUvhaEo9b/Nw
3lZnwqF1+G8n1584Ndh15jZYh4sEesP8TM5ymujo06ZNhVXOY8AW38TMU+4Bqc6QYQr3ZwnBJZAp
5mzJKxKvnGr5jcRsV2jjcG2+RC0PtnB9NvPYyYHyD2DL5EQcRsum7Q8MbOyULeiR/5WJYmAZTeiB
Nh3mzeVpRcjpxmf069d5VvcfNhEpHD9RoDqdMIaBqFXp5wX943LePk25H6wS3D3+Lc1T7tStSGv2
XRuwPfuy9GCWB3jbn5SzvsqDmdUUaWLvtHFahUGBrO46i3zVrkb+gaAZU8V797t3TxVTarPaBv8v
f7LvlwPc63rohp1PgMiM7JagY1a9pOUtk07jUXgPhZD2I4fJsYsrt9YHi2WOsodycnQcqX/Weyce
SoGStb760jfjyVd3tjPdGbkJZgdgDzJ4f3/fNE/fxBu+1igNTNEjUag3zKzA67MDxfgpuEF6rNqf
ausvvWybYlpCu90J2A/f2V3m+MPhgVKqh97wUEBDuysCdUtcK7045RPXy50EJ+rPt5sDh6bue5Iu
3cQ9Y0eZl4DzsAvOqGX2jmnBoEqb9eqJjPPZSeaTepd/cVdYiIeHyJundpUf/GNXvsXVY28ZMCqI
muVPUvJheXpHvOagCNghrdfeZXYcJSuEP1+dJR0rWxhkD5tFIq5Kk/ELINh78WxNnO309oVW5NXp
1upUg6+aWFYUREx49JnMqB7juRv2ebpgzFoXj1vSteJjxLmKtFZq1aoE8pvuhmdiy0zEsl2iCVZf
m9gFPmdnPEBKzJb444EDgcii2zixYSyhY3MariobYlW/2wGS6vFigE8Eer71RXHOuFBZUvEgyRp5
lSTTJTzrhaiFkvnl0wQRhoV+KQGGi+C2m51vyAz3F7sxR8vEEZf2Jwg8mwa5rN/JeF7Sapu/Vuzz
EL2b9QS0HpnEFyaLtruAafF0HsGPgpgSmeh8u1zni1RAPmQyCzF3NyaNb4BfEQGqBDZwBlONIC0s
wYbQEDGOdReggi74cgdNgTEI/NyS7ngbOx1I1LnyuQB55aeuWHZ1KzX8blMcVSCo559xfbUZDCxD
KZ2HtPt1Y0cqWPcEx+zLYcuXeFqRMANvZ/deJjQ8dhALKoeY6xtm0aSpQHPTonlhx28L1fXs7rDg
RcRY5VCfvLR+VGI7JfSSeyfOJ6zmRdoPdtqzmarCO+U2zzQvDi/S3XBpzNgthwHyiahrfEIgkheQ
j/Yf4hpjRpYfn9qgqwNyGmaD9iwmo07BVt1Xx1vNvv/pvO/hJeAx19WRxi896TodQGd1RhWTZJUN
+va6bmJcbc15oL0JAawnJp7jz8lZFjLoukGK+q98Ejx0bbY2NGSiIGH0aw8soavT7HKcyxQy5LIV
ad6iDYE3VcxNQNs4Y50EdNDfSC7Km8br8ffVJfw/K+M+O+c5nMBUw3Kt0ZuRyFGGF3MRO5KXxKlr
drh3IHELJOqWT+fuJ4d1rfswUjli/TYuxlS+29+1djyZ2ADIFQsxAP2CDUi1+kAehyBxXu1O0oXY
cQzLkL2hJtO4zG+jk8KBTE8VVnEx5XyG42zOSjJxSfKNbeHVCif8scSiTx3cStnokTaDCs5suihn
6ZxxUFgKx5FxmX26ej/yF8tPDkqOiU750m7h+Yr2okOI/zlxXYNGl8vZqqXSDX77saCcCvtSa1KJ
+EM0vS9bnV1Cmr0g77CvNmhIf/AMwwwPItS731YRFXJBswCrJisvD6xSHGEUUlmLwcTjGusnpJXT
lk9zLFVkrC1ORVyAJaWc6XZ2Yyv29WsAoyVPOF6gZNm3DEQ/FVanl3IKuI9qV7UHkY9k0w6/auFm
X7+Sb1NCaYB714tmE/N1VL3dFA8CgaWHHPQ+qw5XdOiJR2K3H96UxXiFDhmln00pw1iKjR3OO++U
N6puAM7A3JGVB1LD7JPWOmFW5r9dWWNJXmfzC+l1McA8wFu06fe7WcHadZnwLxh/i0lkdJMGuwsP
jUaLWI7DkwRwKf5MIYFtBS4lf9D+6BHX5jlKrfyOW+lVUnrA6hsreYkskjz6VasNUZSkBS3svEzO
B0DIel+1vejvxX5pvjHPotgNAtTUe6cJkDExR+zO/Vbe9iwvza6jkPBTFcmPxvtUEqLPvN/NXBgm
R9aHb+2Lam4qAM3XK6Iq/tteIxQLcGmuJ0ZzlazW9Kr7e8CZj4GEmIkdujmgBqSz9yJ16hXzXWaL
Tp7gwV74oRpCmvwQ+aHDoCk0kYC0vBur2IyrXj+iqjDhjpemJHFP2uPEtwqthCrtj9aHZKCTEwRT
L5ege6n+gIbA9XHJc2sLr/UvYr67t+VNWvcN+G1FoNv0S5r2/cO9u7Or5SOe8/lz06KFxZVk5xbn
RE3St1JCLQ9tA+WovLfTht0tm94Svs6idlWQgujzg/kS8JkX22Ncnr4PhuhLWeJd7TKEohxOSumr
MtU6Sq3J/NNocRtxeokG0Gi5Jf6DHabeK6hrTLhKhgMjiLKojBgn0up4MQJ0VlPiDp+s9QNXMbLX
ZU+0bW8hOj5inQdbBiPtBX5uJ2u9VqwI0w220rr6+ru7q1Tmch8aup3Fv570R0fDGMAXwRvOFI/R
FQwj0KjR+e8w9BzlavDXzO49bTNuokpfbPPZ39eB0UAUKzbk1YmBm3xogAVl/iWWVFA+uj/n/wCT
3i3CpTgtPw/JPGkzCA8BrKz+gLWyQm8XhYQg1hJosYAnT1aHsBa6dSzXX/6Omsn2dGLkqU6+LK1O
ghaJGbUuDifJ5Vj4fQNW53tBraLXS24tRyAMQGMdrn39YfzdvV/tHOhDhtA13BeziIwm0UjU5Oac
2ufi8CoICtG63c6r2MTB4ym6nLyuvM1mjJeHJqSoumBJ0KldLgsM6pt5N5Y/E/hkJFTGLPW+hMNk
+2YqorY9J/RAi1yqIZ+1xXp8pcPIDUovMUO3pPWphWylVnXpk1XIpjg1i3iXQdY+Wex1fFZgV4Hi
la525WRuFjxvIo4Tn2H9FPRP1De5ZZGKkyvribTC5NMX3GDE6gAmP5JW1Dzy/S5nx4BXQAthLiWv
LXAN8JUZ4wXJ1vqJMdGzUUVVRef36sF/H2lhdDye4pA1UJmpmCjs7U1qDrqVpjauIaanCPOAqKKF
++K/IGl0xXpekH7lOoGb66ZmximuQkVaVrv2OsDl6AMDatuOu3VJ/TZWoLyV7yXlrIMnyci0pr2N
Os6ymKRDG9mUkoiVEdgRnp05WIb9fj4GjUwQLb7B26C3LchQ/ULO6wmv1DeHNnVasaxUnN1JBSee
d9Sn/AkW/qdFgifK8r/cuqLjwR0/P1czv+uU6nwiCljvms4yjFFixbrnWRtyNlVdU5KTJo1Q1XA+
baiNuWW5FwMzmWZmIVc2Ag/TQ+JTPaOiYE0jtCAWMvf00yDqJc+s0f28Iq2vpE/Dov03qKgk2xCr
LDBJYr2yoNqjZrZFBm00nHSPT0+yKw5atbs8apqz748yrR1N8+W7orEObBeM9ww6473o8TnGbBbI
ROA5u385PjkFn6tW871aWB0yHTPGHNRt/2kxHGBEWclo2vlmCpObfzEfe6JqBkQ76l6KSsOZlRYG
REvZTtrMcpNzPR2D9mwnAm07OsgzX5EgJPhiiHg8F8T2AIhd5KGXDBExn+cl9sPZA4pmZtQcUufv
mNGYM7RR2jYZoWvM6s6NAGoWqZEcRGcumFmpawbt7ffbHzsNRPoMIKUPLoZ9VaIi8osOZAAIM5lr
zNHlCdJKPvQyBdx8XQKJ7TtulucPLOzwYkG/X02uySCc32T8iWieMJcKyBQdxFBrEctopyvFkS3i
dP4dXHR1J3kj/Npk6kSmNs6z1mSet6KKJakfRSvesZaN/BRySULu8nncI1E6F05smYQQVynliSLr
JzOwQhKX1hoRl2GOAInnA6FFi1gNIVHHDRlRPBxKsZVB5jh7GpLnWFONwcf/MBlw44pVP8mttUJt
HdAIZUda+tOT/tajeG9xcR/mxkg7rjCz486owFyJatmKwAKEirnN7OcEhggmXyJ2VPrJPVJs7nL8
cteplachmul9sI/0GTEIq4YGXePiD1J8l7SM+oq1aPhwxmlXNOvGyVUlAM16h9P9Vi7c8oKXXDfh
9c/DVsEdDr4sMWT7xYCMD6XJ9p347eKYrrK3/uF313z9Udp3EoKtRnPHB21zP75WF1/Yo8tSHjhP
CKMiEXoezKLXQgVUMQZjYtfikvAMpSbx9CuI6N1yBMkBovo8Ja3aqTdhU+fkvRJmPx6L+S4jQZJh
AHIAqh4QlJObZ0CFXzptXuzu89sE20aAC2i2DphoVmkyTlPTnfkuEExZgjcOGxNQiSkOzcloVcmp
OnuFJtItHJDVs5PPjNaP2WcDFoDujzDnal/Y9KnTXiy2fX0R4GM7gq2aB1H9+0b0up8Qq26JUyvY
V03eRkzwFkYi9cNegA3GRzc9fN+qfFPXlRva8osvYYeinX24NDy62aYwCmM9X1M23cSDZvHTFGVC
R+7VgYueLrefiw1yfJVOEcIMOaVr12tWGNEoLgK9h/3Tm5kDwq5wW1dvlrKgAenkIFskGy9JZ6GE
cEbyTZPMtCe9TD/Xjz8V5lCzYIVehQnJ0gpJ+XLgZhMq/NpPAdlbj4nq2ax5ABdDUIJov/+UZzNr
rtbFKvqqK4v3sKazDEsU0hE8mHhaR17swoaLokrO3BEoWc3ZFM265+xeIHHpIxTtR4xpTZii+7ku
DbIfXO7zZm+RSP9KUDtrkz7/EKAIx7pNmegFuI9y30cipsGCrQpxNhe4ML5wEKj7nUCHHABcW85r
EJFPA2gCuiVATGRq8jQJm9Qy7M5l/70lx1+y78TkEmIR3eWqdGqjCzcg1z+fRmKSqYlm6QaFdbZt
V4gcV5WyEkz/e33q9TBB8C1/t8fBTo9rVxcj7zwFvM6wbniN7Xr1EEgaBjcwR4s1p/902jFbd5WR
kAp77w/I3swUrIFnehVoNQbzy5o1KwmWts5VC2Ns4qd7+MYj3j+THVGaMUi9Q170k4r50ZU8xSHA
xYLZb7E0tnGHhlKVtGsnUsuCq3+rXWdnx9xtDKA1yz1bWIzPiyRXx/nXWTQ+4FLG0fpBflDFu/g5
AeKkRX93GmttQiNu4HOrBqQ3KXVAvfsWc1sjseenqsC7Zt6X24NnSBniyTb/fGj7GlJH7KDnG081
mzmyMliRv6QTEQ6aKyZ5EqK5SBrS4ks4hk3+JN/dNMtI450ohoub/9vjZjeUWCfAJ1K03BZ6kRWb
bz+F3S6qktRytM+SMw4cL/p0+65C6n1GKGKR4/ktJOd+tClheE6Qyw4UkBKZz/GH2dvkxVd1IbkX
jcTLefbeznuBODsKeox5esBn9fA1xT4drEXqw+sUsD0nPsO4jwx/5d0L5fumoitysQgtA2kiKKWa
MMiG4VwxCxV8H5Ty1jNSSn/MJlnp8P0O8kgQCoVgD4WGc1+/aab/PpYOUtIyGKOllotaXtAoTYP3
3awmng4qcln+AuK56DjuBZvsetpc9sBIUed2IASET8PlMTPfLtjF3OXnpqCZ6FnIgTFYjcC30wm6
8KOaZhXtdVeKPc72tKrDUPpaSGKAoSJe8SFUKJUfqQEpqXGGLB17hiSs39ecLkHb+I+s7BV2NxAi
h0WfOPMtCq6fv4CfUf7p6WrBiKLfj2bqJql5PsE3/vVThh7C88SWhyqaBiyuZ1pb1tzerY6ii9GL
Vy6eYaohzX4BHFLUq4sawqORzdU9YdyRZH1GQjtpqlAK0WroNZZoNzj+v+cAqQOa2AS3tOh3OAEY
cBBtKazDfa+bzYz9AgihbGAO7u2WoD3UGW5y3gw3Iw3a+GksjUv5bkz3tS/V1rcyInN47/20Z8Mo
EJipZRkMHaTfZSb5G0kpf/L6G0xOjUY4PsLYnMY3WDeBVuFkZSslrrZpF5d94KuOFEvTwAsbyp7Y
h1Drb7Tz0YCQfxUSRvo6L5sZEyMev3pA/OJkGDvyCBL++O8WMMJKiqQ3186imJZlIVvcX2x/78il
Ca22E/vd1sx92hdn/amQWifn0CS+xKWk7RnJv2okTRTCeY3R8glzsV9vntF9K4BWZ+SYSXA71imr
VQZ2OBTcT1rw8kmXd8p23Pq3uWTvMGhjBLjo0zTu4W3oAc9hxKusl23nDHMCE0rrh2jRIh99/F5G
MoN6iwg0l4z4n6xu9cbJbEMiohlKEdasluJbVLmTYFad5twOR2uHsOy9+4N5W1euOwkpp6Lc4FZh
EqrlNFqSrgGefpUO3kcAygMwJ4TQ8qiIEHflfIUeI7VPTgZ2PxLq7+anVoja0RmiwHitHeeQUzri
wu/P+3pnjAKjyMhWixSL93k7w1bEmajJqyfoN1ynfwY+nL5NegIUfYcr/qaakvp7TVE2MTlRasa8
YaIhcs9fX4dc2z1KaOAb/pgyJ+Z4X/lYN3kHVELAKEZE26+yVnC8H/iiZcsuUhPLZc5udYWTwPrF
xrXrWMSRmpipOblnJveMIH7cfmw6fpdqYeQ1orzYdhOPFew1drFlmniA7XcRlB3R2rdg1NAhsjlv
9tgaVJodfaQXJolsLzKmrj45WCHBpcdjcWc9p5Y4jeLl/zCmeOFXMZ6RKPPHgNMVLFNj/OCb1qAj
tzOSIHeb2OUTVu/I/VwyyVCO7eE4q6PGBSkWSPqMBLY2MFiaAhU0WMQ1q5z5PpQuabeuzcZykRPS
4bC7FDomzetRcIjcCeLm2G1H5lRj6X+aO0qDC2mCF5Mn0Vd5conMfVWQlfcxsP7RFPXYCwQP2LqL
cKqmJ0zRuefqWnBj85gu5ypclvPuDYYUkySHrdASnD5m71CYhUCaCWVSeIbL4izHGTmy8N5Gc7Wm
hdwBCQXeZBD74ZpTudxteoQauYIc1jwccxOEJ9gBS4zLEAO1UoRB5dq8weASgsYACtv80aq6s30x
7TeZA8wcdJ/To3P2CW3HNKvlF7eixlMOdoWZIGrpO+rx+pScnFkw+Na94auNnXDLPd8bCnAdSYjL
uMrTzVIZLF+SoSifEcGFHZ2wASTyDw735hHvuMg0mNKFjfKMiHcrdahENpCKjJqfvcA7+VAHAMW6
IsALqzw2qi98Oc6gvdDACvlyEb27yKqfavrpajB5T7Xh9FxDKWw7VBtZoUibC0+gbsKFqQU8+pjC
+yk7Qjzz+7dOcuPl8e0CEZgXNMOM8RRtbUsFURGxPJJhWXNPOsxhee+cHswfNCfUiuirNI9BRP7f
P+bqR5XBKNdtqcbre04VKFfty/mjUrBg+5iXyaBDxI9HY6IaBdFI0KZ1DMjPSljaMixVDkqfW0sx
DSBeSaYLUn5KqfbMwYf5zYoXt51Vgihz+R7xgAPwc7p66DJgF/IcodaskuiYWriJiVIZ8WiJDzv4
zYv2OC38c8gCzu40DAQs1sdCRksRQHGzO51FCW1PZqdg6JClTjLlwFxK2TpOq7UZaLVVSTLYBvor
7aSBTxZM/2AjUTWR5Zm1TC4i6s7FGoqw6JwiG/DK4LMmBu34RwecWk6oHCvjlKJeuqyi55luXOXr
Js2ejwDfhbsU+LDafAzynhA4xkvK3r8ys2jSaGUPRN0mAVW1R3QWuP4QzFA9KS71L+dgQImNkBmf
FLjgCrrY3my1hHgXwKoNDQZ7HJlvcVCtXpBXcfPFREAN+0oktySB/gvEOCk/13dzYatyXkCrTBS0
OX8yhWnF1Ex+n52Ue4L61N8pbNEHzvrRa3K/92/B6EI7390049NL+rOfUe3CqZiFRo2cXmU2gFyV
9Cu45A1dgfmko2/ny8gZ9foP24cZIzmwjibLCGDfdEJmvcryhIp064l4mOBIaa9UciMK1uJRK+zH
jFd86czEz3As6STapPvZedKFcbRh0g98WCVz4afkYmd5NrHrKMVlELJ8RC6CZmgleYTmxBjIlSI7
EGb9moosMhzuRVYdbtTRBVEDzW31iup9ZE86AkmBr0WNdn9kwAoJI3u/TcbRQ3CLuF6rKkx7dR9V
QlBtxYRfqDZLq9sva+ZXcwiACbwU/4ksr5ZIotQWOVZkqQusXgNGIf24pie53WmA5wAWCCcb1NjA
RfV64WQ6W5lRmaEhEj4eoV/b2lKGuLZZiRbavaxYFk1zmO+IsLWswixOSKqjtKAglKaZ7YdUuNQy
W2h1PeJb2XeUwKPh5q19t6DVz79ndD6JvRB2xiozAyZ0TqI9osrA5QcSmWWuxfxBcw2rL0H4LI1k
8MxEfHzOv8y1UH4j+qRlmizSoU72CD1fLH2q6IGoMdx/ncuY6xSNoRmaQTaGnAAEJ1ElXeHIRTpA
g/9ihV6C5ilqEtpE8cE2aHddEphgBx+nvD/ptI+plPHZMce8tj4Jzxyh6o234mUsFW9pKsZHubr7
ANtsmgA3jleKUwdZdIJ0HYvX6Rb4Q6dxDVR3T2lfQmBKShtyH09HcJclZQvnVL7Fq7yjtsl3DYXR
EpGGMu8WNmkn0fWCPuKJJUawt/+1E+oBYcAA4j81DjDmHkRpklWdUC0Djb5uz2YYJdEgp0LvXZfs
F1fQw4hv8XHiVD9St/zAXXYbBt/c99e4YlclqkU4B8K42aoViZPMNivLod0VhTxAzyRMBxiDX096
2hueP/8lZYPV8/R/9fAOvGj+yTV5ADOkUuEw6bfZSI+7yDvTgScWgWLkexdlfsE5nQ87ERQxLmUY
ExABndMB29C2Ryx8SLWBcSo/FxOegUqvVoaM5NwbxFGdrwObHo0FU+N8ZnA7dcFueTywXZzJJ9gv
za9KqwOZcaYUZctP5E+0H06ircP0BXp2chY6PP4QkyWv2zD23DX8yNxsoY4oy5ZCy6fgFlmw5C71
1fQYWIQHUd2b5sMXmM9lKekzAV2niLpRHj9XV6rl+shH9C0R/TjKHhHPmqy7WxIW0TJ/cmFGBWjW
vbHXu6Jxdo5J6RAdamDkbVGE2jwXag6ye9t9uxet2fjkMQ7nH2SpTdu9oFExyRxRrAusiEN3p7ss
epYN6UDGU+JrOdQHRw3SYL/mwV+544TLJPUFGriwsYk3LVspHG7WAeTDOxRedc8UvdXaEb4Ckcsb
UTj7y+/Qkc1S7uaDotnv6Pr68xko0Y6EQlG6Iw8qpCsIuBCm5yuD8qkxSKKU5XuLy2Yben9BkyI4
Z2ZGwIoV/KqKQ1VJm93FaI0c8QYdKh4VPWHE1myN58/mRthv6RwIO2bZwkbUWcMtpDuHIRUlHFUt
y+TzfXDVro2+jHT7UeqmAXDzkNtHwuCTklkQQwZogshFCEWo1cmlbTBnEDcQjrTCOOVolsFHvFUV
8LjSd64L6rkqu3sArQfe6jo2RY8N36h3yM58px4A8G6C39EiA0c+aY9at0K6yU/RkdGFoGCg9AEP
Uw+zT9N4vuRefSeoMDBfSeYnV/hr3QEJPNNp6bQJ3cwA1vdgTmbnQ5s5VFobBVB4l8lx/zyqyquF
Wu5WCohh1uX2nOqXQeHpYVYLZnaDf0Gq+iKYOmyB//h+hDPNYU/TJTowOUTiYISiVg/PtbbMCj3D
xVDibubay48QaHduS4h/gm5BPVt/BXya/Xz5nms66Azz+67bRJkjnRKJkGNsE/mM8Gz05qaKeREQ
AEnoFcBDzi6vw+SdAXB5H9Wm1Hj+kHRNTwb9mXjhw+RXRHuN0BhgRMDP7g8AoaW6Czvkopbki3Dy
1ztXU7iiaHCkS1FTQJrtvk1DW6ss4/AYVXr/T9S/z8FWxhvgCESAlEzBUE/k1DXurKo9zLQWCLoQ
J46WYyWFijB6iflTfNFHuOzN4bHHF+IydwdBrJRpXsMIf2JSdu1LvspuwKpU2IeW7s5+ktBHVeoK
gT58s2SP9DuPJNeuZj9fBxOXQXpkQAe0d2nYIu0mxgDJozK+G0d7H1k5cKO8moCy2NpVVE9EDPUT
ecy3cfM9E1kakdMihMmqQtrHNPe644BpUZzCV/7fpxEQ/JK8Zn0mncOsS9jyTc6YyuOwduBWf00A
Om9INuqKwtZSejPIxl6HNNoSIBZmbtKJlJoEQdaqhG9HVVdbOjCqMmu8WcpswNX6y02bBJWp1b6z
d/BoqtSbWLpBlL1EFsE3PbaLWNinIkHjMhyiCXT7KBFEgOORpE7vpyXSDn8KLvOi5EAdRsLsj/Y+
rk/8mchLKhwozGLjqHs+zPxDqai3PVeq4FvMWL+dYcwyIGwMbzVYD1lAUS9zq5ub9ZW1aDIZHnjZ
h3H2gGLv9dr/EuvTLSlNYdvNN7EUPRydTx42s5GvG75FhqeJLRs+sPMItZCoMuKYg3sARR3UCt4H
KBbbHygk0j3qKuSWzy7GN4Xh7lYv40VJDoi4Brhy3+RI/2/1C8QtVhQMnlP+jqvRLijYP8U1Vh/e
9DTx613Ypq83hLhPjDHxVxpZxV0deeJ9yUsn7dDSqPA4OHg/5DWMEGEFaAKInKrnOloHrrM0ISdF
+M3GNaysB4aA29o07nyp8yne7sfGStpINwtY69hEjJlt9Sz0B4jBIXOLjbqD5z8aQLkIGLkM5azs
+9BI4LXMWCqyUJ9wyL3BEr7uOYNUlRc8jbP83hK1SFcTHedPHmhetAzUgm3bhzoch2WHCw1WRDaL
48pI2jMG1+NfidYcF8f4j1r59mKhulostgVRwTx5fhG6fg67SaRrIue5HQL+/YjZi8ky+8vXjPS2
y9doY5Fneo2q3fVhUo3i5xa6Se8/rcIrWCL7Selq/Valw2qOj8pImxy+H0hTLqcdAQYgL7YkWb7F
KfpX6MhZ1g4XKvOwvG5MZUtDLMtcYnxwwrCMk7/DOVrdcm/2b46oiAdu5Jd991nqD0rZBdwXMyam
eXov8bywEFErDCWNSMSnW5cQ9JakQaYP7MHWwfxBD1bU2PwPtY77tBUkYV7X3Bw4ZylBi52U1dou
qNSrfZ+gfEkr4dJGLddO6YdNHKAu6Lx35QtkjJj8W//pmcjYa5xHf1M/DF5hO7udjGllymCxb+Dg
yLPpI6AyJfA1E/yuqTXmi1aEBae0Qi3WZnmGdqzHjxwuuaFtbOO5KMfRTBiHE2XEhRgQ5ojjlXRL
KuZbeD2IvR+r12kBJYhJSTqMDTlNyI94YeSMNtnoVptFTaVZRoGgEgpmcYC8D6tpt6cFmDkiYqVP
U3eJnQaLiSz6sYiVAljPQp4990WM3VWgJqTh941P4+PTdHuEEDeu22WcUX/2hs3UREGp2Cfg3ihh
Slkzq32OVFjRteT13CNQDagkNyGZKU6AwpwSdPKJThIxLGY2OHxWy01DuvTPM7J+t0DTTwjYdVAl
sUIuElG9vs/fMnUAIRQhLglczvb2TTYL3EOc5a8mB2RZGhcsCBTwv8LdRblzo04EMaynwQriGW1n
cu6jBjFBGf3HFgH4m2JWQDxy7l4nQsjhAayQTBF6yOHWE/gQDkSl2pLtuRdZr7PhgIa3UpueZHqs
tjNc0uGfpJGCgdS94yU74PD1LFYcAY3PCMp/LLiMSJ56QFM6sH4Yz9TRHmJpcFqutfM7BKTNx786
24vHIiYf7XSc4SA8bNhmrTsnX5UNI9qivF4kbYw1WJgzCxSBw03lOb3eZpH64B+p2so8obN4R/ZC
RY8BDTUJ4l12pHNatWfYMXfRM1fm6mNww8dqP0ILdDfvJhmL2ssVgMoNpRBJW6Ro6gCXcOSOI74X
qfI7XVf9mnJi1nHDUNdSnxH54jMeyqGzAIfTlj06QfKsbMZq4N7+cCmm+t/hdKN27X7J+CIqc1PD
1iaMiL/V7YwTbvlc54fIZ2vq2ZL8vs/1Fapf5bVtP+D8ho4oTJNCabj+2DYr0beu8yg/3hAvRPDB
YoNlMXwnnuTovYu94tO9ACqNFSkbhXdQ60KngMfSWZ31KXAYIWdlDoV48meMUi4/LmxvZ5DL2jY3
90pBRJmCG7Zk5U4HkEmymn3v5uAtFXRIEZAJiYF81Z1vyZsOubKGPt8Xul8TxUqhsVb2nB+w6orX
p3qXK0i7+WTCIZdvUHFqpG7+n140zGMqy3cKcYjjYBPTMuOrFDCEaKCFL1kdf4cQJ4IC9Rx9nuBZ
Vd3vxh/z0/553KDzroWOzZ+c2Z3NVV9dokPvCnAVUf2di6SOG6SMpvScPEC1pv1W7lR+JMSMPokB
75kRLcCSsz3AAmGh8HQd8U8kjjfAXPPzNXeOe30nDbRnQLNDyeMLAD/T5B+BDdNhP798RSUXPc7s
BT+V27vkUqJuiCCJZA1zY72oJAOECb9HWv8WfezGTwW1T9dv9Gv4dwWiWo0IwhIvP9PcERwOkLWO
FsYd5kd6b1Ha3AGznWHgBHEBrRLOHNLsHu5SWxgQFf1UNLWbCEFXXgkM7IBp2iV/Hebcqoo9vJWf
h3pTKE0bCxHwNsXbkUODsk2+WY7dLAC4CDTzT+RQ1rDVG7IjdkTkTyUQuQguokoxVDaFVqXzIWUs
5651MXe1cliGzaWBpEhD6Rqix56BgZ7DZTJNKTfRKzmhFgXqscNp6MJi+Jj6udfj70Af090+z38z
yhxxxNWzuv6HJXSHi0L4TBwAEFVdM5+hhjkGcBTi+Z9SNsd1QEGnKQKz7ia0b3NclNSCE0jZJ+1U
QQGOE011jK8s/DdE+93RrNTovFS1WJkKlyG41P5YTSwW/q/2ahnhJ0c519eb/v+rPKkkh7cC4F58
h34KzPbHc37AKWjUnOvcnQFikPl2GVQk9jjH8fQbo9aCE1lSSKwteiYTbgAR/KYu5itKgpeMrLCk
eTq/u1lfXAb2SnxRuK9AuofiEawxXKksP5brAcj9UB5+Xp3iu4mh6sxMyQhsP+5ikb2gCqkXsDFQ
iQBDnESamBijmslZ4qmoGd9O6xvtNKd9ojo4eLhbKXfG9jNQexCeG8m08w832KJLay9CgI0LJse6
RnnBqs74adAdKlDb0Q9Ifnyw4oITsJCR8hd8SORrL1zyEqZVgJRTxzBvlvtDXPkvyUvAEXI1HUer
OeRKF9VqRN9CYZXTDH5tHKkhFENB287OFSTEJ/t2fnRkbVyVVSZ+iO/gbp1UqjZ+lZKjdFQs88UE
IAuRU6rdnmD4DLsRWEdK2D2NcGWRDVgKOmU/NCnR5pCelTo63xaKW5ChOlcV/crrU7WiaGJmyLHC
Tjaircikkdi8GvayesPuC+t/E3bgB8k5wYdDftEw35FQTbzMiT/WqWL0kbN2JD1xO8DKX6dr9kPj
1bQSNcb/zXXQLkbHuicbVWg4iTGP7ANwkCnqwJ894W8L+yb+y9fXfCBQeBVOsTqa/dpzXWaxVI+g
Ye+PdpZVwZo+UDi/EqGDGIvOkwRmaUtGfrdiQ+RR9Mx1haYZd6rKzzvqkP+SAonmqEoJO2Uonv8p
TfIRup18n7H6I0d/Bd81927EChZ0Mdt7KrDP9L9jQUef6tR6/eJ2k+XtjmCihPl32oqHP//URK+c
VaECU/n5Rf4/KofbscWpMFQqNF/mF6l7sVcFyOJkR+KyYY7HME7u7qR2i1MW4utfMPuhpgMDkJH6
HOk6aCngoPFtve+2suBMxhBZlj1IJ6Z7za+0J4FU0JBufi2bDbGPPp+OvDvmb8RaC79ySFv0fLic
rIadjMJkGbPghzECNJaivTQ7FlhlTK5B2qeBfD5624PYLPapd4KhpcS/gZQXLW/fxRpLnft+in56
xDwKF6mNFcHXYuv/+fokqArevZpI1M9NrkNmb1fbyr2ZUfUe3nIu9cwTYaJczn8PgJQvrNQbUyvA
qlsQekIi2Yq9bMT73Ejt+LNgmMPMRtau5NuqIwq+kmA2/2fgMLptR5ZifLrPwWLetSZiI6MZr7Z/
jIkt0h7zk0ngXfAYnn85fPxICfUpFPWrsNGSdnorJNSkuXFSqCP3/tZW/0kECmPnbEggKF1j99LO
ibKQr+EZNxF5qynh1inNgZBUgp5Szs7Gwz7wP+lD+tMKkPzsBXIZoIu1Y29GMmsltX8AxuXxHjbR
rvy2+4mFvPXi0AH+lg95GDaodnqLQ5X9lts//HtrmnyHFSA4EOQuSHwM+NZu/hMBYh1KKKa9HdxU
MOZ/xgSk2uiShBdvjKcjIoEIpdOfDadKaqbC7LrrhC077i12bOUEAQ12EXqG77QN4X9v7bGiE+vM
4FqE+CwvSOP4BEMyU/7Lpwb0M2gFA1ADPIGCPpjuFzX7EZ9cTTxQHh681t8VLDUE1v9PzOjAMwo5
CN/fhSTyy+0OK6dRt4z8GwbTEzWjtZ5istwCmjZPXdyUoxDQ+pj/nnaQ34KrewlIihWWYjCcHXL/
fldB4s8nN1CXq8MrvVGvt72N5vEv/7fiatuhgXEYUh0hxMdj6Ih5nZAJXa0nyj+d5PCcKIy656ko
IG37/owS0lIXrK6BzOrNBZ4T+Kp3pgcM+aWf/kyhIwnzWZhAHjVv4LJqbJWUPXP4X7uDOR8rJT9Q
ANSrdi0JPO19Gsqj4C8qVaki4UTteeVaHMgdH2FwshU43ilZ/0QS9MNSYEOe3mtKS+rxJm5bnFQ2
CoxQmYah/mY2+Xe7W+hQFIMFK1Vs66vfUjXIHvfw6tfKoJF8tEUA5j41VJ2nubeydQgAqCp46xVE
lxDCuFcaX0OxdK10ryJetYdXvLJRbCLN/u2yZ6qEAJnK1/fktQ8xElbN+GA9AzixjFqHrTJjGQ3k
wIkvOoZ5bzVCFCW/WtdWjiKIGOr1Etoy1j3k7+Xp1LuZNY9fvgKVRxS7NIg3j8bZ7tlfv0dBdEW0
ZadvuXzudWm3jsByLsJbPjFjarf05XrKvdYKQeme8s0LkE9Axfkh0E9mlVjlRRUCdEG3aoaeSQTe
M7svbX7ho4aoF6SQ23Qo1MNohblw/piVfPifWL4p0QVyue4hwdMJYXpGRTTFaJv6wkx1DV9XgOtK
YQiisjLt7DbAUJI+bpWC0BxKuT93brL5Fby93X/u7sn5DQW2q2uBq1qoL7iQWCz9osf4GcsYMYX0
2DVtNKuo+F6MK0psXCEGB+vBRrHjoKRt4vu6Yunhx4yl9sbcCXuL405buVgfg290dOwkr8S3XwF/
hemnLyL4DsG2K1wvNV1x6GLikOpv1pSzuyY1R6UmNcIvYmT6HX2rah9y70VT0IGriI6WgjIsxtoA
o0eVBrf+sI1ac61VPVFsh7ccQlPP0v7NrrLhJfxfKls5BelpQYvCyXwO54hJHCDW3HDw8LA2MFAp
TXNCSheTxT4xnCUQBT1wklmrtz6VOLkj//6DOOz/R3Hu8lG7psKTn1ltxEX+2sz050M/3A164yvE
mjWGF7eehiWAamYsqSv5IYzlrWLtCHGXFNvP7/97AZGvf1jucbs5ZGQ+pDI/DfCFotvtSxPlAok/
t/saC/TsmpEBGnUOBvy4dcZmf9zhxZqvsvKdFNCISBbd16iQfzDfYnt1Jru7/jOed8t/+hnAsOjd
nUQNJC2avIIm6ZWz4pDODMS3kh5lI20yPqhSExQjM2NgEcQ981uy1zSJfvYNH+XCQZjYeEYWbpZM
C8FPYAdz6h0owbhYqeRSXotMyNiC+cZMMdzr4xZ7gL0WU2MontKoKhMzAN7RwHEBlTsJRbDwxdkX
PhoUiwmZlIbT/BtDtSHxw113KEl5WQwHcDmzujFSwPufL55an2MfZ/9D6VExyfpYDLU1KAet7SHy
5SIsezZUJsTxTj5yCJOhx4WhWeUYPlR31vEs9ZCDnxKVEzqMgGV52TiQXzPf7JEqZrhDThCxkovm
VShu5aZGFM401tYDyw+HxTXMR16Gd2eJh16ZORMXEvrorCYsvTHSjvB5vW2HMGbduO096sm8rVnx
MRYmeR/c/PsrxZCQARQMiYvh3Jdr+u0saZWyhM4IQCNl6Ro5tpvQwQ3par1xvE1EunpGMpMc+itN
aSH+5W3XgakNAwFUDEiku2T7iFHCThFKWpCDpz/6BCdBugK+1BZo1tTbp76fTZmOXqHRjpmiSoKY
V5l5DDzB12M0kLQFngDehnt7bS0sx80HBvoAxKhStX2Y5aJ5r6zu3lLKCyNVD/oFnDqjf0oq5xDT
ZML+9O+OrBJwgf+LwDXjaJWtn5MTvvrC1dVx7f+oeBY7zMfONowqRWRZ2genhDLGQ0s55RiwatSd
HwGtGuftH2nE4oKR27EZZVGxo5c5xqSjAmNG030LEcl0gZJmvEAFY1KYiAVFzgV/L941+782NwfW
Ofrk0VCf4OIxOGPgpQdMuvpNRaTwUS98KrTZLLI66xO9qgrwKoJzddwRB/LO3BFaoiqClVNuA2AO
P02IEBK7JgAhyMZraIbtIP1zv8/rkjrlQ3Jo/LfCQ0MfdAs4W6BlW3fGRn+gp4o+XLDHPEz2azUP
aCYUPw4NbO8HWhM7S5UfYguDHjkINZ1icJ1PS5Aw0+qlVXZ2Pl16/2yrFbX7gRT9yo48K2rMgo+c
LCrIMOOjRj8dOno/VnkrVa/mb0tfNezysNxD2u3ksA0mKi2Qm4Q1xAtzehGr9TI8TLvWZOcRk4EO
lacZsCJ3sg25+Z4oJm00UCSRwY5NnHuMlaQdF1ecHNl9IL4rqIyCs9A3PDMTvcvIKw5VEFyX+ajL
GtUA0QaXQSZp55Nstwsi7FemUx3dCgOoDYXmHZkhc85d6RXW+O4tvPN9Rum3q56c1D7aZd77BjVf
6753o2DnQ3Z14abUWe5iolmxlIy27vDDlDTZm/uTg4fCOwxzcz8Alnitrg26RkoqKlPpLd7qGMSS
8PiwKLy2bGPecLxt6pwWd2SgW198aktoOjTf74QkJN9C+OhTOCKx1mgjPKWrEOVj0aksGfbVqjNH
G+5iqqmXgIshaA8TgVfvyzQC1g82ocxiUr0pgFIsY8rQeaobIh9PY/JdbhAIk4++NiYnk1tvIpc/
AWOCy7qJOIvmXNp0T44YXZpUo5adsEcm6KCcNwpVxzQNPHau63nXnDvGUskpBK5BipvhQWBMwjed
WqWHNbmtWfcw78EpxZ4EkmDgfoX/qlqu0mD88zOZgorb/YVJNSctrLLNOMXxMMxbYFfIITYh0/mF
7WEdYuqB0uyTHYvovrRHXfThNf3cOi76qwygjH4TAB2WnS9BenaiPYSviu9659CPPdGJSGFUeDlk
kPjy3QxwRQungg4ULPYm7Sl60PBUMLgPEHZvnQfK1aEFXY3pETsqjuGKewOVs/t6WHSKjab4ezq/
3lGZPiy517CwZ8Exr+78T346Hi0KjqWcly5WOvWlSEwwmLNk1bSs5r/DAzgxKOopyGu4gZ3F5Zld
30+WCSv7sp3nqRHfFhfZg1em13CcS9YWXvgS6iZJsFQ0nKlJGgaRgrwkwO6f0S6x0tB7HpKYv+T3
sK71b/aiy+exMu8/9iZjYmKYZXvoRLEocyJ3EUYmmBpkqUA0SeY9UKzpet+dGc42sxqlbkdMXlIA
JdVSSilHK7H8MQn5cES3JOTTbHdvUitykA5LWZ9mc2Ltn4FBh51EuCJ4oeXq85fZfn4j92b1NXxz
4UW8PDAB95Lq+t0I960SOMk484bFxhVOb4nF1im7I3ZPcTRU6/y/beHjXppIXPClkfWFZUkMMirx
ffpUy2UY6Q4wMaawFY1ocKpdVp+8PmNL91dlvlwA52Do/1wwVp62iJLbrJuHCZVzS6Zk3Lc4wNKN
gayrsqiUgD1h1GK+E3bJzA991WmTs7DnU7AajvA64tIZSFJ6rGTU5S+w8paxvrqCzNbb3/IRwZIt
gxsZttsBiXuLQStS6ZqwZlXmsJ+YxzS/lXxSf5LbJzZpsdxBU+32ORh5d5sRKhtFa44ASK0fWoeM
zg8toHJpdTYbHQtaxF5rRSu0f5wctIxu+gz+SGQluEIpd8nFt9/d1FF61/8RlabjAZ3KkJy1Y5cO
l8BeNTpHM90qyuiYNB11Kv2rB32s9uB9FlY02RtdIkIXJQJBl/zY+jN7HIIS/4wdmjTNoUKgO0Fx
9vQ8FZgy0fS4sUyFvhHrHjIAjpRNjQXjo+gLTtYHoWk87EdvV8VFoC8hGt+cCOFqRroW0hUl4wwE
EWzlslU1hJWSWLIRTeGu5Et38YWXZn+JWEfN9IPYjTjzWVIN99IPdVKG3UJ5p9XoNyqeBp0gwwDg
WpE9hKeGWWKvGEbaP8NisfWZyzleaWYF4ncbE85WY1/reg8C7xN9MticKaBCY2zH+NMvLX5Ic7xE
2Bni24yAwnGrOl79y7vksZs85cCT+Z7qP/jaVJuWAasuwFKPNO7biFpW0cJbbMIr6r7NGmcQswXD
2ruRo7smNxIh6spr/34O3dZLV8RO6fvJhWzViGO/ldu4TcoCPSnZk8bVNrlpCXMfwDGa/0P1yeaE
Qatap17D7obJrt1LqnpbGHXJ+feOm+Eu2gKiQEwaLTYpU1HgQI6Wd99YbA00vaMmPTzIAzuUr8MF
ezlOUcxHKnj6M97N1i8Bzg9LGj4FIYknHfomhIOPwmWiV9Bl1QsGh9eab5+i/T/oHjHVPXDd2ECr
EPJjD01byFGMrb0WlLCdX7PP09dj0pfMMrqBqOhz8scPTHTLEvuxe3HcfJze0NoqAEmwAbd4uL/z
NYvmMBHclwZt1elZf9JJ2nyweL+LZLbHy/dKCJDs6oRV0IVSYDO7O+z7XwIfuixoTQhT8jSzAIuB
v1RDeHxHdSQx+YZH+33OeEp1iggCqyIX0ZRU5FtmACpgfNNjU0azPtPez7XqEWaQvKR711EF+en3
/Ua1Gfiksnw/BfmvN5dVwwpcR7/fG3DEB17F3miSlTo0AwUYBy95q84Wz688u9g/x1smt5uRnia2
p0FtdyeUgXxAWVb3jYmD4CKgUrqXZRFkFI/rQPySsXIX7VzeCfXpLykVUJ6Dksq6VfJZrjaYHie6
HM/hFNW7P+gotD/wyZINr2z3HHvp20/9RuGCW+A+83lfMMfmtq+aB4vmTHePBbvLugxfxeSN3HSp
Julxq2g9pPlEMhf1maU8MHe4QmsrkgYBpi9Er5kXW6evSKpTlfNDqfTBB8qOVtS2DhMki2ZlVsgm
7L530Ej4tFLnnQU1XsTmoBgcbIxaGba3VoHq5haDOZfhD6GyHTkB05Wl+WALYi95IstmOSgNzEm6
m2S31TQZwOprTrJFXYPAt8AC/PVUrfsG2oIL3M8RbE1VZu8MWxMqCr9lrYR+/ACy+XtoGsA/hi3q
NnT0Bpx3XOg45vbHazsASA4oxuCxwjukkJbMudQB8RWtArKnKLgC0mt1L0oB+PwyLOazLbyZQVvN
p5hFyZ+W3BZ40P8rUw9Ad4QNqQIWCXwpiRQjv4Tvl/K9FC/d5/JWqhB7poZdrlFV4cwBsjpoyUJk
VommZPPQuQ7ehTy3iUzprMoG3rgYORCyfy1Zrq6dYjSk5BmcpnExPTaokGA+d0R3Wh9wCak3Frif
/lNfTql+slWTH4+u8nw5swfnPYXG8ukJ3FkK3tc4Auj8OOyFJhhz/LxTQTn81aXpf8AYKGhz8zOA
VyjJCqFnMRSKbskwx4w1dUWEjsQYRFDS9rEc5kx1YP275GJWE+bWminGQcGHpCFuHB7qm4OW/tay
DZTV7kRtEw8rAXDx8NuxEHfE0/Q4qNiKH8kiyRa3NM4555W+6FNpmVoHc92gwzit1wnB9Qdzgj9b
e5SzVu4Gj0pq/ycvyfPEZd1lEELcJOowWpabqRgZqJwnKhmkPGw2q8/zUlunG67WOFZz1aQcPhe4
+ABrpzhxID9L40+/mApC1Dqs9QONTt3pGqhTF8wV9WtJeqUL1HsKo57qUIc7cq3iw1C06NcQNANJ
m3zDEvA9HWjideOwDAVNkZyPLunAToEY7S+sXoQ3WOSEyr7UzhyapJTMxudOGTS2/Udn5IYkvXpV
PY+83TLxohUj0toc3VREgDoRlxWbIajYcx30nhm6/VSDbzK8vRep0AES+Ea1ok739rtl1uTxMzj1
uXMeUj4YrzzxI89rnN1I1+2bJVZpyBHtkx5rEP93eAqoZAbWO8mrWRDOksSJ6DEJMj8GTeoyOC0r
sgMpqhTyn12G1BpCVdTYWpFHxm/xbFUadfTHRh4LhYNZCEMtkgk3rj8W21DWRhiQk2iSrG4vzj+4
d9TldEHWiVYiAQW5hg0ka7RquFb8thGupDzG7dZ/Ao4pGhd+2dahJhjHvyCmjS+WBrYKx4abaAj7
/ko88h2HMEKBpj/cm4TOGyNvF+ZM97+JHXJx0rg9KGidUF51ukE4EowU1+AsUBiypB+JvkR/mJCI
mFXh4rOFxARB1tfo0kVGzu/m5tFabCqqfJhuTWm/sVXYTKEAHVQoG9A/bOHhu/v84e182x8SxoNO
LlaiR4ElaZsKyC3m+oAbsrTmMmZmwX2xJPThsVEeo+WhO26wSf6S7TfgnEqBKw3qJzpPxaaFbEHD
MH90hbodOO582vO/xQRoDa28FSv2td3n/DUaxxlmdH+hxPMKketoLAxBC4MHqSGhqERX6jbOok5i
Ixz2+jfme9OWO65quA+SXjFGhIQhXOASrA/dz6YV/Hr6vH8ElMRIf1xLj0jpmWzRj73xI2w+PXck
FhnwY+vPNwEtEDvyGPk0mn2pzH2ICgnknGHqmiFynxezKBjECSOGCgYnyqeWhe+QtzSsgyfdNOrJ
2wEzDNPj6GhY1y0eQbY0JV9ySgZHjjZKAG72eiPQUo54tl1LgHGiA7CWxZRFaTudal+psFBMJNlm
QuFdh+pni8eaZ76xhxzCdlPv9AFgOOXr89M3BkoGZodocOqpgXTpFHvzGBo+qIM8KDyk/8Am+Eya
kzF6U7yMFcLk80eDeqrrcvhUGQGopTne233nzSj9kT19VhvZa9mi17C0Xpi2cseFmp8PHSXHIkKa
CNeY0wnLbNrk/f96SHrYcemKEhVO7mecLGBmx0bezJHBoC91KweEmV5+XGdBpOnkWPE+OyHOQ6eM
vEQzw79jx9OH/U5NDRH0t/E7wFc0iAh+CCTnQKss2Ot/EOpi6JXtcd90fY5QEb2WgJi57u2lNW8g
tToxsAv92mx1Rj7mqpsh6uf7474oP6+rSI30r10gMrBrsAwPcbRX4NqMHGHCwKi71yRsMY0RfCXJ
9ImIjOVe+U4GfRjrysaF65WlcDAoKTirYOncwRkYdi1FnBDtL/3OYy39+QPjw47j2u0MFd23G65i
W42as5KTFRLRIgbhtUoJH23whsKdMAGxoF4En9GIiWZc2hyDSEfHA+YRdtZLxEbdX7HMAZPhaHKj
hIV2Zikt61WhIDXBclZrSNuvU0a7ujYekiey6MHsd7ntOblTvycHG60NC+29izpFuq523kBKx885
0ir3OboM6rbZGvVtbt8c2E/kuL/lmYY0SOI6136M2+sM8AmckAAKuH9Pcd1dq2LYMnwcvV9OVd6S
V5yojhGV2cjSMmuaSMZtpwHaC0Dp1iNyu6madfgK/B9vi0RXM1po1RWoC2eQUnONlC9VA0SoEiwn
IUfVTcZctqxLZpLFceVrwyWHWwCbtnn79nZfRLoZvUzLMSI112mE2bcWa5948SE8aWHqI1nOXGVy
oCZqGlkas4iKWuhlSag/bS6ijhuU9HYVLYPbArMcV3wnm+WD3zYsj2cEXvWcrqkKko6iQGKPeyUE
HHz1kmY6D99Oqx3+NNs5TW65w+Ov8c2nTqXResXrqVcFP/kS+ydYboKMcTN+kfRh5xOFBxh2cvGE
PZSNq0ofF7tQlMSZxa8eI7NbCTP6m0KmkkOZcMA98OkNE0DLOB5g20iLgwkSb1IgRBZLTKmZoC2l
Qe2wzBBNp5LwXR4RiQTnHVuAGH+/bnvCL550sYSC9ujPSI/GPdGGlAu18OhBRxNS07xoqUAbOcsF
KXwYTrCzVIq4SvV7FyPwP4tvkjILiV4wLavTTrNrOKPb1Wjr7Id3YrjYNbwddzhVD3UXzhy7OX5K
5oMULmUmfRderBdnpa44eZG1lv6X/9RcRrU/IC6WTmvotU/jeJ+sviQ0hWPpnZvT3VO+DPE07J5H
yxbeyoRzcsOgxMah3zkinNpfpYZDbxI+V4uuybCe64kL1xV04Zdi6rIkAaZsTKualC/6pmsWHwma
M7sF9PYXfmIOJd6xxSMHRUik3ZUAKyGCXI+NLSC1qby/eW2I2a53pJzORdQ+1l5IuJQ3J07qcV9S
TihT8l6WqL1ACKuS19c2zWJu65eeaLNMRrxvTyIkoEHhdEmmPajfnVmLYqItcRwYkFdE9MIKbIot
pUNKNiCqy5Lg3b18xD/fmAwrrDqryhRggF0+iaZMs498Bo8ldFKAjGsa1GvwfN3H0m3bV2QfAsow
GefsFNT+AlxMO98QMHn8nuqk9RtyoFyb8CAF39liaKPKam4shCjWtmb2Z5g8XVueo/EDfQXi5DIZ
sr6BOI4TbaboKi6ZYPXKQ9QuaLvFEtStXOlvPfFD/C67dKe89qB6NXo8BNdV+So6p+TZtks0xe+k
41ZqLvdldW7tqRRJTnIPVpAfo6nbXIu0Vk2voda+3Kf1ZXSHhb0RPAHrn6OPvtYCmV8gITtuvlAj
gZ39k4+HKtAABSj3MQfjjOPJLJghhhVoyL1yMt4apT/aLmNiYjVas3wlkx2FvHWp3yxt3Kq0vVn8
LGwtSO/xUsZNI2y6G5YO0LeZZjMgFZcU1s77iNJAjB7CVei3kw7R9CLN2bJEXKQvrzySUa1BclQG
KwST0XelZeKkJHDtBcuuC8bqdeNAnxhDG8qS1ykien7/KFyNiccrN/wbBc9zcg8gLxbzyhoX64mc
2YiNKKdIlT25GR52N0R+g7hDwP0H9B6fxR8nd6mNIh8sdvIX+KUh8boRzdHnN84LoTJpmeHGpm1K
TvCQAoFYJBxUDU3VgjoY0Zu6SaHEChDnB0frG1lGu5CXaxO+sW6HVZbsAmCPgkI0ENrpNjklcWg8
u0IYKucp+dT7EWNW/FP+dcPJJTBG3JINe8phGYuPC/50vq9hIFWaD6btG03VtfgjcEdoYeBtUBr2
Y32Ai2u6HOm6VBfe/Jigt8f6J9T4XpXP0PXdgf/WVGo3XTCguIsSdH3Fv/MkGTLGwmneVHZ2NF7t
YChEIPbHeIkviX/MwyJa5GCB5F1mVqzTe0h+Lw7r1T6AHnVHGygaxUucTQvSnbhWGVt51eYqx23S
GL/ryMtWFUArApx0gECXVQss50vb0nzxBAGjFT4h5gmIVRfXmGHThVvHC4VCSq8xXWJhvAyRIPMx
5J7RuQOAc1nQuy/Ky0E6Obp4ccTgXR1sNbmqTD2BDkDBWYBSGtb0Xhto6mEENqZYBWj5W4zopltw
nIHy15YrA/LMihzVgCIc5Ov4WjMFHSM5DT5nm40mp+gLuMbrovv6adelexff1TrY5g8DBDKVLE6d
0ycT5MFIs0zNcqlkW76z9/ivwwnbSAQG1Y98w+REZgxU0cExyGMgmUjuG9CbZ/7kxdswYpScUk0d
KqgsZavwZE87GuPTWI5nfgdK8ribainPo22qA6QFPt2KO5kyNK8AosMDgE96vcwYTI6ugs8C6XDY
lg2CGLltYz16IHGbS5Ah454HJBYeViC5KQ5dtNyrW3zZDmAKVX4BF2wPQ7mRHjzi1teIonzXoE63
qOk9QU9pbOq3QGHJ7RG8fMjs8mSyENXiTlyQLiNSVNvKgSo7vU9Dz/Efx+lve2d97EKTCDLwIGXC
ZqmHeDj9GxAWeX3BH+x4Oq6b8LmRaI24j3tOC7GEa3kXbJKp2poGedFxs0VOJ+XGwZmf5KLao+8g
wyP4QS7m9oUYNxUd3M7Y8Ox6sMpqWFax5DxuuGB0fwOMUoGpTb/FDKKUqquftz6GeOfsgMIfKpaR
vJsmfYEf/6blg4eYiM2+H0rVDBbSYaMHjmQYOQJZyM0h0RIFOgc2VJeJlM0rk4l32ju/Gw/BmF7G
Lv3PnmDI+HdFplPnRGSWN9aHGr6yxe/tPh9ZaHPTahPSJ3k9sRiwEAnM6X0TgDZ/Qzdf7be9Prm5
73c3fE/FafYYEOllfl79gcdo0x8TRnDIiwJMolDmPe2w2PfPXVVcmi0dEbs5rUc30O4toqdaar4H
k1TwiQHgxzCdV9AONfwaOKsyfWxIJ0aBI+a566Dm1cM8/dbeVMG+bjYt6pLou+P0IbXNZt+Ds4JG
654yhdwUFI/KQXQhwLrcVpLjSTM6D/MsUxS5ei3EsyApjgnPBGGnAUGRh9870Rmy4LgManFanz8G
nyY+lzAWhNfw0BpcnKpCVenCdkIA08aL+8iEr6w3k5U1Lnu6uriS4mpdLj/G9RcBgarZDIeaInCZ
98rSJ9ZfynztOG6AYATWwDnSJC/XaQsles97sVO6cIldqwVGKHqjf119DUYObeKG7Rrn7rjFo2g2
ZyqvboDZBAP37K5LndpQgPjZIID63tu0Bp2klN5L3w79Hwh0q69xaXwKdZ2cQQlRqiB5bK3ySqN4
zUV3GSGBUazsUtx5izDA67nvX8C967J9dcfObr4udtA7WJp4raqT8T1dGNskxwPDAlp8KTALuz2r
KhMqK1tOW3/WxwDgb8eXOOw8rHgp4iedzsuYENVQxtS9864fPEFMoVZkID1yyuKS2dxXe0C7vuRH
b9+UZtWbmUQyea9VjecKKTPy9ucZoW66KAAEMjSCImmTqCu3zh2W8lIYjQ/dEOP70DHbTLKoWeNX
jWQRHsnCjml6+vkfb/JpYx3rdQOiB5nvrN/+FkuiIk9qIMc+inSCJ1HrBj4X8eLlxU2OgYSjtx/3
yGb7dFyJ9HGFU5yp0Eh34ih2r+S60vn1tljIWgE9xfJAykFd9mq+KpkQZgHA3tKgXfDrfkXt0SAI
nqoq/TgMNek3CHRDFcFnFSuwbN1lSOFDla1ZCFibgpP8vsFcaf2n3KTztn4O+h/Hmqd63W3qu6P7
K45HoghvMwSf5iSRGGqpOpVNvju/OAvobQwd/QiyfPxoKl58J2GSFrwh8zsdWaQO4c0lTzpvZpwt
I1SN1y15+bmDaTS9z6iA/GPc/UWd6gczlUha6xH+rHEWZb4XBfRuHpXaClXTZnmJdttW7u9+KOe+
PumfoYx5gqM/rIblLtuUQ8LrKwQiq5IIS/thfh1OaXTQ5cw+cf/zsqS0V6TASUoroq7W0wBBMOb8
I108bOJFQhat45ceG0dYa8/MmmiGCy4WX+7B3sww77zqxbW/kMMEYn2GNsZNv/hnRGfRv8tol5HJ
Eir5rfTr2A1EsaWillJ3MIziE3oet1hcVDJ4OldZ9fvqBWzsTp6TLJxhEHBMWVNGvYXuNInm8laq
C6a4OQJxdefW3T3tWIa1Z6yqBIJTsRG8TSGnEPaiinc5EKJ9WT5fTJf1Fn+ExO3rsC0N7DlXSKj1
04uI6tHKYZld/IFpGdAn7m3tfxrHqM6YqhlCLFZORXZZEN1ebwIHyc0Tzw0bIvWBr01B+jE0u32q
WQzFsHthm19mNkJ5JrzdQK2gbfAh3OYfUO5QRxdscLq+0xxRdH4gsO4iYAudoXQEltdx2jnxzrWu
nvRCV4e1SDEz/fJGSe3X8j7/gTDWHpWi1SO5YmiQs5E/uDXfOL+U2grZ7Isoivy03uUo3lPhdWjq
xP59dl8IFuscn6SpNt0ty7XNQh+rqnRGFagsY9qHEpZn9RJuOPPKtL3WhNiJ/wPzUIzC4l2nl0pe
eJT6RA3tmVapNcJ+Db/ppnuC7mRuzfy/MiboBH3yOj87JP7fsy/ZhAIi5DcVXk+p8Po/5Cp7kVMm
P1oeb/XbFv6xwshrM1UXh93Z2a/qNZVd55LrUp21u2zyLZwo84PYFKIOsNT6DNjb5UGMe4EvhZBp
0G+RjzxSRfYn1IPo3ZN8EgVrqeuoesuJZPUWolH36SxzjyR/3QtGj9zG/LLTux+rg1K+KBY5TyN2
gr8YtpnehkgYvc1CpLOtxAd0S5+BhiK+8IkYlbntUlBqPFD93dskumdV3Xt1mlv0vwB+imDFUwHu
0MZXYyboQg3X1L12UAKWd4W10pOAcq06pqraqQ160+txJuAq763vgayYcfRx4sGQBgNKc9mbqQvl
uYokF7S5Oc84hMoFatDHfa4zFK0PPtAOGQ0Cph+b+KZf69etFFXHGKtOxdqIcrfQDV5bOXzb65jT
ml2F3LEZXFgKw6RlGZkem4F7ntQQt5aI7mwhSuj9NKaJQ703gCD7CKMKvxi/5aCUQB4MKAtzg29D
hQwSu/txZ/iqyiTjO6jaMXrWcpkIcUY/gzenevbfnsmkU0k6yUytoRTPls9HB32YTrfTIJl2Johh
OjpI4n1RhUlfvHR7wZrSXLW+4jdn+1gQYyh2Tvu7tAFP9D8l8ya2We1DPictMyTr01YwT5RhMK87
HN/+5Ewy3McPtlfzx+lG3TNKRy6klX5DpWfjyjS9IWiHueAxjrwvPwtqstQx6QOyNgU78fAU+3Op
tk+WtjTCmz61ZyAiHn+AQF3no4S2VrPGgQGKUXT+FuA1j3LMfWUvYfQYb5q0HhTSbhgxpTvtD9xi
VM6oKBXV3euz5ZKC1pAaYJxf9WL0fUNeAUBbMSzWmUApH6LrNQmHR3frgq4fcT77D3rR2m08BSyi
Jzu2QttDdScXtAJ6t2yjauNUI/RaCBrL/mf0WQqzrFkafvUCVM/BQ16c6NAzTIks1lhn1WvNvIvI
yDwqkfD+5fwwriIaulQ8k1hQ/58R2PnjKqtEXp5DIfP0IFgTuHhzNaFRySY+qxg/yYd5O5QkgP+0
8/htXbCQLTHD1E4Lq5pLuZwAceoXYD5rxe9807SnogIjn7//RnoOkgLn+dSP8AxRj5WD9aNEe/yQ
lmv1DhcesUEdIW1Ve+vKCl7wTz+mZSmujgq6EW5UkZrNsize9TZUDJIsX+G/LQzZOuC0RzjW7z+x
tg3tgZ2kAY22bUCoPwiFmYrk1Lb7Li+yU4MquMb38iMp+IbQ+kTbC+RTiY1rW0Fu0Ki+OVGp9H7V
wSdK/7Q7VYkTlCcqwjxOvqnDbg4RPxEUIE44glW3NFsPu58C2W6y6NdcEt4PGyZHUB2U3D1uwznu
ZLLuZMBCwq4mNIxBVJEF1xE3xFQMhUmuHA0bvqMnImXyUezQpsIw4G5O4A9iPeR5cDGiF/W3oIOq
SYZLjQDLzTT+54NdYH+nWsrV4qL9OcBjnKKRqjsI34f12GU2IYymZoR1P4zrtB6ARNiSnS1gk8Fe
WFQHvmVWwGwgswDwCb5luTDPKKtUV1o84wHaT3Co9TT0xNa8HCSyRzr5u62+0ld8tZYfoVaef8/Y
uKqW/P8jiy3BFqR8hHnZNBIBmIVWeeuNM8/1kH7abfUyv3zujysCerw3fd/6V9YUSB+6pb3oNMli
uCVYTxsH50X4fb8w4TLv90KfPy5mh7ijzF+Pl3VwSpCd5F/x7m/MXAVK1aQkYnoYDp3Nqhbr9rsI
nhMxeLAK2b4Pmu9C0FFAUcldgFdy322wwl/LedrG9vLwZt1WrNf5lRdIrmx9jVkb4grIxlNIpqhK
+CtX9ppeThw4fnfhnoHTcNeQ8S2BGO7hGT88JFbzBqRgWGl+aiXlciW5yqtncsTx9lE5S723LSgf
n6NMIfmzValNalJenGwEkc4BTCskQABifEuRMYE/dQN82nkqNJFaaLwAHebOLKYE6cV9pTFhmXxf
TgswfmeD33OifC3+vy6gPiZ6BMVW/c31+hnK1InTDV1iW/176BqNj6SaAk6128NQkH4R3Iai7N8E
uQ6ZV4ZRhqdFigoWYoWYdJ2BquWwdyxbmeeS8x4ejMfg0Zob0vpvlOwNjnm3D1KYWKB5FH/9FVrX
l7LiCsWY3TueEETHlArNW31kNAn0RHYnWqD4ZT/H6ygcO6jNK965ytck0oX1DnWRYMCfjgvmhxqr
WvH0Sj0FRGJV5floEXqo5nlobLQV4QOovJJtiOXiqINotD85qnSNzpIWc1PR8Q2hUCJZJhKLX3Zr
QRaOFdQW+ecicCGydBXBH2bRUvbjoxVCqxyl5NmuMYho3Wuj1hmnvZ+dyLw9kFxU2v2y1K5ZQ3d1
jSTJfUjt3PmSM4nWVXxvQEFw/KqYu3RGJdi8eIWzO0F0AYw5ULdo96Dg5ZszN2fdVOeaPpNO0RCX
jdacQX3b3g5f7aCfIiPAu1HhfjYKL5F3TMOfZC3Lp0nOCqLzU1hU1/d7Mf5RSrAD369+b2QEHdbb
P63ennFivkpkmRn9JlQ8pzUkEjqa9wLSCQeAA4oHsaLPITQzWsQ1SaZYPoMp4EVbF1f9nzcSRX6d
pVbgb3pmeDQElo6zgOH7xkzntcibmbXBBOR7i1pTVZrCPaqiY9qziHszr4FPiH6qWHcKyTd2dSrm
N2jestFnodTBsLCcIKl4WO1HeT1pODoHUlIxBfgw29FnrYtqka2uwl8lFtIQoyBEHOxpnrC7IhYs
ne6szQZM81ysrrH5jcDJzKyMKowuH2ZKVwIlPxdu9ElRcwenJ8D3m2EWNN0w8+hNJJQU4TKpcgF2
YOp9sXqdzMsJukbUoFR4xzD+kHcr2WlofwN8XO/R6loRv/W1QrAWDYAHSa3hFsJaryuve8QrFBWs
YSPrd5cCZLjHLhsQAx90/dhJ7MJIfawKxU0yiMOTsDIwihk/X7xWsOjs5xdws/R8kexaB2FiHiYg
W6QRRHpDJlmEYhW//7gmhn5hjY8IpERUf8RuYtPOEIrROb1orVRvUN1FnTPc8GkLhJw6tlmU3iUd
x7ztam4qHdAdxZyGrFCnRRSR5nNdq9VDyaYnwMJ0+4MznMmptUdf9fSqpXEgk2C2jYTSlRsSWhLa
T+O4nJ7qn1PL4UdNhL2YOkcWQfPwFnBwD8kkMwr03B47/k0qVkpPW8LYiUGQCGUmdax/llkWfsq8
a14bKyTfm30SHOBuK9mNAXiR2UU/ACcjbNcT8gTJd4XBywYWJx5daRcmzrZRMdhohUX+fYKCae8D
cs7b1iU0YTTAjyUMXvnIzcBGedjKKYganXgFQRySdnhXaWx62my+KGGbZUrttxzkUoF0zsu1uRJ7
6IlHDwUUczeoFzm9NXx8L7e4SZwNsuGNQWFyrAoJLauQC/iGkplr3sVCQ9oge4zj1ms5yomNB+kn
dWsG48Vq9myEJhuo3NoKTtAOb4L2E+aV9D2LDn/UXtyeUYsuaDv5vK9b8HYDvjrH82Od74X+SJXd
jQA7qCxH2kJ3qSShvn36EipYyGdBw39V+K3/OiltaGuWyaF+c4Fk5VAq7yvUYBoVgUjqnNOWuoHE
R8FCWneu/pNDMiAw7H9dLcQe+/MpHD+HzX8hHYlvmnD8Q5HjNK8SAnAAVqdYLSmoD23y/4/XBIaI
Ya0xns3oSHqjJl2mw3GN8yxz6KVXVQd4M0eDth6dvkt5Ppf2Kv7V+cjGltUDX25A99s/vPlsJDKp
6hLvff6nP/WgqinDGAXhejo4Q2W2PJdtBOsVdMzgsAM71NDRjpI3fLKGe+TI+1QOn7lMxoz0txSb
iWqPfCfoARi05zMj6HM5EyNQxEp37zYuBxuhdW5bExYoEQtuo6Db4hybboGE/Q11El41tLIu9dFR
seGQSA5fLaMHoRor8Q3vDRrsv5n5ft6ecXGvAsZUvVYyJNDhcp0tzgo+a58fpLQwNOdFHbrKP2H5
zypHlLDOKFQA+VmoA6OvngLKdAhS2sXA6KznmvNhj6z7Mx9j4mFdwC+3px0j1SWZ+ZPi0oyjbp2Z
jF3paWDLK+8V1W3uNXUs2Iq3Gd/p8hELCzTLQZoI1Gynk0PfHWNAO/8EMUxbsLDo//c1byPXgzAR
XaOYy4AkL7w+rYkCCgsiERT/VAVp4rVQrWhS7Z31ZnPDQPhqdH4VS+1DLk+TiueF64M22TLYuKoQ
XAyArpGG/sVdTyjjBJSdP+dohe4Dw2LPNfqX2GOTd5N3+wtfoj9IqXPROMOiaL2ByHUtt+/S+WIC
jbei9dMW4BH6hcY0xlub9Gu06CFBRYE8b86615ejEWv94L6dVcTs0u96BLA7vhbYGX19WNaEAHUJ
gg/KqHUkgWPi/X6DdU9TqY+T+eBnXAle3s42Kaffpw2SSHsA6m+r3c4SvG15w9mn9X0/bZyMH998
m5FGqAZ6wP2YLrPnMbVTXCL631okhFBJW6G1a5ay7IBTZXbnUZdpw+45XP7TtlS4wIDMFxDvJGMT
q0Zf+NEYVUIeaYHqVWiTPVG9T1Zh9fTzXHUM17yNWbuvrAn8GMa4jLXmHKBNgzNr/2NR1c4HiRGC
tjnwlFiEqFdzPb8WS7h0runCmTaOjZZdYDnPRmkIlOCaXbWEL3kUrHAfwjZaOhM20q0Oo4YCkLOU
O5TB+ffn4PLrl/rDwMikPNZc+3FsBqT5rgBpwwOg0EYw3l4DZwv1fGyG7Se50Nzp+8BOwG1vSzhF
sLVf8CF62dwiCq3Oy5ITXQuK3nGlgVKsGc37+oAAhsWl/9ReqqwiEdPhsyzjatrEb23FWS2/i/pQ
4RJnSLsDmm7viCRCFpR8RHABGvhZ3BJgYdLF6AJD9iZ3KjFSHhbmcLLKyVUeuQLO3EQhJRCHlvGh
CyqwRSJ5lUaxMyabiV7/APnRdRXhsFvZ+xfO2V5MGFZzh41iKuR4DALkP5PGjma6lE1EWjgqnrDp
PNd8eXJp37ldA4ZvKqsUQpeQFnQzBErjo4+kqJKxrwavxx9fKuBefvQIlBGPl0Pplp9n1vXX3939
UB7TPT+XphNXq/kWT9QL5kh6iEmfcwvAwJ0tCVsdI3RIOq7E2ZN9/ElM8/ls65HyvZklTuAMi9J4
jHVCGVA2ZI57LEzqw1E802h244yzpkLcbr6aCOE4ya2QMXZrHcjJPCYGWUdL60V7nsPf1qL7pE0z
CtkX0sEUNtAx3tjdoIuA+P16OAWpo4eUjswHmIlpWlQC7rQj2WdPje8Y8WUEIup8HdgzhxxeLNyw
MGJWE0HiiUhk+srdqOUi/1kC3sYsACHqldJ8WRR6nYmWe2hiyZLAovxpeLfbKNoUzar8Y8IjosCM
Ar+NNCcJ26bqNK4za8EQYHtBwc+rRmqWFrBHaMPQMKuYL2C/8Gnkg1xoe+sfhsTfFSgSIn4CasS9
1hW9PLnwq+iNFWyMjGrGS890z665r+dl2C4eN7yLt0SRAfayG4d/JQPxFvzoCpfma7D+xwiCP9p1
2er76pwCgZUhhvUKhLiScS9SdY/s336ziasE1ouIl7OBF9bcl9AuFSINolKTieT+x4TZDwEHDEP2
ZBCY9L9wT8up/PzrwO8Dm2yBZDnBZUtm7u/eZFCvcPawGeRvZHUPI3Eph2IJgJvHFPKPUKO6U+HR
3ibG94TwI8MnMX3gB5CZigN6uLderv0G7lgrqSWIzViQYdtstQhfps99ZOycFmK3P1+Ph+jUdUUT
NWwsD0V/SBSB2VcL2T+zt3YVV+H2Co98jhdSCQgVxM+mK5WjeBq31NyVXdM/2O3Un9S8C/FpaoBd
+oq8XB2Aatcs9uuY6WilyJ9bZKAHo7x0R4+gKrxLr6NqqWHylCN80ajnRYb2BYfuMXUB/7lotB8o
yUFYWJtcqzvfAI1KL55oBuzUzHzzvAPp/llb2q4UbNn+1ktF5CCGzb3JXhLhCjSwgJDs5PEA0qzf
2So5v4YSM8E9cXIBRl5618nCfyBkPZeUxWPzLKfK5aKD01Lm3cUg7FlXTe0ZwR3VxDNQuUbjAZM0
RA1DvEnMSnfAHZBe6efN1Dri6ogyivq/zxBhL0xAk8b0EK1xz04NEmEEsVdy7ruRRhqJZoWjStFn
3LRBInwrfkhIgb2VCvB+mIa/ojdCBO4ZG9qCXNDCJlIEkAllNAravuqHbVtB/TAtBSEjGPcefL7M
7PaQIdmulv/VPY1b6XqLorUu49ekkUR0yzv6twEVEL2CXvrJkCLByFUA1yshqEWuVPJH9UxoKpTF
hwyE54PgNATmEPvc6nFgJ7Bq8dupDgF/b0c6LSDyC7JnOEcKxaZxUD0jAmRN/jcovMVhd3OuFwMQ
xD/Twn01vRCRpodckbT1STlZ9osUMMduZR8ySwfLzV9i1lsojCOL6MjJKaynOsi16RJe9BYJrtk+
JhuqxBR0bPP/TAI++TqXcP/iWavSqHuXWr4CX43L/d8juBCxveAFDKXMtGSTkrZPYW0CzX4oSfK/
uE/ZjdNwTgnhSsCKkIRumgNOgfPDjShpcPb2emOjVF0ALBQAYd3qNJD2fTvn0/ZlzsQUwNKwDaCo
+GSpCSiw0eu3Jh2l5mB6rGH+88UtOh9YOz143BRJJRw6Pl7redSv/C1ZNTc71vIuwiUO+oEE30lq
fnioE21lHeAjRVXNql5MDb+umOXJb2Rs1jJEZ28om7Vj9J0S4KmzITDhi4duHCsUSHKCKyrowrTf
Ide7KzYCZqLqHFNkRrnzdXCiFshlrMMK9WKdD4cLbIeOmwqX91457caIl3n/jJNgTCrPWd3SJyds
PxNSKn8zuONoijqBKTbXaJzSltdD33Gp7+UakZWxg3qrDHaWsXE96g8xqM6+0+BBwJlf9wAnleju
x0e27eaJounGwNOWpqW5AJUZmlgeoUsAAnXTQkZi0e7Vq8lJX5EvVSqQEC2OhdK5fmd1WREe935U
ErN49/aPypfGHFlJXz3GDdsKiupFFAXinc0Du0O9k5SAvGAIp4ApsVvqtHJaf2Ut8Dod3CflU3xs
mlASCEah6aazoBs0pgWT+ftM52PYvb/+DVhe8I+Ga79c2uLmL5hmoIrYPMTKWFT73H5gfZNzytHI
qYy6ynSPtJgrSPc0U9rtLbB6YzpcQKAe6Bu2vMms4oas6wkKyPRtvcg/3XiSdxSTOpQDU1KqpVc/
vSCJWysu488xJRVXP163hfEBwQnSmf31R6muf4jHWAMxKuyhl584i9wuz+Aa8k8SLQsMHVfEofnm
nOjTPScAAJgXbbykZmtCOGZ4Kv/gw2nx5je2WU/DxME79nFhaoV1gWtKpOxKSdJhDpfM3xrcAT0m
Oome+xA0aSpGrjkdUEVRuLEcCN697ERMAEn0aSUzD/XW7RlnNFmthECQZP+0Qx+MFuD+c67zmCfb
Uxdm20X3UMN+cLj8kOrvYg+sWEZifna5JB/59aTK+ZmUEtJblxi6vDub041aFiiXBcPa8vC6c2TY
HQiIsyoMFPI3alpqiV3fw65ZGR4ei9N1PGUMmpnfgg8mIls6vND3wX9Za7i0p5fqCGj0cWyZuTZi
0FA5DKN5s7AJwB1eMfrn+qiKzjoMj5wHqAXmBxf2TCkymb8kXpgqLVumAjkvtNE7x3qOcTR9yTof
Elwut/l4lu7zkskUGGFl6iRuiByIh081dBp/XE8mlkMgw9vVLuuGRr8RyHmwDfFKeLLlSGmqPh3O
xAhT0mhV02vZlvqLVvvTTUTURQazSjzvhoHUdcXP0fSwaHxLhFumnQai6gSrVIN04130Xplu2Xlr
L7H4vHVtPP+wqExtzOG1g7a1uxKufK3C6PaqRuOGH36yimG1msBeK4Bhn0E5P63J4BP3oKn7Z9ij
x/8pDT+vYO7CDM1g4cxki7Ejf4ZAc2/A7pg5n//gtrhAr3DaH7+T8uJYfmqPc/Qq8eBDVftf7IAH
+LQTNSw/NtEpkdbktYkiwItXM1r3SFrtY/M+4DfW3/wqooBLCzgjVK79pZJCOgCxVByJ0S00kZhy
rR33LaTb1aBwaN5W+BpU9il2NLcqtxnXmUuQsxA9SbbrWkuOuQHBXGjdCsc8SVp0EX3ULyiONhL7
uotwzey6GVOvp1ClDbQlB5a8jjY8UjssoKZgHT+QuPl7CVWMD2L4y5cK1Nc63eKI9veW8chCNbct
uo1pFSV7TZTBWhH+3mVzRkDaMpjRdSemKErRqdKYpkA9/ypvp5WhnhLd420o3Xokd2RUlqvJ2WCl
kNDEJO0V91EKOXudE4Jx6rYQ7xEVdc/vqpiIMjh0E7aB4DKIVEa2yJgPSeab2FacVJShnYVnc6tO
iMEA/fw+f1QjOC90Y/DmxlcGWoxb9iusHyJs63YH6WgcRnj/MTQ7o6mryNQHL03Rktf7N/7CcFRX
/N/cRumm5vDYzn3bre3/djAW3FANo4Q2SHj7T8X23RaOcdaxfmU0BMxi7aG87vnYVOuz695za4Zv
MDJXlVRCT1wjsYTXPQubDS7WIxAlXUocre5JAyg47TR7xYWRbXrhxMGXS4CLK9J8pIV/yAbbmYIH
OnOH8P6Ib4tt9esyBdmBASAmPDfFQ80UYPT8rGkjQgN6yq5ZT+jArAWfY7MYtTsrkydbui6uZfKX
xwAnsXGHOSTTI88QJ0jKZvHomLuLS0peGmMsiqpAiI69Mqp1iRgClxNtsjhu5ieiDH1onw1nz1mV
tQHFrituKnfpJBWWZmx59LMVlQ9DI8S4EHn7Ablgec3DXbuphSF+Js7qWlHYQQpe1IGcdARrszhT
c662oCJLJvDD8/6a11U+/8LKXmMc4BneKG9brq5JiEfj/eLwiJ8pXX/rX17YjclolqeLqytoolC2
AQdUaQkVOgXcdrLIl9ROnrVkRlZjcDLxe3wFy3TmCFvusHXbuXnKh4KmTskmbGdtLwZc56RRtdde
P2NyHli8Sg1IMURMQSrVrMRoCYJEKjez43FU8MQwTEEEGXstGqielaQWPxh4h80hlFaERb4sC9O9
edgIPabcxfBi+Zp9P7JX4MSKaQ4ut2uoplttkd5jeeFKsoENbno1RZ6U95butG2WdJZa5PQlxug8
kyIoauVrZPwLeid+nC/nxmquTltgJxZSY0yNDbvBLu6Nh4ixKCsaAC9WJPUtTiwJc5G48sRzJ5hC
5XWC67kvJrvmz5TpJ335pU3UoLylTlMjRGuCy0coaxhpvHFF43+alpawKWJvqsVmqUXQgAoEeoug
gFiTOMBl3UV8PRr+Vnv+ZvAZcLy8dNrrTcoxx5aNTAvGOHuI7FhKB09WGzh7GiC9SeMYa9D29vaf
fTJyVGIomS6KTton9yvQksHKRwWC8GXLBhTBfqRAUvkBuebq3JKmFchxczWvoEDTRYA/KMXFd+nx
pnxmraCaSIFgecXSDgwQk03VkmGZWniwl23xJcbzzJfDq5st5KdNcaMf6vUEdDSlyeGKPaST4nKY
mYLs+HQY06VS5BRPw/BE79IwV9J+grf+Wn5DpNlJh7ScpU8HEEmINoO3qtbTIycjQfPofljRq9yU
lPGMtYE/W8sXKDXLEs76pcJetlcT1hOuO9GIGiM1rp8dUDNYDXJGRfBYD6zZKEub4cJf0qVXCWCx
sPMMCyOZFS6AlryTGK61Xf68kr9H4ZHdaVkilnYcZQXXoN75XkuIA74rzNa+CffXcwdAQlUrDnMW
iH27EKBo4s29F/f+Pxc8Eqqo6p9W9Mt8Vwcz6ENuiuQPvboQh6XDwcfG/MFit+3HCc4hV02fXPN6
c6BV78lsckULYXNTg6txA+ZFhENUngB1DprOp+U6lZS9JgNcPKr+DCfjZ4CPGDcChnM1ZFzCOhCw
Xu4UAStyZDnu5L3qe1uN7gZt93Mz7SQG+CfR5ezfaY34rAUqM9Jxrx9t5t6Gz4FEY00veC9WBjzL
6/6X5KjLbM0lBgSZZ2iZffodn3bdcM3FO+Jwyp2uI9n99gGiRmij+TbelaeDZqhQ3YsNdimyNzDi
XhrwfUO3J0en5nMrB8y8iq2MOhrQOycs4YyguXBpl8n0fm8DmFL4cRvKTc5cFVpBq7K+wViM1jM/
c1UsquqW0T7BkAned6cUrR+m6/h+giWtnWoAVCv5naeDerAyvBkQrz86rmGPivJmFlnzxW8wBWZB
eroo8HW+djXI38c632nH3alnwnL4St4uPco73Tht20kjXNtVt0iSVqSea9XzzeCG7YSm2dy7eqCA
UNZBBmYvMdf/eIElMMx0PqM+nuEq4We97uk0gU2buWt+5E0HMYBG0QxCacOkgZH33PxpUuqmu9bm
qFpeWuQ7nHftu5l1kYgNaQCC8p3FZuA4w36Z7hUfDAVg8+QWTtCeIiqgpvpp7QGPGrM8zO+6FBTR
kSRzwWaHDkHvHjlcJCQRZYvKatqhyHtuFkNHApEQsSq4TD6ZRO3beRK4D0Mw3ohJ1aycW8PgCNvE
P7nxQf6cwTHTnjBf0O7K8H6h8OXC68x6IKvIGoaGHHiCBYya9ByWQNgUnlep4FV+CHyKBScwyVpR
qzOF8SWZh7EsyiMPRivLQdNL1AEyifdUvwLnfpTE+MD0ifOgQhHXgf6TKJq2dbCdIO8lKuv4htQP
y1lsCwPHmLTWOSHNmcX6lGcwiEZDoKUq9biCG3Ml/I4SyOub0ZWBFti3fsf4f53b7Di1AK5ugnjA
mfdf1j53/LWg3r4bCdauZ9t5JQ0g0032CDkdL29Mg+aoH0Q812yfg9f7Q3SwwVZRX+JnCFLfRTO+
J4EnfSlBwMEOYmCGW6KQB0uPwhZVMPztbjhiFO6EnE3Jciv4d48/lbUQEbnoB5RKMOvQehck9OlD
DMnwfNpQHpTpprVgw93kgZQZrHG4Uo02Pru7sVJM/dweXNHRAeAdzenBBI44xyPeRA7yiSZnQHVV
r1jZyndO4I8eYrRMt1X4JsuyruYQ0SDUtWsqfDP5m0kcls1LHMhFQZ+W2MqnSGVYLnn09VHkJ17x
hGNZU+DCDWgLaceIJMBJusoZ8HFEvJbsTKnZl5gQPk263SuPEZinnnl18SB7WcDw7pAs9csRLVHh
uUb7pjN7jxZkruShwX/GpJdLKfYlSbrpqCqnEaN92MuJPjFm1IhlPkYcxorxpghc6Tbl/jriZ2OQ
w+m0hP6MwFCAG9wZ5lT+SUrvT4zcYh7JSuMI2pJZruQHOxnOVCvGISv4rEcg9mS75JvBFVvePAsZ
A3rCZfb1MmLObSRABcEl2QWvWfb/IgOlaH4Vhzwk9d0EC9kwS/PcYjQA68Wk+30FOtlMC4MX/2Cp
H1b2PXewrHwa3fGsfzIU4+fxdczuLLfyx+eD9IO5YTzOFzROq2Q7416bAy0ZQnjQ+Jb+EF3w29Xt
wB10nBSmynNGtVv3BUMbk99UHpm/YUHP0lfmDZFSVdAEwDkNuj+hXHxNHCuozod/aXT1w69Ra2qe
UEo0dQ/zC3Vz7dsUEHgm2mwtQ/XaEjMkXn1wwmG2zZW/Yp8XrTfnr9xODDweMmRjIrY3q+WlllKa
b8u/2VzAaYd9RvyCYEjnkbusCwUHUO81B4TyMkZKHYpXHrI/42QPzlY/IBtDtHFAaHW+ilUAXbq5
DD+IzTbnxEFPAKkU7g7IQNuslDkB3X77efUQpRu5viko9MJO6Gmonj+2UCzhxeHEz91B7YeQopbd
wOvinI7GpDzA8mD/fvU3KHzfHoc0ZkPDE/xZC8SyGdMaic/A9SmQmOBHJnKuLM1EsgbxMfmog3Y0
O56sWzdkk9YqU4tb0BNlQTOKSBn5Y5rofk4bFb31/CqaX5BsO13lCk3M9Lnt16NKQXYuf2iR7xcr
4ciV5IAaJDCec1QHa11+gQpPo1E4c2iknBbZgJXabFhrFTG+QNfzOhgp99sr/NlWwgonN4+k+fji
wYFRUGVJqsZlUth66Kq1SOz3Y0eTmik1m0CfQ8PjKrAeDm09/KtRJFXMCe3CUyc0yzQlxgKN5jIK
JYkB/Wa45GmYOTyfE+R2mUE0IspdZidmFJnMk8gPRnj8rH4lJb9Oi9BJcH0nf4Q0eOimWlXH4G4d
ZFZqpDQpWT8CYoHC8z1iCYl4yFaTky7r98Ni92/iW5Ouqh03Dy/gt1dtYDTiFUXkVwT230rkemM1
8zxtRvkoDiuC0CEWc/THdzmPT7N4+7tlWg6IXrcnhsrX0v7wPGOd1aU1hPbiF10Eal24GIiMNOnG
bWrV4gInXII5Ij8of1N1EyTvoHBMn3c1rV2CPAO9vu/UI0sJPJZhlJbs5dHTXmZ0S44+WRJT3z6s
uWKJF5TPhSScvPBhJFw2V/IxI/6SiHam48pZHYyeD988gvXQqxsjc7y5Ll/FmNQPfRv0KJfuXH8I
yb8Vi+uDDqjKuX7L8dastNtPng3Vp67JVm7CmOqpHBoAAt3iw5PXJ7T2Z3fE/ZT3hptP/nfWWtzJ
qsgEY2jhnOwJt8sYogxl9X/pTk8jJACs99NZkPmM9DQjbbmvcG8T/Zfr8XntR9i0h7q87oUtyYeV
JpMddQbiCdH4/w8E3TLhOlw/rk3h8PsoykJGyIgOwlTx8eD6GBQPfnnMfBAqYaxYyE8fuVtlonuC
T1e+ccoQcKG52kcwN5DEZSyNHWgcRdIPlnr31MX3/x6bBS6V+z1W7k60/DQRFTxl7AnrrTBwBiXj
P4Tcz7UaKbyFddIfH64JITLktH+y5dkddHNwXeLrHaXrofjcAkhwXhZi0rFJQq/K1Q1Jht0XZn59
rBEXmAMWkEIChM0WTKgeVpJqHL5mrG8PiLy7LZr53q4coNxfveLLs3MWuX4VdfehjiD4w1pMvQNd
pS1T6m3IF3XANUzF5ruQCy6pYQRVMqOpeArdha9ev5wm8FfzIsYjp4jzTjiimMZVmM/4mgkA3QBT
Grj0eAIrS6/0IMN97ZFp6JTwHZbdYvznJxjgX9CXItoN8Gz8f1yX8ruVdE4itmQfhtowGmrUqemm
WH2arJV/htHhOK/LoJCCc9aRf6B7klxz0k4IfCtgccEyO9sfHwwBR7vXZYfPrLMw/GV9wFP05H73
EWd5eVR6lZwsODI0fXF+E+tclh9w+NLMyL57zmvv27ShoUJdbPAndUKPpX6mKKewqZObte6pldJg
FikhW/m9clttIwEKAQ+z6fEUzytmdc0LdRp+4OGo1wQHIesNntG7NaWPmuG1Fphj5W8G8BYladE6
U+jwk/ON8ogKa1KIfGxV2eNeQKsJVCh+yHlS8LFT0W3VFZshy4gWpEs2V91tdMa1zOERgvIIcUu9
56ZhYhH5MSf1yJI9Yfw7PwPWSZjNfsQi+Gr8LRYcHLbQjAxqVAdh2Jg1ysRA7/5iCA2W3bviHvzZ
1Pb3MbAXYIn9zAuCdX0HRM3GYvLcBi6ANIbCLYu/3NbyKWo/5/N8DJG0/RKq30WelBWZ83vkXDQ5
bQRvtlAqECa1+ELMi3Fm7NAreRIwlII0eEFg4C/J9GonakbUE32ghXYCaZnvTob73Q8jsypzd75H
ELUPshnI+aGJ5QW9AKzmr9Vo6xGvS9qBeqNXCaIIQBOFevMSKfJpWBgERmKc7gzIyvIZovYlazke
z/emCV6VISGCxIoGDnFa1TjeO/OLSKRQB3UyoKwHk5+87IvZHihWj2u5QonQkMXiUVk8ub3IUKga
ix3s+kcaJlloZVvDoKiExhp2GqEhw1l3VZaKQ2YOxsHEjPl1rvMUDt4xnJyBqo9k+0an5vyN2AJ+
kERcmxxWjhOY8pyIT1/oQrC5gEWdvpvBxeWnAs0oc3gSIgyFrqAfT6oPn9LwBGuYBiAJnhSpA7eW
uSZF/gd0H+k46Ne9fhD/dX4XPO/KIfx8RD8NHwXL78qhKd3lhwu0FQr73zpwpOv6ubtvbevLBupF
kYLs4RntqfyW/oRo7aY0DCyK9Vztv/SnJnc0Sh+NYTjgHJXBVkGLAWn1FpAj9VH1aRDO1BTVPdk1
XcMDsjwTRV2FYETg3Vo/GIEQk/CcFs7HS7JOjQ1k7uoIGcuaHrSQad8tAxs4XMJKhDHRxni+PD80
W7FlVvuzcAeg0PXPsP0NfFObAh0JAV42rzedZnHgiPUP/VyQhwpWTxDAehCpnhDHFQvYGhJf/+qL
fzFs1uyvy0I+DLTQoJf/b2nxlGDaapYqO3NeXxaA2XEvHXAdXsAdmF6wEUS2K73E3MRsONU+ZXQN
wXmyz/OBryLy2JA/5t+cht4/56EfhfITIFuyrKxnwLWpn2h6wMcbG5OLva79ZA4IQFGqS7QUW8Hn
G6XkGW1F65J0Ou9Eez0H+5ER57MPhtjVaUtoaz2I+b98ZZORvuUJKJ2yK4PUhLgEAK2p2gbuRFcj
7LD5MTEN2Mkiya+cTVQqDnL8jqbUub1rjr0Nv8eQ3uX4cBypYpJH5zMFUnioMZW9lQ/thFcXghjt
uuNnreF6XSN4bE+QeRHDQP7rqavnelphc3coI7lUmo4UM+JmgwoVt37KgUit/BPLrY5wyzpkwXcb
T32kpVBvw3qGKhBeU9qxnggngA0INqU7jieflA2dZcrVgikfypvnLTHphmScABZWjYDrQ6pBjvLR
/NI/+QI1luC0lb4Dkw8Z7rL0rtaiAYmF0mmpFJ5dZ6yIOdtMfOtvzGu5LUiEBImNzW6xYzqM3BbF
PPue7DiDwDVNbJaeiLgTf+LzOOhageF8DX/esXtL7/YFyWlksMhp+I4W5m3WSE7Dxb/1H4lFXthW
pXwwDhhzpAa1lmpHOXURO1XV3/2xZF0V72Q7pE76F/kY+Ya2LyCeRVW8ZDWc5jIIe2te6LKMYPpi
FsEloJPHNufKkRdLsJ613VOR7X9kcD9KEOi490C8yNa7+uiVWogXgVMU0Nudq2woBWaKqWgYTMDQ
3Xp3s9FGzBp9RWO2A0OsC/4qeeUfflXuRXQWDzZ6lgVK6mO04kqUfBvHNls8Rax8M6dVVfvmGhFG
F94lECJAK794OdrKnPGVjNeqFoReo56nyJ0ImRCnMgnrDkP47oa1u9HkhfbmPQ0JyaEFaR9dcnFU
6Y/41ax47Y7GLb8LzcQWPgNqWl3CZls92hpWje64TqOUJSeue5qFbjEzoPS4jQXW5iKUwYnDPf3g
GOaClPseuLA/eaQ6FTFatsoRpTpUf9qfyZa5dO4KZBRM1lB1zzue9yiGRmgsc2mRKXwq/R+yUilK
f8JtJAIUOvM+1v7ICQpORNBLo91Ohzg1FJUOkBzmx1NpGPxdSn80fHETzA5D5FrHQjQZEpWINTCn
3997E1zvunkR7iPtNZn2GFUgqzjRSSzwrhZH30TbpseP26akxN3bicY9M7bV7sy8+1Z45U5mHIjB
8/l4BsbHbRuR8HRMRJuGempHFdkPb+YOti/56Yj06Ye2GOuOdIRgxKRRNCfmW07lsEQ3BpnK4jmL
N42snHJz4+/A6U2v9RmW4gggDb1YlJ0zO3smZoZsYAzePD4NwHrU3My4RAymeXuBQxkzWcVRiFi3
khiIUPKA9WE0XqbqfmqcjjUm8c+sDV45dP8NegbAjg8Us1C6Vf5QW/CoojgSnEeliPZzeBL6kpby
65FqwbX0fNVZ5k6M7PMVsYwQELdh4/HHE3BaD2iB7xcaBEmRdFCcN2pe4lEWurK/+QufkDzjVnMc
kaBms7HrrvPgjD0cIVEyLVH4WKlbyygKBz63CHI9cbMOiTLR5+hnW0ZV/TPXdTDZVH4OJj9uPe6u
dtnI6Y8H8RY4BigUO1gRc/C/lgKv8LCNsn9+Q6mj5Rv0d97yhbakDaS7c5SmDMsRiDRbsr/di+TR
M+j9Vrt9R2CPxQ1DS3fQdCLNoPCYuUxMdmpx2F8Erp6RN9UqCKVckEpzJoJ9zVN491mw7+3VeHbW
tcRypV/Uud9KoyaZ+5/zZL/qCHNVgoYy/c+vH4okKE+VfItyOxvQ4Ou4Sr/w4yWIEhpek+EEs0Vu
WfrarBjIoQ/mF57/weQUnZoP+Z8S0ALzO2Q6dwJsytb09TQOVKh4Fhvmnp8iDrew3Q9ozhACUV9B
KaYDUPdCB7r6BJD8IYAw2xk5Cq1du9wNK5jvU7vobNOLRQcjaTrUqKVMrFGiYuEdpsveewo/vioo
c/OlSqOIecCU6rNuGvb/GuOse1kbwRguVVtK7sQEBdxK6eaILaWCSQ6BH5f/tIJs9+6DTax5VpGg
xkl7wcFhS3tj+nTN/A7xo+zaqxk0yfKVue/locyyUlQXc/Oi6PKY5M8b0dytK84MHi5uhM/Qp9T3
elvYe8Y3SnqqCQHihe2+dPpHXYo0fwsgYjs/xvZt9P5A2LT1UzOBGX5g/0T/R0A79PZ5BlNNkJny
T8zTdHILpiIsBwrZW1+Vgao1A36n+Ii4kaxse4YLuGhtTdoatJDV40l9zBNM0ORnD/V0mtrLaMeM
rJwJTyOASRiaET8llpxCCbYSLiPszXvkKOZsqAywHWd6OOIOwI/HBB1yA3W9xhKKLD98OyGEHNwT
izq/MD2Ayy2i1HlYfggq5p0Hc4rGLTVcfsfCjmjJB2rJnt9az1YALMyxkUQYFFt6YKmRFY2lfexb
E+J54Ka93MBb0tJCLevg+tS/IyGKNf2xk6bLB/y20awMkLzU0urgK4WFXMHu7VGWlE7Vf3zJ1gMu
ssgEbQePzTjeNB/EMMT3wGyR47u6CuQ3dgg/9mRXNLulPC/XUFJoFxMX34QNdc04sYcXJ11qU1VT
fhO9LzJEokG2hxJWyIeDUG2pykjF8+Ak+0oqFhDokQDtghZH+D3CB5WlA46QfIV68qjb82Ybz9Vf
qUH6Xkq5yNwQn8QX0k0KKMYD0SfGmq83Me7RG7tUDWinnkZW9rzCfTCZHLZKKrSI22lEWfBcfd14
H29p8FXVkHRTQvUHd6V/SwuXdFk3yjM2ZiXZOxoZ28837v19eJSpOIUpHyU5l5BHJOB8YxruRUSU
5Eh3MmMWYuI2jygZ9Y/MILRc1vbOyD7xAzhrdE+uhJd3EB+eqC8Wu8c0LSdoec2u+UmvqKPSMs1M
lKKP68aXaybyd5eZtUeuzJsPbgKU0oFFs+MF7oq33D0uSwLgRgCCgfceCrJK6q9YTvHN0juUlZ/O
Kcq4x11vp7oreKRRglcdeFbM14q0jfQL4zsCxcuK3e04XEicO+SVrcJ9oKjXXSloyw+DdYmoMDoy
h3bX1M/GVCNzKY03YYPEtjg3xC2nVszbhd7iG2MO98kigYSo5b8yHKcVjsjGNmG9zjxamZXY4GKg
Swfm32Wj3O2rulLm4kXeA0zIfyE52rVaZlFlA7BxHZzQ6XMpkzzakUAzasMllW397Z6g+ahDTiXa
iIAcUMGWDEM1g5Vw5bSShKpS5zsr1zLztZt0a6vVGkincf0OxZFh1pmYKFCwdvrh/rtwskdvdgJ6
oG5gzij3B4xmknRWlqKfuCHq0pz4To6VrQP/OlKK97ZxRLcaCd6fPR/ZXmQvNeWm9PmbJ9XVcow3
OsmYIx06ba4ItrA1JyDw0mbk6idxu494fT2SnO6b211dJhSAsqidkoqR4etODAHQfks6R6GyT6/c
z5cr+EbqHRRXga/sqMFhK2RVTYNaxOmFrM894FqFluFnuIPFBwwN4Z46DR1CH8CQMXFVCgsgVmh0
OOTp1WGI7HRTIw2Rm/XAPPRC79D3H9GIm/Lgyq3wGMsXdWlbhDZw17OdVdwm7VXPBSQ9bYzHN+6j
fyeBAt2l8ax+y4cZ86txHP15AT2yjyyShJkgEKrB3nXnHw7xFjIBVylukcGqHMVEaH27qIvEXMN2
DvakCy8nulYUiWWDNbjnUQMGRqb4MlRGNez6y0ZtgRgWn9pHthPsN2m8U9u7DUBlt76H4r+bLRGh
oyHAjc7ddTL7cC4YBSaectmIZbZ5zK/jlf1Un4rHv6E/WO9SUV50UOkFsPZgtk1EtNkBFrb0nS+B
MVhWsgDrkvxCu8WAx17YqSKylkZ8YRgTDGfregvNCkIRip6fFMY/N+1JA8H0PezCM+nUj7wGksGK
0OICrZEBnN8No3szJdu1t5yUsXPx93gpqfzC32Uu4oCKIK2x6Xrwrs4KdJ7IJJqb4ttbAlemGXt5
eO7szUtg0Y+9PmgzMw8JwaJcPHAVbPRvFwO/chqILCd+GbRDxQLT5W9bhscrfg0hOzcwRiothNUQ
gHn2lPizxfAuB2AhMRw0bqgzrXG9jpYIXvGXmiCANIC+WZkdqcOBLMFTf/JTaiI+8s9myYL1u8aN
U1/FDUodOJ6fqClzhysRerCAWpZ+2gDFamRRulJY2+zeLzl7jWrZHzYvpkD8XY0kHEFi9Pd4niwu
0xwUZJyOhDaGTtxQfjKYjsHApwK1KxewN+O5BcKXFNV6FPItc3pQcJNjjm6xNHuAgfezzAWZe2QG
3CSUr9t8ZetA6ren+7UTAHIykMkgfhTIQM03iyB+XNTMTl5fLcgyRKJZEv4NtENspTyeUmWucidk
S5NDVu29AOo0gjDOD3OPsOkW2o+NKjPr4t/7bl9DuzWsiJmKRjHlSviX3il2bqaLweYQBerFoj8r
3BPCmYqr8AMkcroPjvsFStka0UR+ItpdAesAK2kMA74jW2wB0x+GXUcgj4Oz+1OH73V98IeBHR9L
W+WJ7w8aroom11PT0l3eaz8n08xM+12SEie1ltHpo262jChaT3GBd+FUGx3Jw2I5AsB0NIWu4vkE
q370ps3qkU6Zk4VNtYa/nVsR9j++2prG736WfyK74dhG7TgHRvIqHqvoJESCNwA0MUNVIq9xDZek
sEOEgPMQeMDLW/dZSx3KvwPXqzckRF3ux1fMFBlZ+cbeaJ2yq26rhUiEC6yrwAI1J50NjblxAgrZ
N5X21HDU+ZSNGYPTqlM7NbpRpY6iin7p0SYmRwDdBrsnBIprIgZVbiQJXED79CmKgznV8g8wz+S9
dRrZq64uRNzgtbRuDwk4npqLVL2d2zo0KGLQRq/TlicyEdZWpaqkZLlI/5+MOsmyhU+AGNk41vRY
4WI6wY6M++ONZIVkYGnp7Z8EOI+skdsjbRRKtOSxNMIQTrsVV6Z3uqNqW2pp04Kjode9Ru391mMb
wnhG6A7Ek/W8sNaumDcHvxeu0tH69ENKsIMukB9aBGsXYoFJKdlg6I+3lIZ0zWAF8dUISbnH1Rpx
qVjRy7K7isr4XZ9sNcsZVpzHAAeo2321K69Iu4CmwZ/ldG8ofgqMbckpkMnRxICblOKozJP2GFOV
0TNMliKLWN/xG8yvxcdqoDEHU4aFxNX5/eEqw/UIORlyHP9x4WmZOJ4JSzxjOxUQWatKOSWhC5o9
6ieD5Az9hKYyFV7R6Perr99iadnp6nfgRFSX5uRcuoI+HVBgH9Hy5bChsnYF+4bedkk+woptmhVn
p9EH7jRUdjDVrOd1xnOI9Dqo4TwXgPsA8LI6urPPNP/OSchv3aPlCVTsIJn+T79JsvRmi1uWiWOT
UzknypYNik9NBEL0H739BOPtasRz4fuULxHxpK+JFeqbZXiIfzr8Sfepub+fNj4lAB3K91XVoPY0
JqeuLEpnlOPz8WAJbGx2nmD0LdQDjU3ZqVgqHePFgmxnwDF0pGah87j83WCt1beO1Z6/x/s/eDSZ
mwlBVEL9fbqRu8qkH5EWUA1MMPnRyDEj/mQ+zWCSeCzOYWSJ5C4jLb7X4qqVN1u4ekoIaO7nxgTJ
NLVkO1JTdrsLw9HnJGQ732vq8KLcbJr9qSG1Idc+82c1fomn0uOOChJhVmEFCaVGV55uM4UhFa2Z
RKxps1JiKysfMRF/FvBed/iau5Ch1qPvOB3F2Z1B2fsDNRDmBYLAb4j/YB0Q5a3uiixLtpvOCAxR
sAt2tnb9IVLblFnO9fejFaexT6DWiiiMrtx+XHK+qESC/NmbK+fkUC9qUMQKymUvM25k60Gyl/81
ztuV+sZCVegmuAJ4B3sWPQgEzZP/Ap3L0nSu3wckVxC8u04gRje6W7sPmpp8zj/Rm811b7YyJSor
DMCri1+9p2iD+L/bV36TQFnx4tiRGeEvsNKlR+TR0Irl9B/2zyAYbZ6wnVEb/AEAlOwhRKgdwSXt
7yuvIGWHJ29iKlfAY5nMWK2Ehs/0ehmeaKpYbg7O8vd9/SCz6iEApr+gsXSyXkIvKndW1EDYbvpi
B2kBYfBhoZ+7bBkssmZtzS62uGbV0NZ9hLhteJAWNMMkHGVNC8JX1OY4KQK0+S2OT2iTE7ldMdrf
JgMlmXC6Y0rb+miNhJ2RvKspza+Jpf3kjZ874jtFa8Y1PtQCt0YOOb9pwZrZmECKHEf05bUQLC4p
jggbbm/bZrImPhYpgYeeK9PXvuUPLRa2Ebj1krOCpN1LC8FbqaC1Wpw7MTxVS8ygcRKbOk1eu60r
bUAk2o/WpVKOcSwqqEpUz7kz4ha4LCeoPlp8Vf2PdR8MYhS2/O6aSg1cvhTDXtAxjNudQxUVzLGl
Tc4XLC+k50tfaeN8PkEM+fIGWu0huy7a7LzV7X+w7EMmA1ONzd3j02BfxPpOkUObPD1aIolRxbl5
Dd+ICgUSzzaacV/QsOH8LUFDkNUM1V22BPAJffz0jTqlVyeZQMZwwxprm1D72V3RuRBJnjt95skH
vdlZ8x6XlFTsBcjknM6goHXBOqun9B4QkIwa5UOxq4XSbp2+6V8xBRPPLQiesH8gfjDrJvbtlOwG
/wLjrNTmGS4XvJKqVy4VsWs+AT0p00oRE1diJT+GOt5AgjzPIy9s8WB9SztVCXfYMYx5WrY+ZSoH
lUcOF0kSXK3o51rNEFpSDQCbdV50fYyg+rTQszF8q/OGkqjEKL8mWRMqAaLD2PbrEjl4oEEJJHbn
9w4zskNvKgEBuFmS1vPSnViuXE80BGk3ikfm7GEt5FxE4PaVTFj84zXixY1V3XsetvJ+t7aP//vQ
anbhMtPa5cEo2B/9tYLIyuYzCY2Hum5ghz9zf92p8oWrh5m4wqkEHBLCL9dGH54a72OltlPKWtNV
5X+GWK/XgYRKUsBa6yWVXKkemzXAIlUKifo0jQXyldLqbnmZ2txNkSNG2Azzsh/KIcjDAuGNP8dg
VNK9YOa6Rdnvfx4Sp7U9BXNhDtkC6o0OeZNSnVVPFS0rwHqYOO5Dh6hFaozlySorKpyPEl+6gjMr
UHLCy8ucsKqnE9zGkm4rlJuYdGsXP4fbYuU+yd/LBl5Z0b3NHE1i9f1CBq4PXqH/70qe8eBQqXTa
R6ehpEZF/xsVTCujh+GCn5OZdl3a/8leGVOh5gjMmK10SRE7uKTiOEbcYEwhVwVPTD4eJ8YYSQas
Spj/MAU/UkfkmjVLfpNbFSPobSEuxFauJK7D+94MZgIDvAOzsALzh6g2mjmJkldj3GtwagR9t3UM
4F2/lsk7BQhMytUqhnVfwkOv+V/gwX6bJYK+Oq6gh4YojU7uliyB1OHU6OzWJ1iI+nUPr/UJ7dbc
DvIlkvxYEuhX+ByyTLod51l5iDZR43Xv5OmiXgziiDDmQ9oLOb0GDXQmUFw0utmv63/Lsw5rNmDN
4URE2f148HQrXrCcwW2eyPCa8yQhk2vv9rYOau+R+of5dITEYrdWdHAo5jUDvzT69KmbLftaVcKc
tFo8tSB9iLYL/AXEXra1cxUX0t+NEdGxcw1ZWTfXAE2r2ht/QBe0r6woVpb9gt14n/f2CCIiz96C
EKvePC61JE+SYz65D4kqwqJSVL8bWi9Aaa7oUeL7gV+ijXeUVQlZbnHS1bPZiIsTTxMzEKWLjM1K
xS9iA/JfGKGAU5T1/MzNweGH19smdC2yCoTDwqRgcdE5U0jS5YVurl5jY0k5zygPL0NxAt/OBCsI
S5gWywXfXur2v66h5kYzvjNPCFx3+0emwQnlm7qBSiw+Eu2VfMYuL9XEe3roEhZvzkaVQs4UuQTR
2ZKHL1A7UeT6Q8JVZ1mn7z/SfF58PfS5I1jbz7eiyuscNNWYQlaHccaLmMHidEv+mJde8303QRVH
+1gXYb3dQ3/rs6kXvatzQiSlozpmpHH+ugxAYKbDIxop+dkuo1mUWq15c//lJ7GjsiIse36gIp0L
8DDA7+WounE5aqKA8gXj/wwXaJyjkmZDprSpOgcK7CKtq6PT6NMKv0+Z3thubnct+ygt3bQlL2Iu
flZtz84e5oA2HRBFWGCl8NzFG5n5J15iZE0FTia0BsGSC3tZXQPTeFc95npLp0ZQAKD+D46DaPtT
EDgzQt1W5wU0QUXrJg9Sq/PHm9IM/WwR4Dpd5rRzIstqkBRigdbJmf+VRL2n41e5qcGPMWFvjuQP
MqyhEzUk9aLS+vEFpYQIsFuo8UgtGzGIkiO6hkgsJKPLo7yO5rhTc2vZJsO+wFRwAr/DQaTsZvV9
8Ayfqrxrp/2yVN7DDZhpHbJ3qxnnczSzrr6qKsR8rAjkuTAgSRESwokBcndRo30KC22PJzFvMLhY
wg4GGzLv+5OwxvZ8GMWeTTr+2/OAFidXdWbAnFMtak2prQzHLRqEOSMu8HZEm36N4zJQoQ8+829M
yNa1BHCeMkH+XlJDm92NfA/mBb54AunbyTptza3kaiZcVATshJ/LZzLdmyg5SLohXvS8LerrRtad
jVs+hVaW9zD3Uf7HmLj4KQZBvQs4VeVrGrnnMQLjprA61qiWDOiyNlqCABx40viq6qHS1VVU8HN+
dX9TP26zFtE33WiBLyN7c3WRuCS47J2T84ezX0vzTDzixy9Xu/mSbWswWwQlNpVcgHsDsafJh5gZ
wQHneVcs1AZa6bcnqg2AUbZ+NTDgUM7Ff4I5+Ey5Lv2imiLUCDD4GF96WD40NnukfycPLmE0Nch6
U44AOHGW261NFyEcdc1fy904cXeZoxfrK0Ttlurv8ldG9JU80xvdSoLWjQ/kVbGMlAxgLFfUxzrq
VQdxfmwSRB/pCtRc8WeBHYn3Dn5W9p3D0JxnWRYyCMK7R+66w/p2K5B5MvYlUHjnPqvHexxqZ3zF
GZUkZaTdSm6yl/q1JnjgPwtFVY3U/gdwXlHHlSpi5oysHsE2hbIX6EwiGH2lRo6xl0aCrQhRFZie
0joDc+jRV2YNse5+ouzm+LjE+s2gPXQZKiwIxTQBTQ7XXjWWBBXKvVRQRkLwkB1gtPU55OI0Lfw8
Biq2LmCjOqlYTU5EIaOQNl7MCVYf5DE30FgV72nd8Y9fS9krxfQyFliT+vjoIlD/9OLgcmQDX9UP
5Jqih26NJYfvQQ7n2WIpO/x1q9fERvY/lE56Fls/ieQ7NOH0jMyQn53zDQSD720sS+fJX6P86JYk
AR/cF4uAgE/nirpgQ5sSxICkKiUAbWvJ3zr94ezM89Wm2Y4HA1RrZ6bvFQayib5yq6UvEh1gDe3x
AxC5b3SE3IP6dSC6HgMoDKNVVgnZU/lhrlweScxWOfN4KjwxHBipHax4CecdFegE2YcG4JxT/dED
3nUuGNx5fQfGTXZykgnBVKwu5dhcgne+UfpRof0PB3iBwHsPh6WXP8n/ElGXmA3PSj0AJmgL+6/h
4h6CONkPzHVhYg5vGGsoUWh4JSMZS9JSbNZgMn2ReGHiwYi5Bq9IwKZ54XV/Fx9SAU+UdpqszlZX
iIIINs/eZZ36tt7lX642YznctkUzeS0cfojX+JtayarwXuemt0qUxpv9J2QGLqSu+JXPP1AOrb8E
AmSeKDEnf1pH+ySyv8BYD0fmVRjIhc0fXuG54ZfAW3BbiWrAgtN3CPlJNvNdpcjTrHu0NRTTwG+7
XAyPXhZtbzjyQgnYnTAYOVM/lnpn7Snx1b6BlGooPMf2mOnah/Wi+tA7U6wze4BPjSsDBiKTIBpG
PmaQobd09zM6L+nrMGzfme2NjW9mB9LApmhWr+gGxMpN4GVxxwE+rVzYalokFvO/3ZXuxc0dz3HM
jeRThguF+8vGPqoddBiH/KBAa5fAEM5DM05bb4he/dAFNdK9x0mVL9mXj1/AOTtOGiwnAUq+zKpe
a8kmCjljvG+xTBSIKVvMdPOAKFTk85e048g9cvIBznw/tCaNHH0R6qDy781Q1Eb0tYTX2lBMlcqF
ztnnOFUJPkoXK2WyJQ6f/9r932RbHahkza55aVg84MzgoDHMgje/MYpMECZtqOpUEL30uGUWbigJ
b0b8KcJEtjNTAmJff7ih+KVO46bAcDmH0q+xwz+FfZI0YilR4pvBtnA4HHHrFxPlcIvOrp700o6g
2zLCbEuohzRkeqiyMq27UHZHlqyUHl6F3ViqAwNoIUZS+hsH2YfVxqdB0iVMXB12x/+NFayRByds
00aKEj4cIM5RtO5pQJ04TGf5k8efkWhQlBTei6mL2hEmhDpFv4AXzBWhQ2UWD4CDKxJR/Tb3m+6C
gISi7OfaopH/tJs7Akq1T77PCYC+bnk5l/B+Z4KiBdw1sUwCJocxYF9P+3vierwsOzxoc1xfbxK3
V7DfQfFnmODtjHJ/jpAGLh6bmuFqztSk79hzxS0srqdNgxOxofQOUyIVWJDBak1e/NJsC8sbT91D
3nv8Sk3g07m2/vYmWx3YKKx2nDTOnOhCud7qSaVdextjqY93uFqJjmmfRmPDLk6dBVCIT30cmNOL
Jpgn0GIUDl330PR3GT+t8yThpGzN6P6N5LnR2b3kbD5zCF5m+Vh8W5IXsLz5NFyZBTimvFF0juAD
+Al+Np/tTgxWRg1zstj9oBhgTRmXJvc0hRQd5xuYnlVCoRW1HsojEFycQamT2YFXpJfltSRkHfV0
7U3yNWfw2nRUgaCqACljMJb58B4z94SY2H+/5XqWVGtFB3F8CEAMRjpDv3zhhmSY3crWBpWb65Vt
WfxDrNtgTkwZb0UQl2VZn5vR4vGk782v6wKda9Ft6yHlZGGXJUvNBFpQVgz+JswFxNHDI2hW0Ohr
LI4ooPRID/CvgxFujXmjTBFoJ57+2ssHDX1WY01a34MxqXpiXwAmyQf5gWk8N9yqxt/8J1W+MqdS
b4yoygBw8uJKnIiUAeW83DWLA9A/zbJYa2/vgjGVOp/NE2s3cWfxGYAJPoF2gS23WT1sMxT3s59l
8JKFV4ad06OrWQjBUgY2Nz4N2qW4RTbC30RVR9aOWBY1/LzEtDKinNEZ71PQb41tm/0TJ3K25iCP
2D3qa3TsI9jempqVCXV+N1mHXKUiJUBdYLsgUw+U7A/6ArYtuH1p45MQ4yEYYqjstqWl+IWbb3hX
Q+psiHItD61RowWuRB0M5ROuCbTaP5dKUxh8kldnpoH2AfQmSBA1XOup7Yx8XuGeO9kYVXj1nfga
RciiOohij0FbO9arLv3+b12qr29X6K62UrnuWAkAxPG3hipeTFEdrl8IsARUSX8lq/Fs/c8IDTFw
TMiijXoT4SxWJfJKp96rZwP+Rtjutn7mcZyJv5Ip2vI079UnUWIkPFQ713uK2m99ucvWmys/bTZR
IBqfXW44axeGplopRyQyDdW0hUidq5INYaOdZpMWhSN+UUpIlVOEZyhJFQE+ABOz35BOoZmoPgNA
PhCuXQYWzdWdkMMReR6RUoZw0KY1WMgsJh5Wt8DGkDZnkLUsvBxDHkK2HNnWP8Ji3dBUKQYVFXHF
wSiuTmLV3qQlACuZZ6FCwjYa548qNoQE6IafVFBW+4o/PeLvQ83t9Mk3N13iCRg9wj6ma9b+u9hc
9hO9Z065OBsz0lGzsElgTmIWmDAbfRyRigllWhF1yczlQThL1D1chuV6p8OMN1z6wUcav/RkXOsu
TWpgMk9T2HtMnyq6MGWkZD8kaJrM+c+2jAzb2epzaVBPzabpE6UWh81C9B5zm/Rpj9v/S7oxfKnB
vlhPjMqDrMRwCro9Bk9LR2vh8yEBxRc5dStOrSHx8ttpEfnN2NCBH8+/fcxtfTacqiTK3p2UpT2l
IODydQR6CR354+O2bkVreLBf4MvuEt+W0S4p/QUXFF2NuzWiEuzli68z3UG5NYy7mbD+J+gs6H9R
hoAwbxhIEYoGX2LdJ4cAzbSqY65rJt7A5qFH2vr31suZJ6qITBbKOs3vbN6i6ojSa2PbgQl9sKJN
w8ztUKOUU8xsfDXZOCwfWfzlNVTuWvKyWoqWzicncXfp1v6tZrSU5UXDmFvM8fRidITJ53EGimuN
651P6Z3t6AyiYHEDQxms17OCRwZXmKEwieKS8mrS9FYJSr2Zs4oTtVVoUMR+Ec50lWxNo1RcIOWg
G5bOn2lWQt/Pq/Vo7IOS19h1W1wOhb5eZWwBi91IySKCLdZI0EOIsJw4XQ8ukoYZhgj0iRAqXiVk
KCLKZN/hiLpYh+MrCpwMXI2vsdZFbJGCw3o2FXj+I4dJvfHHLRF1cK0qyj5GDbplQu5xOUzI7DLR
GkYreaFiWdSt3+Uey+rA47IDX+i2nKEeuv9X0X4iZ0ZtCUQIuXA6BAQzhj67/e8Lo8onMQGn6IGI
/Ddwft32vjJMrAQriF9XybDKuvswYX1JBzHrGM1/ZLBwN+Wrn3/lEx6jLBuoHnJOJ11BYHPcIKuu
OawX7dcGGu7ZvDJOs1KXZG07zvCiqYBhJvb7tCQf+8316J735qo+lVl+I2QRh7zCUqldT5g5ZYTQ
shVHMi8SyyUs3UcLyrI4sToFYXB+zUQQutJ2P4R+lKrWyGBECEpd8fuWZ/9bHqfUqCXxfpPsBjvK
sEej50yq2WpPtw5GnATg6aBUWNjC7KvmV8kGnTdf6lRoC6gagsjW7PO1zv+0DmmIVn8Cy/AataDT
ZXe1Uh8Aq3x7sA5hdoB0rSg+BJ+ZTFYJFV2l3lCVxGVUxOTSIFeiFvh8qD31zCPo8uBFlIIRV1Bi
P22HRpDhMLqsbpLsPFq4cC54m2f/Ju8qC1wan/+XTkWTX2vO5uxGHxcfbCHCwYcLHBZ3M76NGbOh
fk/44rUs3T+ruYWcHMuUL6069U9q9uzYiUzw6ypibZiPLG9uxj+FG81DQA0duZ7y8rRJPjgrs9NU
Q87p4NqAr0tUd6Aicn0RbfiUXTGAARMiRAkeYzgXzGE9+kR7PFXAPpkyULL2MkaF2rJQogjof1U+
OG6gagph5Zpk4OfVPbFfO4KN1QDbRtqldKWv0PR4a2WmY3YvX3pvw1opvEdouGTYGTzrqy5ghOHE
MvxWxpe6uCnqCbnJi8gTG2lxrUCjW74hX5ZFxr7wKFLxCKBupUsTO132GQx88JGHQuGx58rEKHnn
ZBqDOIbDqWm1LfiyCgSDyr7Z4sI62z6CD3XZxbjlnIduCvYDut6gjZD68PS9z3sYsIfMN6E1iScy
BP0odG+MKvyxL+fBHrVRX8uOqs8HR45aKfj/U1t+x9fp1wUttM7RpNUap1d4slK4yy8TI9IEchzl
Xhxhm971EXWWfYC824dJJQR6mX/xqMfZLaQj1DaERdTAGNPohOvkswa4DT5IL4vFghLtuR7XFpM1
hXHZxmkjR0vKj8qdE7cf3p5Cz13yU5iDsNb2nvsWWE7US70/gqolLXNj/83l9rDdqDSRen/AEleP
xAN4tJIWrbdQ8Ycan8ub+t99hzLr8SjYsTUqpqDFIWWM9QGsBDSahVnxBU3j9pqvgly2YEh2twBm
96BpET5hdkOQQmQTnGxKCeMbIOzW27+ZrkEhYAW6O5vNOdu3jb1y8poB8x1pZn0Fbx0T/SZPUWNa
vS8+TjUychtK7negtTckU3OYMeTK5v/xWkc4TStfrfqbf5rWvBrRxlsqEODfeL/o6Vab96+L65mH
Jcc965hEa7WtfyDZHMX8ROvKh5nFwU/oWw4tpHh/Vubg9AeiIsI12ym1BJt8JXBDR9jAuTZUrTEF
W2CdxyGcMu9JU0yxLXMDQ2s/qCUAP3SY0w0JSIlHjeDC1PzBCXGfWBShbxRAJQQanvhEvJ5jqlzH
8fEtHx4Q/k5uDZz/J1AnqVI2N2N9+ndL0VkncK88crbRTFWR4f8dh6PsXSq1bHHzZ7oe789B25rU
PaVevJrBZZ47N/3HvwJ0VAJaYyjP9agDJ14D6AOiZTBbuKnYpyhFGXgwncLFFaboDzf1wrpbQws+
CZWZbb0j0T5/0WX0/Og7f9bX6lzFDN9hTuYqwe9wlRKTySrth1TuRvkQeVoWfDtqJL3B5XvcvRgU
o2+jG6mpyA6/lnHVZN/0as2pJx84/2Ufb0TMbk2EfPQIbfgDP6OjrDGTwK8KAbGIyLLH30Y144DM
yQzFvVYC1YQYf21IY46GBKgDlhL4NryyiEXD59eO5p358QkUyMHYm5wlbUUKMEzl2mGY1IXqgs85
tRIAlAPuCxaBfz5j66N1hfs95NggcWdZIIbZ9ZgL28lOBCb16yOag3TZ07vudx1wUTg99oU69Kga
7bIkgydbsxNZrv+ZgdMzoXHw3zg86MBBji97XA5HDxHRa6MRcwpkkobXpY7lP2Z6lb9RMMh1kIOO
yycI3dx9m6Nm1kRqTAxbKlcW1zEcvGwxDPbmnZ6qzehwyb+v7TiFrk7Jp+1ADLdYIbNtCK3S92BG
C1jXWMq3mdK3nVyixx282XeqNxtvH+//Ic3bfpX7TH/SFlrYV1kmtV3G/QVNuy6NSigM3cy/vN2M
yVzltXRzexxTaBgj8FIlLWwbXDjlt4VweRDx4OrXO7ImUYBtxoFeSyXeQsKiejnX6mGhLXI6IsPz
EipcDSLcbBYWYm0cPn8yQlgO9lqjSPxQFnbi1qDflGHVNzBdDKPsjh6Fm7VkS+aBrm/YdRiDnJmf
vfu4zywr5ke8GqNJuT6I2GQ5o/9WHrUp+M+om/XI8WagjLVqGz9YSqmbm8h8eeG5j9OPKW3PAKTY
4sBg4+uuiMCj8cFCvIqgQDB5Nqvm2TOuPe5Az3/NIq+M6sPe+T9+70TsAwTcHonT5QReCAsZyJ2Y
tOIA1riEifBmXFWoyxNl23xj5rKdinSFRsBKnxNq2nVi+sOXyQ5SXKZahpbjhrSC2zFeo63LTGVU
IEJUbyXQgbnk89ZEmuEHI8fc9sPEss/7y2NaTcGl5qW19lki0O2RhWuhcjn4L/b+YDjkpCyyqGWP
WlnEU1L8LWZKKNFY0Nell0Y+QyITsJCLgFFgzFdhsDqkYmUyVarZGhdmBG6BwgIB+tfniBJ+ym4I
40loudMA1ZEUeRxiVKmlomZeBbXCkloW49KY9hVyAXJyg1vdFviO6qx81u+jen7p+wBBiqtCx0x0
BwB70EZHVVBxqGtQ2RK61hVhJp8CNO5OYqL5eu3Lj3UYICVNiVLO7NEJxCaZbKW/5rDzAiHEcpuS
1Q3zteG3+k7oNwteFdnSRSYsyoMyA9b3ujEhlZfgjV3SJV1uVWrDfrOnK2DSq3/A0KTQVzvt7/4z
LxyD9AaqbFYhExMW8JoO84drB/UUBXuI97mjg2e2n0Ic96uuR2qH4pIvaLx6h2wf28uvRJRrquVT
jIghH3RA1g/h4dtaY08jAUOEuUQPhNOdj7Zr7jX9RvaZB+DvCouGTIwjYhNchtmc+Nn2dSvPNfZg
oADy/cJGjdbCgjfSgKsZlRoE0KSAy6FotDp/qKRZ1te9AOkjM4cXEX5cE1uiCPw7m1apGQcta5dY
4XDSqSLgl4HFt0bYGE/jVqNuAQ5PLPFzbQmnbGpe/n4EPdEQEOwod3n2Nre/J8gr98s11TDnOzU7
k+Lt2l218UQn8YaDbyso9jpcsS5j28oe/BRA3UwgXSb7R3r/f4j7xew5T8gk+kaUVRFO0+9A8G3u
fjUoWMu42tfO6TfbVzjZ7rlAkhLvgblvhu77pDiv58VMqs9YUb7YREOA3y33NkTQh9WolYmDIvFg
442hf1wyROJ5NzL2KtGHHJB2tNLYApQDBv1k6TX0zFbCP1WnYr3FI+CthNVotri7T6OG9HCaewi2
MWHjdPW7fijw2li4sxI27irpFotOUSf7LPEK/+5eVtYOeW3/i3ZC6NvBCT0/ASXjZqyArhtV6VUS
A/asDF58oHUWEZ9uEvhpIdeQEQ6xZBn5BnaravJOHmtWChSHZNFOqLQzbkJ0dP/ZLedJQVzsaKpB
/BJaqLg3y2vT1ILQRQ3nDKLFiTYA+AesQk4PJ+1gOo1qvB79VcslV+TELbgPNSgABU+sX/WIUhuE
3IEG2qx0xp/sZDNtsWoXueFXkYD1nZruiv0vmf2I9UfO9OqkLUK1G96VNV5naghIUJFLRUnP51k4
5FEAWAAvn0rVSeQwr5/xpMBAfhPYaWU1Pp60aJV46jVEWROJXZEiKyoWTp9zf4EtdA1XeqNlJ2Mj
yAEroes3DXKLNqlYOmEGTWc1/03AgbV20lqKqNGsGVHVmtDkoTCoze3jN828xFo85QNW1uxtPd+T
UpaANUyK6jwWkrCEMXSQlyxxLjyGz7gbikm3V0mVrt5pdmraWRn5PcZNrLASNTPSJk7J9Vp+Anz/
FtqdfFJ6279RBXDdSaeqUSWlnsz7Y2hoCrq0+rxP3FPogb9rKxaKBlrB8QNFkVrDCLoUlXlEKB3S
20H5GW9sCGHFSTpgTLU9QeRiG+JXdUvBfqR4RDDvPiDHZRtu/3THYxe9Ur0xqnK5yXgVylf2PIOH
kpzXqAlPrN98MrwupHNeRPs8Lc+hUoEqg/Ytc6sne5dyBZIzCtHDI4qdnFhaHgnmOGkitCIr35/n
VHd6yqRKXSLlEyL53wsXejwAFj55BnOJVCj/vxtFBUcdJZxNjBNc/4ooAIyUFx/t7/trLQgXXKql
yzzjZhfjvbTljSjxpl6O2wb8OVfzUU4ZSdmblMDyqDZuVnGxFe1WuRVqu21LOQardWRKJFCZlmlF
R1mF5ozkYEytkXSdN+bJKk4DQRss1USBFIxY9EEQh8SdjiIBYgYJn3Sh5Sk3oJuPiADDD0GHtBpB
E6OulFYz2hp+BOVgPDT93mMmResyZsEB8auoworr6P/m88PKOiTAyQs7hxh4qiprTQ/gJjeI4frv
QZpYdWgZXoFmMMuNK/j3LMefuYhvBmyUVTsM1A/kIlZ0sHUGPSpGAUZu4e+06/U57S+9Ha76T7bH
GPzHEuSBiwbFu3Wy2ORQ/eW+P8B1g3Rsuos+Mz60qihI+SD/KeR0RpbMOEmgdGeV9Fd1gs6rdmRq
A1RshBo0DkwsJrCiGYuMWASxVO+zDqoEj05YKqWYy+DHRmyFrY1txZoLMEzEfigCOP3t265TGP2d
3paTp14kR7kDfRPeWgvoiCm0yQ+EPjCS5SnouCWLeJ4C4n0Wt1Fxj4f+Bpy8OuwyedWYIv70dxnI
rk4JJ+Tuh2v1Gu365KAbumixQ4riWBiDuzYRaaBkN/BSwi9pzXQzU/+r0+YB7L+y9qvxdiBqvDUw
AntAWDgXjjGt/OayA75f+LWE7LWA19qjJ55gxByvPNf8SO3v0z1eoCisLdl24Tp1mm2sFXy5y8sN
fzQZxeFLs24ccHmAe2GC8z4AHAQ5vXHTk/S8+o+eXntdZmnR6IZaYRsYMEyIjINsuiErU9FdLK91
UPyM+EWuDlKR+aESbNUINm9LGQ2IaWfWv7qT+fELhLkx68q59b6grGPdBK/5tiFFHC3QGUQhF7/P
9yhKYT1KjwtwH88viAYGu88XHpD5TTJ0jtEKSsD+XWmHFbYq2Fc8njkR2FLL9cUrBt0TTWEdQPyg
P1T5bcPvcTHhgxLPOf88W7NgXzQasfjW8IR7zg/d4A2oA5B6Z7rVpGLmoqFuy7YwPyneJunel3H+
tWdaru8fKRBKPTG6QIMFn8dpsvPficW8ID7Ho0RY3j1CuHR9vYKnXBhIX3V2NZ883fOKSGPKfQH9
DbMULprRE8vznj0A79SEDBPb4McDIAuwn0VR8P3nqf8gGmSKMIR0cuJ0cfWmHUd2/8zh5Ii9tPC6
CZj9RWOXB0jEKLuAXGpXkHvK51v0pnzGMrlPu4/THfCtea5CDy/u+S/Smd4GZsAzYBSa+ZRnXsK0
aBarRp2WfiL2EDgGMwu8tjZa/R+nZ6PR0mgQ5bq82heYW449daD8Om00nFwqrVlEPBIUsF9f4qbH
I0PqfSiPnl6ai6QKQXVOt/tReMgT5awgL8CsK9DNRygwPhxLpqKdHIiaR6M25z+GQbNq6IsTmM0b
WJGacVqVeBJICn2iFqUNYJFIa0X4510VLf4a8YVNVFFq9GyY0adkeY8haNLeisGdiatUv0pDI8I8
whMTohZvuO088vxFe1Noex+chQ41NfVZP8g3ebIEPvo+mLWnRuRC+uyr8Lf/5eh3RHaQ22NIvxAq
xHS+wcSpUtyArOCSQa9HzvhOwDPSjPnkrHDYUyasziw6ZOC9gRumSwUutALyWVEl/lzOkwzYT0Nb
h22sF8Bp/j8CVgACGqJfiprSC+Ky9pkUntsr09mHC3WFM1iKGBRdgGV6bBmR9Jpex4+8r0R3C5YF
FonVwYrsNJsQlDnKaNE9TpL9rwB3hpz+eyMq7A9xJM1VHufX77yYfenx5Q+CDpU5sFuBdRcLUdsv
JnJiCtR7iOwB2Yh+T7HCMyAdJ0nmYiS39QM3fVedRjjZyCm+XNPh+xCsguwZcYh5zjIHg4VTRj0b
GhhdjoQgPuyAhDPWj6D6RTt8bXXxqLtQhieeg6e7B0cmyPjYP3lMI9KPF3PPa5wCXxFamboE6nkR
LqDNqp28RreydQeJygz5Pwvz1HjZH6xT2o3XGP/4TZ1LcCAqOxkR0ND4AL48aFhsfMDUtZZuXfwx
yVF+E+uaLZS2+a5m51nJNSFZ97QZCO7L+AhDQ6S3GevKunyX0SE0QjwIAKtynHzzjEsVrrcIEWnL
/vYHgkHhtggXyDU0jYEPXVJNYP8FLP0XCQ4ZwuS2MR9rNqAhQQQhc4OiFII1eNvO1WkfNNsjRbhQ
GhT1fKJ+YEKjJGjVUpqGJ441NWqrHiCbjMNl98McgqeDlIh7kPke5yO/uWOESMEJ53kemeqcr+dx
rWvpyvqWzL3CQVVoO3x2niKf48WzV8h8Mkr6eUGXMxwzAttCi9sfh6CuYGxuqNmcLLPIJIERI2fi
KTLmKp1Cj3pj/ZrPDcjDFb9DhxUzl/W+0uOmtoq8+C1Qo9qtEw55kcsevUlriHVkoQok9bwPR1oj
6wZFs9/PT9JQyFd9pHOLgO8cV+VJi6SAfJkQdv/Yv528ZlGeWHlTDCQ9oYgGTezfIiaLvXEIFqVc
6dOGNDw6ydR4vkrloQ0EdPiGM3XJrEUExyZaYJ/TKtaclGpcuoAduC++vaWajpOPds70rkoplnoR
muHpBZAa8eUHDzaL79FW+VvT43TZnxtfNQzpGeR0bz+If7GqD8ugWaFGAv2VPsOS1ZT6bIWqp37V
hmmiWtITqxfvj88SqTUZaC+yCl8QUw4ggU8/Xaq/e8vep4rvCVX4IkpA3wJCFwUYMXaktb5O5FR8
3W5XdUMxIq8pn0kMDKQB608pm5RTvLa3RniC1dpSBfWV95dlZDehaDec/g8aNmktmRxv/t2SLga2
vkGRj3isG9vuXMsO45/e7qZ8nuumvVPTUWIEtp9ZumZ+vScOrEVv8wydREljWHqmTqaKY46J1eSr
3qAO0OZKgVc/KeU48YabSNyR29SDnFgSuk3eoD7aR2Nj1mcAokEhtDEjcWRpY/+csAHD5sn22Uw8
wWe2VehN7GWMqh8ZAyjayN67NWICLGO5CCOTB7PQs9Ola7lFRZKRfiKpR+tWVYDKupNwq5sz31GN
+jWpl5WLSTmLxlrL5az9728WaqSvamFVd4n/xE4C2eGZtv4HJbyfMFsJTYglLvVFDQtWmed8hNiN
w9b6KjcE+hMYVkXMvmGc8TGKkNX9ouJF+UJX1gvI5jjP9RUOtJ6AFqSP/QNM2mutZJZuVSxYLnVw
5EEz12/iNuPRfFwfaKSb9V0hGTUuXBBOZK71ILvjnprRNMeG8H9r7mj8rANrvHe070IIgl3eXZSf
EbZOVnux8axP1bIr38SFJN+DoGVXPOOIhr5VCpzX2gkOU05hULD/J3HP8pdQLqaDYGfrsLmHhBee
rMkK8+Alfoko4Fv3kCCC9unEHozhjJI6JrEDg+SWyRbP4xOarin6p9SycmNOWDFN56YcHoK0dc3i
5R8tKn/tfv2MHE3GUsrdC8472bOFg2++ttgG8550a51pPgm0To3VlBrX3ohGwJGem7IpVjGIfD5j
GI9zj4uT4OIpYXSWtVfkuftDBCLtlFKFz9LyghzEprw2JCRnPQafrc7av5JYJLusRWh1ZFC/BWk3
xYwBEn9K9z/l0FytEVNeDKTa6DQpqETSLGpmxVObn72BVX7r34K5hwMobMEXxby++bmlPTLxjHuQ
xfeEAfSUR5Ww90RaTzHBT8/T21pxaA/SaOoXY1/riL1qBrgnpQZ7q0GieAOp5fNHqL+kg9x4PrCH
pP39E/6DIfB1lz6e5L4JvrluWl2F0zPj4ESbI6g2DV1LWzS+15Gs0jmlb5SUCwrnfqDAK28RX/2y
7nr2H6UY1YC0RCRauAUgQcbmwAXikL8eS6RD+fslD1W10dmiNOPapFKd0PZzz9BFeonGqnq6LY1o
kTIrHdi8ZoTl2gvZx/z+DUkidtxNqRmEAB0X9X7fYruNKVHzyN4Iy8NMkNgqOZxxBy9bN8cX24UN
WHCmyvW0IizGYA3hBJi0B9iAwEKf68Sz8i3yE0DBfemVolHbcV3USITIJRou/bBT8A8zS2ibuwN/
a3l25ZV9IWHeUZ1OV6sHZvftRan7noJgLg8RRqbFMee52d69LLkSZx2rt4SFrNKuPu/FVn0lXWri
tDDcfalF8Krj1Naa3fzMPKNQYAbHkNSfVkMIV3YIpi8cfmRJbzT88QRrPfvqEMOAInaoOFkp4yNP
xG+1M1GgT76TzLHpZnzPCBVuissN8/GiK3t1vXvzj0lpAgRO3XgAvSS08iGvpl8j9fia61ooRh4s
sIPQPAZwB0xNEy053zlcjFBahY8qcKoUz7D7hy4H0NtaGoY1GLCy6S2ICcT+vm9JEJMzel0FOGRH
3F7aFIlDaHphdqFXOOI5E9U/b7oljcD9OGyHD20gQSt67OeoEzsprGgJRGeFL7lYiZI6FdsmYIqo
CHinQKjjDnXMiFzou+td69/8Wl0laxDjowSpHHTSDbaHXgJMe2TpsZVsVHvm01p5o7UA/o+WUbrI
Q3/IY0KmHwoUbbeeLjHozoZglPl6oZuN1gsTD20e5yxLAUaIMerBP0xWWymG5+I3+pcqSPVHJlSA
JtIhU46LD8uia/yWkD/oz0THz9xCUHjodTygK4Du07sPPM7Ph0poa9ZzFRLT58GND5V4x6embMEq
I8MIpxmFiUP+PBu9Rpv1cIDiRfr5kH+4e54YXdhaJ3xGTbna3vVtKVmkUyx4hLMHRXDd/IcqZ5a0
vlp5dZQ5iYdOLI7ubCi7OvjiQQNmzPmemUUoiXacLowjKm0kKLHPu7z+peXIeBrx2zsq2xpCTirG
oBmTUkqGWpNNHHnYar6ByTdFF+4vbs9RSWXgVud9x1HSVIRK0sWLA/qGItFPkmaFntBuZwXw9lpn
MVXLrxkK9vK2FOtUgBV5juhYsXpbW7IkmAkS/wiBnDBy6q24SBiViv0rImmVIADERB6zZ9/9y8uU
MU3xpetgVCSHtArkBsUgPo0JUSK9Qgka3TxXz3hU2ODdA7Ur7+3fXEcWvDo2/EUEhYopFQuiscc0
+L+s4mOz00VNWxD8+O8uC4NhrsKd5BfcWdc6jhSzqLgPt7GEThMmfOijKOyLa2cpkqI28tc/gZJN
Hkuq2TvHBM8zoI7Axn0FOhxwWaVwEpwlil5E6v60Ges4wEvoSXZOSIKAhWQtdxLKSkqkD7X2y2+z
bwlo7M/YM2asZ0gCw/2/3JywWSPOVLYlosjmNr8jHwtMAR0hseOsWjmQl+3i3yHLxVMJ6BLOg3tw
+8bgzENwcTBO0Gp7pdgKA6QLBrQ0VjDDBPv0DigCNdaM2lwLL/zXJyXSak8VpWsCV/vv0Mzl7nTh
vw7GhP0XpM3XHIGCGl2FShBEcjLfJdl7gB2ifRNzqZ3qUUZojnp50xPaxTVjGybPmFSLPRoCQ/u9
9ncLy6V4BW0vHwt/rU5uZ1bFqhTyoSZspYP7e5U/uRG4ZtDePOllCbirVmzuolzFeVHkOMI0x16K
B6DJc/y7uLJ0WsT/xd1gh97PaKAriAAi8eGqrOGZdZaV5EAz6/flumKTv5dM/iPrE57fpsaALmUg
mrHtrNY6ehO/tDGki4l3mbvMgQsPCw4gl9qdQpiH48JX0S/GEJazQrUevXW5RFDnz3ZYvMSb8oAL
dbfF9VRFbCq042+5D9TP2XNPqZCRdTFkowb8TrlhVzeSS6onwMlsMEBEYEChFw1x4oXqt/hm/LJi
fIfpJOlVRM2JhbNr0LgROlI2+8C549vsvPzW/ZHoklCr5JP8Em0KX9LFp4DL5KmSLx00w+5MBRw3
Ma/5mFqLrjcfxzWogzE2zFFkjf2UqBeoBCm661PCsGVHdsymJ0EpddMtO6ye/YEljpy7a05mbQg4
X9mcgtJvqV/V2zZWzpZ8O4mB+mvvmdzdcF8Zz12c+BIHF8UwBe8SA7AzNEeFTssZa5EupirT3SgN
SXBgcH+Fc9k9+GMSkQJ+nWOKr3sC68JTYpN4du6qonkOwHHHjI5zqnQrLQSGmhhHn9rziHqKyooy
H9zJ8FjrBLIg/mcxl9MEDw6Kt5sxLaPna669TUmRg6Fn1oQhEBA06bRJg5d84BhFb1YYEZP210XF
3OqF3yUr+a2zadQAY90iWXVlQMADf8ifp0xjJ3okV1g26Nmu0zoWm1S74c9x+cRrUq+LVtozrwed
+iG2AgMXpYmRMSWQ2v9m83lHQAhvQwQQSP2jV7RYN+iQtbZQv1rzgm6EGG4J9fHDrnGYDPAeVRhe
Qh6AZKckBKv7lUuqT1vNm2hipzgVmwpsfKW70sdZGcGCKsh9esCz1FRUtl17J3jvKSpfQNgm6eq0
A0GF9KnlfWc3lhKVnP+Svf1MRIPJQzGKsDfdDsR5eUCSGLgdo1w/LSw6MWnDX29DV/UzDVEfHZFJ
M590o1zheOSmjXgsPGuETFDsz+1I+RN6usiftyvfUUoPBKOwPuwRtYG0iOs+leyNEtl+HV49i4+b
QqLoesKRDc7qxnqnltS2V0aEAdPCp/EEkYF1LWHuob9KjhE4hH1aZnqMwju4GZyqh/PCG0+qfSWW
DKSPm8zworzwjtoBMsvmSElqUl5qV6UbX7sCsg4UIdgcJfWrZXs3+bbw6Yk7i+YpvQybATPN50mf
RRkKsfyDTxxVU6xaxXv8D/SYmBeQtDGG/VSJfwAOoJYQZwGZ7+/LnO01kE4rd3qvHBOuiz+3P0gE
X3PCTvtI4Qf53pWZ5PaeY6uZiEwNt6Wk2d+J0UgYuHnboPdzT9wTHBGmo+v70axSHR17IwPnR+SJ
SmuufF4kA7xqIqeDCgNfOhU6fDwL0KApSqXN4lpCi/JTywu2yqIntaOr2aMEZ1BdznMp+DG5Z4Gv
f4Cvdq3oBW6eiF5dF6QhbgQfQyt1VWcjPqBSHJpaAIi2Kui3fwb0cCKIRVYrpXuAiRdVQZ/Phxaw
eKqyl2YqOhMS5zP4FNzH2NyWMRfphYIMy0ZHRV5fhvfVkiXr3ZFMSUZp9d+y3kJXg0dqJ4kWDKmY
Z+FlecH/AFGqQrUOTCItt4GjVBjfzdxgilSNbSW/gU9xLON4ML3ywvEI63m0OFEZ6eYH01phDE2l
XG8KGteB+r2Zf/Kuhy6x+OGh5T9Fi5IU2Dkb8+ctJWow133FDmHA+nTJCY4gfmVh76qTh12LJ2vC
iAgrIaPCPki0W+sKJIcOfRhbwiOPMDhfrY1wrTDOuVbZw63pbyL31Z/vEE4LqiZDDHFOfmZS+FCg
Jb7cQ7qOFVHaRyzlAteUq0q6qPIneU2EuwSszYUZfBPpmP76JLuU6NI+dpZUB1SYsuNQPB3Lo2/R
CKAo9urFIL+MwaUL0eij2L1puQLSRoo6CbAJZXIDBWKYroMVYkDIw6yIC84dfkHzqYU2pGe8eT5v
XDSG9Z6pjls8Jez5OfPX2YVgG1Wp0fwAftuoNfnMhTqs+++9YQDwzCDFBcZC7wj5EPXBLMtTscb3
BF7UnLW2Tojnx2UVUPrsyMUlopOnefBTLlYEx87nwvHDcK4mYJXQFk3WZMizXWEHpQebh1e4DeFm
U6BEuG83IDw7xSZAxi7a63xDazuq31WREEkn/TAd6qeBVAMxPaptSfgaHlitz/TptiQ6G0NX1a7w
Ty9ZaHDqJZYS5N3KKdQeYnUNdE0SVWl9y7EkAnfZBuOFuoSHfSpfXpqKpYau3IRhRZcX09JAn7sD
10yKjbjHCJWe0Q1Z062ZhmQJiaORXRDC9IsYI4Fj7S97JZf8VIr9Zjp30LpxJgyxvCz7EN8g+x2z
BCzJK+w+wq9X7jj3H+8BTjlOywJBIQEVgvpmvc03EuW5YUBNVkWff+vZuIwKKlmnFRAP2rkWOWsJ
bmJb491VgM7UkEI+c9TGMd0hqU01NF050o1NB+isP0/hLAj3YduZD3MsgDP9Qj6/exN4YutPZxct
ak2F7s/meDIm2o6HYLjlAx9rIkSp8YUCUrhqQvLUN3sgI6wlQgJy0M/u5jhw3369CbQNFhCVYZz+
n7QXOH6ksrN7OVNA0b8gXHmATtkRQ+XcsQzF5zqz1zieagW/T55uKNxCJDkzPQPnWTsq0EokyNIs
wLEwkyLIau/gDXK50JGM5ZU7hBSbhNMRN2LTRcMB95ab97UI9ip+rPVHolwPiSTNMHV1XsqJ3zBr
TbJteIzy2BLyzHOpv9MbcOdJY5BbozzeJmsdlgYQ8xPjFR2IF5dEIlGUaMsXmvLUl08U/4JZ4AGL
aHS4dQSjxirGu3Jh1NgQY9c4ak+dKUIJRv/Xdx6pafiIYmJ3ss0Rc9Ss5/PGAou5SESqG+c/QUNy
rh5YtFRvbocDLCU24DqtiOmGaxXqAF7T6HbQ6a5GnFubXBuIfD5n9fSb4mpERTio6t0sZJ01d38T
FoIm58pD56nUfv/gU5yat11+yUEEYZykfPp83dedvWQSVaj4T04rRsabKWlBZhm8TnogLlKLzAMx
O8u7ZYy9opN1ISTQDVcinXiQpMTZXJ3AeBxygO2Z7QzSz6pxNKkgeUwtLzId+hEkN+n0BWgKbITu
vGtQMkRTz6Jf0JonBq7lzNsfQ/0QML9/ximUVurtvUbDqqogCPvi1PjXPepi4NzkMhXPy3Z3W+mg
MlDhafD6MLyeJ9the3QEjfKpnBBpcvLgT1MVtZE4FbORv9aIYP1vNgBGXxk0/bLKKFKzUkyH6/CP
ZaIcjAlUBgJGcq5+QnyN0bTvgLb9PWgHh7pDmx3BNupp+uzl072OaOH4ZDYU56VXHBdYUBbziF5c
ghgfX3WM0lBqGdb5pAaSKQutALGKsB5gb+B4y+9+pQhi+1omCgsSekvj9M20IgtLtOK9U7EvefpW
Hb8gDXPrMBIs5G4b5yhfuulVxx/p3G5YKyvmQoT3BaqvQvJbIyVLvpkPD7VJ+61ieOGrbPK03gK8
VxVL8+qttUqucCYn/94oOGnT3SwZhYoW94Qh+yEAK3Ng6fzKQlYVkPYMTFbk5yS0K0I65RAk5LKA
Urjb41ujyxzVo+w1udOcVPzjBbo1ErnSczv+lhJ2Bko2zgEntMwjUQ8H38oXZRAqTTJA/67Rtayd
nWkxrIRTMTXMglfkjHzXExmO9O/AKUXIbtE0Atb81ChBlqQTjFX/vY6Cxoo+Q0EmnALUlNyTamwd
BxWk7Y5ds3tf8k3+XVHWo38L79WufU8ILTZUEEDXQOvsZydaNwZvpAxKvgQD5wLUoM6zeeSpYVNC
r69Jo1GsVNi1VxzDTcGhSK6tEhw8z0pqbg0Mrh+SbuVjluDO7VttH8GMXxr7lCaSg4Tca5wzHI14
HBsVshc4G9VuLFbLEZNzvHWXlwOquoFHX7eucafgeZif5yOOME595uZhdqSizQswj1UlfJlA+PqY
expo5ygwRVIIIE2GgbIKkxvigmxuIK6ZitkG4z+nD6Pvjij37jsNAEdFO+HCeiZOa32nfHiQ/w8D
sf+LvplEI+6KUNQ/bu2+QazVJZI2seU+k04YAT73klNi6uz2+67fQ6dfh3sXTFpOOHsOJtXodcVo
tQJIuKt80PRrPLj2rn5EI7+8MmkT+dp00909YreEr7pR7sclVPQgM6gNyRFQOoncWwEA8Zu/UxMM
yVmHmBn0V1IKju5N8Av8pknm3ed9M4r8fAo9diXlAWsBxfyjhFuDdPd5I+gdBJI1teMh1Va3KmJY
AbRoBpCpHJwAxT2JM/s6g31Y09hTkBdBKLbHJA5u7vtFVE9P8/VBd0H3svbcJIzF5IjLATXP+8ur
6UjAW4QZXsCvfuhqXO1ZU1t4knYkRyuuwl2jKN8sZj+b6ZnHbAqoEoPMyKc97ka16pdcDCUneYHN
7cb+0GalfaurYvcXtkgRmSqzqczYavbol9ekMbEMO/LcWvgIaaLVxNrnCr1PfB5Xvcp71O/bCtVd
kr9Xb/BEOi5Fka7GAO12MRPgBrlR5KiCKxLp/nEbdTjCwUmcy8VNUdRqAbDtWTT4G7PgmQYtiZD1
v5r28jektGfTnWxg764jety5fYQUO+ekiBVrdmwTuLu/4f5v2MPwsmh9DotHkEmIC91fLm99FVUN
7AQYOcey3vFBSbn5GbCF6WcPQR/zAUPjGkmJl2Jv+aWHXcWvpEVArhVP0O395go/wOMWeRNev8VM
UxPh6NA9m6zUREe3Pr2oXnJJk+b0Fej//2tXxInsA+zkRcBW99xwVVwgwf/ETdQS+XIdr6egukE7
lMAfIJm4EdIgT7j9ZUeF0KDg3vfO2VAy0ZQ1nXung+xommTp8tbzuhDQt9KuQDF+fABEs8OrAupI
80zZscZVZNzYKOfPBOaAMXWq7S72YPNk6tuscdDFd0ZXXC4gQLAxQhwlVM0L5Du/nQy7bNAf4wWP
+9QTZAwb7U4jSILkbikVCISz4j2tPniG0QhwoRlKoHu3hcLSRooxu4v0UDgWVBz5L/xu/+e1a8lC
r9KNRFMDJmnHyEDk68O3LPhClns5jA/NlXId7oixk8VicXu3ScCRt3dayHvohJkg9nasjdwAOBQ1
nu9qHoSYswQN1uJyrFf5v1CgNORQYTj3GASnJLs10hCBhLQUwZ5cbbXJG+lo/vu5syq3umJxf5Ki
kLTVq/3mMVhpYrG8oKNcWvpjqrMn3Y+PjPVF7/s1+mqmZ6FFfAGaE2cydUzsWD6HF031u8LIK0Dz
kW2hVZUOdXiNoNTSWRr1uosnakZxsrvg/IRkKzaUKOkUn1F7+a3dmACynV0xQnC9ZbrmJel8cRs2
ONV2Fveqcysc93w0WACFmyXOla9wDx+og9Ef9uK2lAeGFMRNSWk2mnjfEyVh4itMHYxhzDi4JD5b
mCRK3m13pakfxrNR+JE5SODfWFFOEA6j3hNrq+bjyE5NXbLSgsdFDwcmO4k0rjswUHpEuEp6yNZ/
YvjJ/QZdtrP0kHZXjYcUHsWplTBoqLxZPaLT25NvXHahgkiDEdgte4rw2/xTb4kFyjqvLA1Q8hdV
ZRjLBwzeCP9ZOuXzSIZ5soZcWW6gmq40AH2E/RP96u4vacETfZAm1mdfesZvmt3jo9PdctUd7qFB
9dGMkSSA2KQdDsRQy4cNj9OlkmafcTzuewhOobaPZoNECe/N4SAHL72r2PsFk401SY/WxNgfUqQZ
6QoKREBbbAFj1/Qfz52K+l5E0gHs1jX51MqrKYYvKF9+G9WJ2JSRVEojFDVsa6O6WZgAl2OA3LvZ
zHs2pDHiPGZhvMGGT0jj99B+OBvN8PxxLA6E8DAkRkCWFBMnqbRudN4kVzZBZ+vVeFQvunQ9ly38
2sugU1pTGEzo0rEKH3Lsv5SunH+A6wly1QU/vtmbP9KDOOBUDOb9wBgtRDOtUDewfrTF/RHMzDLr
8j6TqIkmnTr74O923cL7KEERx8N8X1wA2cBhRtPhYpyDlzLH6p5ZH7//fScVMbSZHlxw70c2j/lH
ULeXCmS2ESOAN1WDJXbh7HVlAP3yLRH2QF6G6UsSIAFcSmrDxAWBJqXumHHxmXh9fE0Cy6wyO/hJ
u2oAZiWAgvt8U9gYXnYcAkuOmAYvDkTcZdi683le7P+B6beo//dPMQHaZ+4Ckqm5mjSIcRJ8zhcO
BnJxcLBEffO23wsnG2cndgUVNd0fLrYEh1uoy9tEBEgxBEHixX96DcdeOKpex88QsjLDOzXR7ebn
IRtqtNQarkSnVWF+mwEVv/F2WnQs32mnBVH/ddKUg/ZxAhLd8uQRecsESjXAAWgMIfWkxNLzneRY
OdUcwktRjiyq2Lc/rwrQAcfTbmd6GkZP2e4D1oAu2DJC3YfL5/X1voZkw6KgfoQkoK9+ZfQ/8067
vscZvFj+tnGTdv3ycIdYZ9MRlIfOUFP4OmqjsddcR4jQUluJKQ7ijo4394cd8wSoGOeGODgzUNa0
D+Ta9MUr5hBcWx37G5kpS5aFJ9FSvkfPCaNuPs9Mv00lgDNdPxvX/Qmd6n25mpUpmmiHsElywY7U
2AY+Vlhu7SrLaFZ8SVjOwikBP0Y/1y18F8XR2gTV8dNyYwv0Rqckan4ruSbJWr9U7wpXWPbNlmJK
QSmS5YZI0GufzGtR7t7Sv21exL8GZw+ATnXo/Mtum6XYqh6KwdwjcF7pEa4mKV8mndnqa/VkUuHB
dMo92jbv5A9geeL8R+5wv7pKBQfWm54kttIGg7/l2vUkJSFiO8KkzF0I/EHN02EP6rBnfJazx4tM
8fz4jfEvXmIUFa8megVsgwG8OuAQDzKLumv2U5poDjSeI8rcbTKhF9HqPwYo/M5KQ3QeS2ST/xAM
Zsl2v9wiltPmuUm/JNFa4sHrhgxBnvYA+wPhn1kaV1CaV1rOJqav6SKxkRBbocdeGoYcwNaXLoUz
ELnQucGoaAJnXNzBY0Mmwyo71lnhUGIm4kKgXP7zAdaoQYGJqu/jMf4e/Fo833SG7TnbUY1YMTgM
jcNTiwjcNUdsrX6vvJ24xWwNS2+QCuoMlSfYDufLlo3AO6qp2gP7ciEqAYHJuo08Dkr219v4qTGS
9KJ6wCUTSH6WW9dy0EhWuIzEajgb7kWCk7iyB4uuuxdhjU3+43XEG+UBXhumzW54rpQOq0osLiGr
LG8dcNFg+9QCbH1tNp4uafn2N1YgRwqwzoZoB5dNZ6bbandwBdmS+ethT6SUpkPrl3KYPOGFdNT2
McxIa3qg5SUxfkzBxw7tjxlVn1VUCe5TnMiat2JUZu5cdqoBTmkot1TK0f8p1jdBBBPEhnIy0a9s
UPjTWyVMPb3nQuOypPKwwl8gDDC0/HiWNVDciPHCUhvoUp1NcnZchk9QM+ItslsPMa+HlowdDgO2
tZJOuSdE01OIxoyXBmiyY3eVmraU6UzOpvMjXm9lXlVv42YaMUJ2yc48PMN/84zACeFwWSxMwrE+
KHDGfW6jKv9IXq/UfM6BmJzA8GwQ7Ukepd9yNqJHpwoGG5dkrmoPsLcWN4FKc6G0RNx0QBT1FzZR
jc6s070VLUUrEeevaDbbpi0c2Z1mlhAwdKyBJemJ7+kFlvZbV9rcPuPY7j9X2mgxHDi9yb11UJUO
Ezsi2gUupz/Iwz3PQsChmwFHCMcoeWu3TPTk/6NpgZHwAhJGrtXA9vM39ELKNu9c8NOQ8v3tR09B
8PjN2oibyo4KQ/KvAFHKX/ALtVFhMEerRnWhdQUjeiA5qKO9f6is2QuR1yZT0c+m4naVhPMCqGIl
uduQuHK0SJDXPG7zzIFBwZGmwl102ufEbW8i1CNajUXhBqEs3qKfJD4he/FkxuiErJ9OQtgN8v9n
+K+7p+e9WDagwVJcxMweH21ig2959Pk8b6jus+9RYc8PCtJmYbBlbgD9BHsTBCKY2p5sCkyNzDS+
/RmRfk22t/VG3HMVF9vKI3YjLpd7hPSYJEfDBv6yB6rP6Bz0KpYD0dhCcsLJY4PmKep7vhvL0rzX
jpJeAF+pUEZ8QnJqnLP5ugi4rqYNUy/q0hVJfe++M872ES4OZsQ6wvwlWOs5eDSIhJv0Iy6Ywxne
FFe7SQ+4ro5FGH466oEaI6AXEaYRG3x7DPPbcoMIlaxKF6DyCGH/AnjBQMJ0tHnvZVXeAR/bWHDq
dpiRV22PmUqZF6TbitzkdVikZbmVfiOIqZvuGz4xxmsESfYO37POwXfB6e/Tsh4sQAjA50QlYsw/
wBr+wNs2hU9gDxdoLT/Xee3xswZFCzmHHI/fRTFLowCtpjcAcwcVZ9CcsrgFCmsa6m6ZRVR2ONlM
bwo25UnaTT1LfNeYh7wRH4dVXx+uks/AhgIbYQw3MOC2TCxrbbESIfZl7qP70DLZ+s86A/fKNY0S
7O8CSZj7fPf7nAMw+Y72e4vKTrzQhehrt1unCbYmXvi9bh+woJ4FGGtZKr60PDaUF6T7KFZNNjMZ
UNGcinpWOhEdg1JDN/KcqvvOoIWrred6PiQ5SaQt9a3L5mnEflh24tEpORhTrzqtLibJ1c1ich6v
xjNlYW/wJwnTXFKO0/Y2V8C5mJeZvMeBaZt/civnMNdAmvczBY+xxPRcr25QC255FuKz+TD+pEtN
HIVLY6kH8YZUxUXtTD83sTXI59OYVCoKE9D6f0SfPczYwCZowpJDs5v43NVZs81YZ3rMIuug5EfQ
h9Dn5Zj39u2d/qgQSqT6GF+ZJovVuIVC19xMehyy8wRjNRb+vSvCFGE4D0ZyEyO9/k1CB9Q/RH7F
X86UKVKqY27GTVzFh4Au8ylwCli9Q7Pn0A73GfrGFM5n2Uq0BZEj1yPKSbgcb4u4a2EO4ulkgs9Z
92+KpWhIyV9+Woeis/a9aDY9WZEFToWmT17HB+UI4ng+mhaE3wDUHT0h9mycgBtX0JBfiZmIdudZ
9My2DBU8ZDTRMr1cl4nX2Afi+aB/FyHu0QwijvaKA478cOBtGiak5QJYwZEvcj24m/iZ0AxbJmuo
m/fmCOW+VWIOvf3fPwD6aRlnxsYOcLkI8Q0B6vLe9P1QJbcq/v97hNyarZeSaCnChHeGpWVUzb+5
QvzOjL7FkWU9S18uMM/uK8xScCMAAEtlwfnd+gHqk9WfG/FVkJfSRB3Bi2cXPgRR3XOGyBqvaG9u
42ad2vCrVgZIQiXnZo3YG2tKR5O4IQFa1spuMmnHeVcw4DKNvWuCi2vDNAs4Fl+ktClF6wmZKAiy
shAVLAhpQ0sU5t6oAiM8q/DLsJAby7Pcg3oJRfuz/1dtO+cSAg2mG0Tpu4whA8/jisgHeth15y32
7GDrsQR1RpgRXSgG2c/J5RL2R8WM1rvrQe5ZOM9h0EGHfPCt7xnXlOxEWWB24eKRKIVb+jqXEMA5
dYyQD2hIDQQcaXzMWEWN96ZGPAuftEbuxKM6ub5zKvoqUgAnuHTYrU28TSqARvkPKBw5+43Eo63h
lfIYXlFN5om6PBO+JSzE+P4XaF6KgYKJmaRI6JVfkYGI/GS6dBJwwI6NDhoa87EOG9afh8qvAldC
LJlEb0k0ZMlKa5p2xfCGHrxUQdnxgkLXuHNHdDwrsfr6IBXVsHug93DRNrdcURargkqoru9v1tgT
VokifnjAaAZ5jr2hBjMalM1SIwCfWwBuxlnuLyM41wbhTRXxgYVjX01NvfjScPwsRIb3t209bLut
JhI9QzAN6grwhFKQ3Jgt3EB8Nb1jsHpw3sCFnf63Y4M8Gww5j9k3qd+z5W735KFWfyuHyatUvb23
Bn4dXSzbvkBytikA4STghk9O/gD2hPlx9FqVgG8ie1i9eZGdHihFlO0QwDzt0Yea3rcFtE+Xe/5E
+FQdvhBeXbiRmke8ImsguBFhTgILLekSWNNSSnRW17mmsYPk2gC2Xv0uarCvEwnLhvgV5J8/gUFU
PdsZveB79eLB68lZcfyi+xf/3VmnFfV88n5HsFH+/RYWiXI0t5DGn50uIpr0BhH+Cry9kcqkEjMq
f6fkSk6IW7PsvTfrS9bkR+z7A8EmR21cbINbP5HPiHE6Zw7N79WzywChA8Fpx22s4lkINkK7quhE
rUUVgpn6LN+qLYSLq5dUcfODvYGhloHRjxx4Zu0sFP2jCE15cHMLOyHCPA0kjZo4bOFDNkkdIQCd
k7GahNf6YrTexjH9FlN9qbHAI1FYY+cRSYbGyRm4prKCzLmdQh7Cu/48In606XoVP4O6I5GG+TOn
E9sKOG4ez+VX7k/HcD7lRFNCUlInas6NYrp9ZUDoN5LDBT3n+2qfXiCFJXVsj0/usutbGAiIBd8T
ehJn38j604bHtIIpSsoI/qkUoD4FmL3wF7t9gYEhf4FkxIKli1hVgVGRTqxnpLxchMiAZCH2hWSY
Z1ZYu8S7zm8QjrDf1WkTDA9a9H0YZbLHyzXw6w9XQBIREp43i3xG0WUYliEg2qO9hujf5f4MX+Et
O3mwpfiO9bqZ1BkWiSqe0HFg9G9MwZN4VGwWYA5LyXHJsamnfoSRxlLy+1HyiwCOiC0SKG1W/Eo1
9MryHEhGpCGbFDOp9uad0NSHra+gw7CUZGqGTNYUcNToIaOxrtKvddq0Kl9GxVk2Wxjn9JySARv8
df0QjGpPep1ffA1I1fdVi3Z0yUvIXbqO21MAjcmMAqfyeX0WGleqwYPhpRAmg9Y9Mx2/smiuig7I
XD6qouW+08sznyFbyGd1ngXaYiOAVS21P+L9gj57wQkHaVDRoR3E9+Tpke2XSupCY8UXuAZoclJa
Llajudl/jbSyTnNae9sMjC7TpQsd6wBS4wl6ChOiR7wzy9hr6VUtntxgXR58OXwmwbxcvir6CMR/
4qkJudKhFPJleiTYQmWSVRyCBPZSIUUdnwVLk06X9kN4sxOmZVblx062oLFK+gaStJ+/B0SVpvQa
X5Renfjd5dd0rOTeSescQCX9XM0Sqmi6wZRTTkgtM0YmQRqi/mKwxRFA23EMS8Hfj0RhKkZ460tu
XWZVXo25qCI8dMh1ljKZrwzTwy0ZY5esJd8nihNvbdACUg7LA7LnWEO/EsrcjeRuhJUW79q1dRBQ
uRwXiUJcpiVa3VIy12KGRf5WsCEHx1aebi1I1ZP38j2zRo4j6Jkqtjtk/LqTYGlrNdYza+lDYxzC
pEoguijUKgf87Hnnea3t6xNLeZH+lM6dTwtvLXpCTMCXEmbES5bb0jvWuWlP40AictT25rJ5GpQs
chf9Izc+VeydmyzKhNWN0RR4Vr7cPzgDH1LwoQhAjQbqZJIPt11xEcjz06PmGxMyHtX/2UUUucB0
f1AQNYNcjgwExIeClULHoaJ5e6eC3csNfmzpeF0WNwsUS7wGR/3SjjO6K3pKX8fQ7F+XOAYyU9Hl
ZGoI1VUCpM6RG+cMLg+nyA2UpDLMPlTGERFbn9MwuUZL/REYUijpITl0jCI4nCLeuIE7BKZ79vTX
hk9/Lcmr9j78KMSx3zfLGfE0+X+Uy4wE1WzVdcWE+dG7L4E3RnTmrwGJ4+lhaGW/qnNHvoba3f5H
sX1VZXE8pP0mvI5Jd+oWYkJ+jcOCkyFYYxjGpyPi0TbS6dCKwgazgP1hjeyPIi9VBOJd26K6Aita
bsXQzMaL1ubnkA+6eOV2lKZo+J9MTGeSxU8jccfiOIwzZA3B7XA1x0yuwfRL3iznzN05vbdcMGRD
X03VUlmIujcujvP/Ab9AcEeQz0opZeXvif+7p6TxoQR7aT+auHnY/Q1Wzj0XEoONaHxtTSCIFwAg
A3F6hk3UcUpv4wbwsl5/H17J92x3/8EJXzaJzQaM8f3tgIVQTknV3eJvG++OuaIEkZt9wLTpHX8y
jT3Dc1IBgaMlG1xlCNJziWs6idJRlkBi+X+wV090Mmz07v8SgkCIb8Jov1BLeICn06wW23fRQZlK
bBotbNuN18Ynk8q51hOL7phOQHBxhS2bhUyHqH3q7mEbxBx4nw769OjTcp9Jy7QpcLEGYdDEtkGT
Rla0D+dYpErr7jdBkTs8Uy/UmQDVjtpMmNotdHZeWq1zQDgOjRpEKhUbogoBcby5iQORwTqshob5
iroKfRIjCFQe9quGlJhXR7VXZhHWyaDyi9RqkNFwsiQL0xyopaRsWtY6Tm5dDuCHEhCZfnvlpIvJ
skS5y8RjA1kTT/cwzr8F/fY9MF6NMGHW+lXGJWmTcjlsqIfvXZuRQl8bkpIpkmAbz5kmklEtowST
UDTD+mkyi38I6O5oyW+Q0MYyfQf0MP+TpYSTfu7ye26l3LtbkPHVtef1JihoNG8axBN7nrmygQ2Y
ywPjxKnV3xSJaD/AsjJx7yFEDIF+m3lwYcd7rF683U/z+hFBZ0FEr78A1Z4/t4s/4FvyOKUtV/cf
x+V6yzbimQ3aqRNDGcdZASJPz8ibAH2juNXkCi4VIixs8WgkRxltlTmrQHnr1tuSNrUXtxm0hby1
LFc1ALkgWTcPRfaYBNtC/0U47mYZuFIkY0nNeE68tKdgISC16MmL+Ja1uiE8PJjVh0L7phPC/t71
vtqE4XOeOO+VZg9tno7hYGRKPROKsuqJUXU3BN5jTcAtJFKzVZtiHd3UmIstp+DydlZLh9qETYC8
U3/G6BZC8Fuf+U/+1No5UW2t2ZvouSp+JYxUh8EuWa6VSHgL/3vnuZBgQzfmuyxFXoLJGbwxJPu7
s9Hxcg/fL1NYLQVRuBBeQK4pxphAVZ/BoluulGwu0cbe12yuEfxJ5nfdN6NXkRh9j3sOPihzz2Mw
MzRnGi2iLswOAACvYjeKkxuCl/5B46q57E4Od+KPTvtbHqmEzgEfB+FB1brDgVt+yFEJbltyuv2P
F7D7p9rI0/8mpJuh8TSQaZvj28SYRYuUD7+v96gwlYN4ePKENJvvSIyt0cXcAtABbLl0pix0Q8u4
+rcY8SFPrCNs44KI6I2Mn7EaMd++6AqzGAa+H7jLye+kK48sWW/M767KJkpnhv34vj2nZxY2Bv16
KB2akgMUNby1DV6TH/Pmm+L5dDmqXK3pQ9R766EtdlgU9CgaP8JxpARvotBnAipDMwdAz0PNfhTo
7YFNl7IaJgj9HqyKNz9XjJCon0haFtlWIPix6X/fanrJXv0MgBW3f+HV07hFG2CpDh59mb2YH6zK
ezMnjVnjB1IT5o+L189dSZDlcO8eSewgoL+Gz02lz2oN6VQK1Y4ZR+gFkdAv3/POWRWzsCAQ/nEY
8bQZnXizV6HhlFT+8mSAoPwTUfjOLyp663S9LFEx0V+HOyflxRbvhg8l+EC5sQ23sVCTRcfQ0Yfk
0+nDDiF6zNEXjsONwfCUyzibF6Iz/KimH0leIk5LSksd1mk6RtaV5Vua7n5SpOGrodQ1Xvz03Gz+
LiXPSp506MFhWtypmXrGVqI+DCNMYPDSjECGBfTCWhULrc59QRUlrooSUjzxznbsStQaIfFY3EeO
AzATOig4p7hDWVUqBeM1OPU7lR2mQNQMMNIIAnlHqpURxpfZjCuVwi1VolDjKlfw9Mp6BQV4+rCR
kWn8y2oTCvNxbY7d9i/Uom/BBr3KNBEitgy75PQ4yp/h8CUEmmcsG+zLv7chhkNElITcUN6bmCqv
jidY/WcCbkd+cksEDMqw5U9g9COXWT9f871zy615PAtibHZzQVQcOIAEsTD6DNxrZORw6weBQrOy
prWx2DwTQPLOHcBm590BbzB27MxBjSAVKAsBnOW6T0ReVIfesm/ol7HO0780vUf0jp0/jS4BNBCK
6PdVh3Qk9axwj8mx4VfGqtj9i2aM2fBF2becTFEi2w1dAZoLEK6p1RfFNrRoc4uYM4+Uzan7RDnB
jjesfTwL0vpgtdHdDyYYVekvK0cATKTD0Pr8RG1brU1SNOEH4ZfC0/R7AWSv6itTLQjAvfdIDkjw
B2MI8+TFgo51PuAVQXRyAsSHQgav4AQocQ91AOgKtq+jTmubPtz1K/A/vH9cya1UHDk9tGgs5JE7
sv5YOBWWoZx8xoXRbPqieZB1u5KGpGC2xLBy7EYtoQuu8k+WlwxU2WMoW//hwz21cQwiD/EB8rxb
qTZ5HXYjvVhumAXHlOpkg9PCQ7YV08pPL+tOE5/KR2F/iH4KOB5EEnOhBmilSFqXFX+PqamU+BfS
8FKLIUFDnoAaGl5uRpSbDJhmYWaVQ5k0qymGNzD7N+Sm6Lh6dEoj2lRfHOR27h7ZHFPTqWLtv8rh
qBZlZDM1zG+/UoKL4hUs/gLCY2Jf2BEn1uAu7+sfclx9/F/ZP0MLr+RXMnGF6HZvdzzbiPfN3pGF
OJIsXvTQul2DVIgror700H5ZOpn46WcUYcMp84UAFXDb8/BiMJfW9tqs79eVLNPSMI+q3JmU38ae
go1oPDDGUO8eM7+8hKcYRxdPRmU0vdEVBGb0s53oq0nuJJ7bAhdEvcwOMzcqJl7baLLLLcvdLjgD
lVQGIRY5pA/6sSrLa7LHoeerv3bnc+OYjec9r5A6bp/DO28tUNAJoSpwrkCoIkjQDwahH3K8nREC
fkJRLkkViPriqA1RiKfcfHc1ytBW2QegW/BY+cYtkuZRwyeDmPZfqobgFpyyETO3ovc6MkSsOM3I
3KUSa+vNC+anc7kWa3BfF3gmpe8pUO/9HRI1qFiW/Y52tdDJ7pW8KiSj/N3owkt2GzmdFNaa7w0v
VJbg4at/lh0Ib8yxkb7hM0C7T35orNdczuL1mToAsd5IqhTALB8Rakr3W1t60n6sgqe8YM6s/+69
T04w/fUS20YUMAtrb9c9aDNeE2sUFEumJuX3ltwTwouZZuLW2LpGhNxmxFtIt70+qHN3b5tbeT8U
ylsuUYdd0aCRPzws9o2TllcefdX42VPXocMUCAn2XWRt0jwZLI8cfFyh44yT1rIQjNgC07zpyyhi
V4auGCSnVQYsOJGhBqdi56jUv9xucPa/XZktjOkJTxWEiWVQlhcNAVNC/SlVQjoPYDWbagtGtsTY
DL3DsjSHjsmMt4bBiN2a+h7WL91K9FgR/zN/2tWEk+jCEwkUFmZABOAJCaVFYnvj+VWBvvAjBIyy
Jd/WFXUtFz5fFe1yoiJ4Jc2PIGwLGGuNgcpScEX9hym6D5YgB9sLpHvdozn7jPSPD8aeagOju9/k
bnHzTUMpmd/pbh7i17CtWqHhZ3aFgB8Bhstf3Kb6XDRguVXG12YkP9BybvC9zU306/2In8IYqKw7
h7Iolgcx9hUsXDPg8tyn7AwaadcLQZOxqt8bvRErg9XikU5PMmYpo6RkHDElGaI3DQCdRxUBGM8n
dR2M7X0n5zxz/UfU3Dpv8+A7mIeXUz815IXArkIV7lIn9Ooz9lAkPpVehU6gYf2RFJuFPYSgrYSm
2S38ta1IuYAwUemHNHUJ4U3uxucva9xNhPGLTBH0oKcxn6Gh8X4Gsy9xd7cliN9Wd8NdN3gY+BR5
JDQA/GVcIIHulfV0xJYNbJ1k7IdU/7kNgz+28YpY+IHOkk/2xshajyFv5sBMYAAHRFVDO4nOZZ+h
ZlKJI3BvkZBuJuclZbYos7lcpjLZ5Ic9dhUd3hjjVy/c1ATlpt2ilp2XTbWFXc4cGuVVF1jO8jMo
bfGymRajwOQ/5UnMP7exp16K4nQHfoNnYn2EJCKEsNCTdhWJrVDP7O4uWsjKUWMZxhydTg3nTCfO
GGUxsfd7V3NcofDKlLqT9OG9An6NvBPAws8hosOrd6aUiQA7ysHttUwfU7apCYOvOcXT4i+rEaok
RyaU34/dKX9/OqN/B7DRAhYscprxUhx0SewniZqhW71+ssik2qe526/+RRijyFZevh2hqmAhTDsI
+1jP0iVEJAmswtfLIWQ2U9y33Mjm3NCtd/ZEbeziB/+hgLsTwpubUd10KRaZuhw8hmoQ5btErqsR
TcFPaMSWE9SlXskFhyLHqimZB0g1az1OZ3Ney/oRg89YUaHJj9yxaDVfJTJw023io7RiZuXfr4u6
JX05dpzo4CFDOAQwabC68sM2brvhXZzr2nNzJTjbtOdkSZxWbQC1HA5hsKJhNkQNCPS7jORDkoC5
Gu3AEm5ZKdBrvv9tW0oGvok0C0AvgFBgoIeMJSTLRxrvUtSjkdc5XTFynHEntMpaYxKiivlYl9Bb
6X+MxbtRHAPjGw590JUwuY3Q8JiNNSG7QxpRzy84nG/hu6/5y3PfWWb31BwP5YnSXkhesIdfVhR4
C1WzP7oM+Y9Me6RGCrakvpHttCBX0pkimyKeLVTq4MaJzBfxdIpX/Y+0HtKYgGCRvgd6iDodugK0
3WAp3T1BiWsFjuSi+sHPX55X0HRTJQrjG1zvNAhtGahc6hODNItq5OawaPgHwJKnThgdYm2g8gCg
72Y7ru+0m5tI2OaNb5k5A6GrjVsMH5MODphAzR1+L45YWzL3GyWboNNqCgV9UXCcn9HyQqGnBZG9
OYpcP+ctiBxNlHNKl0BvJQg8VOSCrltmJAQcYGS8r7XKJCqmcrNEthr5mRgNS/NrZm35TMfLM4d0
+bO9+prUl3+jAQ552R0D69h+ou+C60B4lYtMotZFUdDEEOY5RcEmtiVT8QbDSKGrnkNuah9KBfTm
QEpas+Mg4ZA3y9YEmZCagBPxxUjkyP/Lx9l7RHRQTlT8a4C/Zme7x+nmHWji8l74KgCJ3i8+qYgH
kx2bqSz+aZqtorGzNUqVlWwC5DFLGiA9z7ZXJZD9cnx+089fTxlbGQcbtBp9TvNjhK26nGf0Rua7
0Lo7ib0+lB+rDTNiSnJC/Lmyg9UlhyuxkeKRTuYmWVmMi+rSRF/J1gbyY6ZyZUDxdWNaQDF2oSFX
/dTF8yyPqT1hYtGT3b9viaW9lc29GJjxqHnawASxqjPp08BQTQt37uSRqfe/vYJ+TH5+GCN00PMK
QIiGP6OZ8cnrxwgE//b+qXiTD0dPQkERVc3ZoafTCjEuzFZbgOAflhW4e99bF1Gm9BfRfEEZnRk+
21HrOqqrNEbWpIMzOUMpnMBttEDvXtxQq9TM4qvdEbXNSnLlzVV13CBeZ6gLCL5XU11Qlrh7j45w
gi9plr2nXbhrqV/SlyRQf/qSod2OwkwwN0Ey0l7rRn456ISVgwYh/Cti/flqwcPdlYK4Dbo/YV/T
twLHAzR+zPjyW9FUx+af4ziATzH/xcinOsQSP+Jcn6MhU5++XO/CT+j3NGmN2EDwmANEVDbDztU/
lfnHPSTpvKXvXXM53jmpqymI24VBCtl/+Mazfz0zVCQ4412w19cfFXFYv3lQMeALsOba03XLjG9t
ZkkSXM8fpGRLbDPrEaHKDL2rn4l1EIx3Ek9VI3e3joE/cSHpATxCmwRLF+T+yQuOTRsPP0ZQJ6y+
h0rDosreSpVLrx3T4CkVTriDEN/DVEWNvqz5I8dF733A/+hMuNpVeSLTJm6EMWNaJV/nryQ5k+UA
pyfeeVojUk1+C/kBJ8paIUpIKvgIp/cPkhTzBzODldStGblkaWmb67dKjmuuNND09VZxKTHOBqoY
24p6P5N7U0gnwRwMNZ6CHbjYg/Vaebf8GqGJY8XUZG40AAbZyEtTd9W7JMvNN/Lr5BxDkuiFsW7R
OEy6SUnW86PFTld6rHJLoCcCmW6Ac4kaQZeU79ag+Dh7fxMtb/KzI7SIoz5yPFf1LySRBjkrr4/p
EEwvmPT5qHoaR2m613GNVw6yuGRSNxUy1S/N5zDq2MWENYYC0TKAVqFcNkirwEi3GX0t3jRsCZ0y
SqGFEizaT5MR8Z0AAG8ZZhAXj8kzRylsnwZ5rukI4symX9vrjt8BjO3TOU2ljaZXUSZeRd/QTtQN
3ghhl99GBnEUdEut6DrMAQVqzsML1YRTvAQbBk0Oyw+8OQlCFPQNtTFKzLYf6LehuVbhDf7HlanY
0cQhXb5cdDFIyP51R/zu/BFIhIp36uaPDrerHs2ucI/GI6p6sJV4sB+ylsOr1+YGhXsQJ//2/j9i
TsfiLK0a0S3lZ2EuXmTLZjQBeoTrzOAHT/jMm2aykeywHrGoMqfdneKVTObgnQit0z6ssaNGJxcr
lzNC3O2nxa/PM1aC+BdeA9orIuVd9z+NHLmTxI8fg0XaavjTz2+/vIcn+oiG+4X55riPH3J8JH9S
jptqc8X6h6agbFJ5Avh4qROakjMwDfi8n7c8UPeCJ0kGLDN+wcUytUfb8ZB24kJFUtXFEOPZ8Rko
bT1FaWJsw26X08WVqFFaoQhgktOo77KaobRlSKicLbz2n2eAsEan+Xhcjin4ARRSGMstIGWY8tc1
M7tTH8xYJJJmi0BekgNLRQU+D1w5hFY7uwlcvuqUmCsu2ffr4syKk0OdYrSoj8tlI8DQQZhVb18I
F5Eat2wJnE4AYmMMJt/elO0HXHSIwOOYc6GO7THNM9CbJnCKXFXXoOuLV+pHu27ezg6BvO0eghir
+IgyrdqGKs5PS4aD54VoHANbah5Xnm/KgZgtnEWY2iDphfRFlWRMFpdwKrXc4eP2oLIlO6wMeNpv
P/HGs+PtijF9SJIG1juOZYqZtpKwXsOf7oqVEe4AusAvquhvHkT22W7S4SyR7F8aIlgv6orIhLy3
d6i3jXN2EAf2vngk3vEMggqirZ3XSIhdXPJ3GnIXHiPNQgY2ecNmwJ24FVyfQDtxhmio/mvpnSic
gn5WkJ+UTD5xkoowOlDuE/Bm6lMQOegdaqccJ4EeEd9U8twsiuzM+BhT2b5xispjZwkUZvoQw7jZ
bpo++KySsAIj0E+APcrMXY2dgBSwXdz2VbmIhKXBnDIZ0vQ6O78amFhG9ofxaHO82LQq44mz2AFg
rTEv8IvhBNoZ608uEVbpAxREUu1uKh0e13XHO5JBcanLa3q0RaUtvk9taylVOnhcy2B5rvBdKs8F
VrTdcLw0rpHmIsAv0X7y+bVE5ygqqD31YzDImbwII2qh3G9KUj5z7RCxXt8l5hCUMo/6y37TKunQ
s2VZf9GFaNkxRwjDafsHCNJOf/9jMKhajgkQZ47dJNfHUBHSq6Id7VxmU/0HtgMinroDy4s7NhIu
NGNiKYktE2kS2PObnmfbvs79IbC/cx9vztjXcxE4ypuQS/4P4Uv73ujn/gDUvABOsh9QKmFhmbpa
U0F7IbDS97r+7OS6cd/z4MR48ZohU4BOMVNt0Ca/3Dbsr64XJ0sSh4rLvMYGjqSUE8ghhLcqTh6l
rfJz7pYLaUkhx7XjwGicqEbORAEO7KGJZPbRnbpyTckkOHKPkv61MEvl6bTZubETQQ19sJDcmEN8
FeBDMK9heb8BM25CRGv7SsT6YnU1DyQKHI5fg6by8SJjObfd2i0AqMqdCtykyhK9XiFP0wx+CYxa
LPyr3IebowaJ3TJdmFxBk6akZu/6RLezaG9LW+HXy9Y1oAPqXLSw+o+jKEE14ft1ypp63aHCi1YY
4MKF1DwhvIXRJ/HkC1OCkhPKF8+2zU1L42RFNIDZcCx/Ki32M38IzhYV6zheqjgrxqdfra1hzRiM
9QDfqhbd7zn7BPljGVrq1fG74bpiccddhvih4zVR4W10jzQ+PocsyKC64NdJz2YZvpmz6W4fw34t
tepgyVsuDWQCTSwNNY/6SLZB4vRB0ICiB57RyOJbKw3bBXfPTKPfSwwypMd6ip69DSC557u7RYPL
G6PUfVyuWWmpnA8rU3TREDHJSXjJikNJnXgGgdNhYcOdYvKyqiYpdl0MnNTJauKBtxSVu0pnV3n8
qfZ6v5E2tSibbhZns2LQx2BAG9yrUw1uL+N2kTn5D266Iuj0p1Ko95I9S5ICxOLgMmt1JZV/0oUr
3T93R/rCLXFj/NqUuKdmzTouoN0KPF1nYyihSSC9eN4iNyy0GT9talBn5CiGBCS8yaxXDWymSffC
e5Ice75sIlDYTDEYAy48clU7xV71R/IzRAiPdSFyQn/j4GxV5wosRKPMmVHBGfxdzGspeLMZlfk0
u5oEgQ2A1EkDiR2BUeXF/NUvILsDcXxZuuHgqN/JgRCeahZp1Wiuv9kUNxVO9NWVIsw1LzRANQCv
VesS+KlLDaaPyQCjy7irxbL8iUEe7OBQVfRplCvhvOXDQjtoPb3LPrbF2IogLYV4bzsBCuIyqacI
MLoDZ76scDOCR/39HoLnAseZoad3j8ElQ7nWKMabXolKjjz2m0LHhCg9AGompD+zPLxGfapmil7K
9E9IF9vJGJu5JA6+Q6t5BK8Gg0KXTagVzqObGTUpXnRQyNdMWmyBPx8ynoxP/r7Yx7ajin1QtlnS
h2jbmPqcgZLPPErDqO2hZ9EgBG3D/uUKB1ofYxmUeVLnDWJY9CPeNaVfgNIAb+a9c6SCnp6sNaRw
M2UuIRwBLOjFDF4Pao56ZeEI10JXLWujzGeHPFaJyn/SQwT+34gHNKTav4hEvG2fnMPCmjmrXeOZ
kmdA+TIm+qXbDKJlimmCMcIeCLXKXUQd9/HDQoAmZNk+aPehcmvsyJ47s710zZF4GTIdT8xU5u+o
K8n+6bTdiPUpL0jWCZkoKbVMO1TMkm2OuSELEQbhqKVighqIOpKhA0RPjbTM61Pz5heunKaqTGW9
/1Fc1PmoO0ccrcyfiWQi24abxelWo5AKihnPogEQeGJtA/Vt4KxtGh3KALwWH+c1SP3/SKI724AU
RDY+gIDf4zdWq/ggeji05ud5n6kLctVBOwOf8K95DT/qNI46PSVWLzKHRzFwIY219f7d7F/MQuSu
sSmySTvIjvEa+k9fFoOkEUuKT0vJUXeqKZmaoRrDXDuNBUsL/aFx2dcClVV1GLR8WlvAuEeSE3QS
Jp8m0RXTuvWGUvX5tQd8F7QbSYPz6b5l1/d2r0MYEMlVV+NZUKEtVl2+gfeDbJMhmjMwhk2lzuKf
Z2DD3wiv5hQn+X7Vh8ZU8VGJr0uzo++1ic8VgIAakAp/UdJ4UGmwjsPWli84awcrMrOdUV6dqibq
y5RPo9scrdT+PRvCMAqpMrruiJqkCKa1HgUQIrpqggEbhdrZfuyVKxECMdEWnUFjD90AHOOjhenQ
qKLaJ/BgWn201rg/gkb2AYCkGaLjstoqPgSaZIo+seCyz1I5FvEi3s3wMAfZAriUvDgBi36tNUXS
UVS4evDQDF4VjXgX5rm+7LU3hD8dTjL88taUP1K6nxwUmYzx80XpJ4SO5vahMqSa9SUexnztqX2L
Qau4uNZVQZvFQJFfiN6iXPEMlEu5u42O/6JVZznwdDtNGfaMbf+dw1uVynk8h1aStPLBot6lkvJn
4+3E+bO4F7KIgRj54hvWi4elI0sRZBBV67qwX/h5hxmkZWYVXewcIWtLhEaBDFS9st+f9xbBokCA
qdsmFWVE5VTxewDxkF+Aqa16LXOgO1UYIICkK1oMcWa5ntQJX3ctDGXni7A39gN37aEBH1soobp3
6YlpohQcC3KYP6DP6/o/sUMKUHRehNePN+cLTNY4VSx9LXtQZpI0XCJtah4eVjUwVmYQUmkvBANg
NuJw7aVw9hmUBFHJPr77oX9DqzCxaUzBS1/g5EmPMziOAlO9Ep40fcVxJHHcHC1YA2vb4NZHgHvq
rqpiWFeJ3FztXd4iYWRunr6RcBhdhywO3ab4C9rGIsmxCIYmk+1tAx/YB4eW33wOa+wtaGfstXQO
3RnxOHBUCebSvyn480wk78KZvW6TUHP1kktjhVys7NNs20i2xcPhks8VRvLDam9p3VmtHo9LZYRh
nlQ5WSC2wTI7VHKOayCJkZnMqxrYoU6TyWwnt2cc2e7JnS9Rayx1VHdF9AKWd7Pz8FrW2xh9I2nB
CnOkS7BK3F00zbYJEZxBm0EFZhLYvpzwf5sHsLu60UvoQMwJ4Cyau8RG2mwclnvz9BBZIfR+rBuY
vETi19LS65z08RTc8ThGJRih8jT+YGjEcqv3bmcKX3r68nGhY2rt0Zlr7q9XjKmYkzYr81jzwM7F
eKROqvyYWiOgC4zeSl8gpCkjQ/7MxFNKOcFGrZqd6zdaaGbdulm1PsLBqfbsjcC+nLcmscY0eHux
X+/j0bqluU6PSH5aeifaApNJkraZXBXJznrfZlRBwzcl4M1OqJinFwtvu7xzBxB5G0r1o2spATyZ
Q07zm9NzgmA6H9GB1+cflx0Utg8h8YFJm74dNTXY07hpgi4/j3V+XyTwvxJ5Qb+fbOpdfx21BkOz
gsENG38IWIbKyjQOvy5hiUhzc1XrEywN1YdRoz9oTv15SdPjGY1nXbIcqjV6MuStwXm9cVo6/dfE
i8G51U/M56AvoRuYlQYJBn3fugMHlHJiAgXPFek+zM0uQgm0OD5LjXTJbd2ncXtoCzB9GlPGoTHb
InyQSzkjUqzX9hd0cik/6qen+N+btErmRQd/kxl5zZi/zzjKm2kk1a+fRDZJEJJ5fIYOTGPe7+Os
Pge7JCnGTwv/w3PeRh+OLQqSrSdJQ1xfYtSIj3Xa6OatqFkoajz12z/hrQReIuQdB0ETaP+kW3aU
FHcxB+aqSHrXowu6gBTv5CeS7g6qknjLnO/brHl3m0zTnmoCg/vXWz/DaP7sTljxN9CDEYquG2Nl
snHDxJL55Ty2E74wpIcPn8Vesu2uRtgMFeUWrKMerAavIQbIWm53SDYgN8fsJV+uAw8O/fxxsNUs
IcCCCge7UM0LX7mHkAWBgtforwxsblmZcx13XI8cVg91kpxVE31IbeVbhWszlBXqkBhGTHo6ObLo
Id0X6X0kzxFgMW24YGk1RgHbDcpmFADyrZNr3x46/GhespxvimGJMQWz7vYiv/KUYHL8F1Vhp5+S
AP0dk+sWGePKIlrK/VcDrMutFm/AiRM6HxQ0n3X6KMZYV3Y8RsOamrWu6wswKUeqQ3M8Tnsx1tC1
WK1Km7zEWTzSP3NiR1w8jTdXbYwKKE+FLj4AchH6igZtbZM/X+2l0ZKUWSavvNMh8HwH5zJyYhRY
Fkr8rfG8xkJtAtQpjPI+tUAdFiL6JVsBWGEVgeTQAx7VOoWk6Qru0MHXHhXb63/2ygeaV8F7feQ3
+h88R9806ReAPS3PTjc+9G11vtq+DOl1lCd1yPOWxl/5gYpxGYOuGMsDsKMVzyjgMqEIQRQBXmXH
4fbkexb5Td7iyZ+cboHJVel7Nnw1lui2RoQ40p23aFmEssemMUOvNTz7PpxB2Cg5kgV1BQeNaiOq
GcSpgG1nZJ5mOyZsP1t6VNE+8/JhJR1j70s2fCs/qI9CnW4AFO+src3J4anQfSXfOQNtiKaP+DxA
3zU7kIEvlbjzPE6QElnCXQzycaHOFXR/H+5FNwOq/UFqAs2Pe3/O9QiIksI580oVJwjeIVZeyu0K
YlzXhClasvmuqtmeo89zMLQlgrgxpYankimjBiuCoyx/VVw6unRKqF772x8YytBh33H3epnlmotQ
6AU3TqDhedmNjAy37es1/z1rvPV/9YIv0nXGB8MqBvbeuG2PLTzb3b3y0nv1oySp/l2aqc1sPEPa
YYDHIGS2a2cH3CQ7dRjcnapfDMOxNZkLQeQ+kawomO57xmZbhIxrX7JtQX4jn63QmKZf+wAMLkEk
bNI8B+AammPu69hsGaWnr0DXyWWFYr/m6FnT6HJyC+Ze8AAq/1hWT1umqydU5wPzDuwTR/XtCs25
mdog2/YenlwXXhQc9/cjAYeGE2QMr8bN7WvNCOhOpiJm73waYY+I1Y9vB/8wmJrrjk1TJ/OckLTx
ZpWWKwtnQskjLx5tQhoOZL+IUop+iK1CskOzR4+jxBvTFodSJZmv4KqWUnnO8AgIOqF8UyWbQmVn
0tk7BC+uUGsw7FQ20v6/xyYs6B+s34H7E3+3ozcTVufjDfqUfCt9y/ad/yKrRIHTndSRA+zPSm4i
b3jFGZMUXWmzmVFwxq5ffzvLvLK4g5XadKoq+tpSR0Wu2uNjnt9H2mLBVFDiX5PRvRv0M2xA2lpU
l7S4WyDO7zp++hIlv6DgxUyvcakNTXPhEbmDLMztm5izn3kSH0yJh9YUhbvrenXGL6lEyng24Y4R
Be6Xm8u6EZoe3k/ppjZIz6aTxq9O7fC9BgM5lIBt44W4cdxx0o38su3IX+DIo8gsfI5wK+f5IJiY
KC3OdLZRUpuoOLZpYFbc0tPR5DTEW70d7Nhm+mpDQqYuPG3EE5tNTfz2c+oKNgrf/7pe3+YIsIeJ
c3fC8gM25nCm/MJfnYxNUpKv94Y2uGavCFXmWmeFskvSX6XuGZ261iZjlOpy46ITu1277eTnHl7v
+ooZRu7wCo3gigbwiCdxom1oxV9RnVR+rPphBH5XO5QtEFSXru5ypRQ4yeNSkGqhsphHHNRjKCq8
HlZmEFLYLHseOtYgaAHNWF83pWjras4buNW02ms6bN3FWKr4CvXxJw6EmAojkN/m4Z9dHI6t1XEA
mSy9uTvohAVwbXXrQjdAV1HfAPAOnjqyAS/GPBKmrWWetGl+kTA7M+RVqVIdcFUHL0W4wY8EwkPG
TspUosqDE7cxfQGiYmKW+OROvHi8oPG/dO9PwTUTigWa3gacPdRE/QeOTjPRauTpPp/Fjdv0BqGC
jJ5N0tcRdx6rwW2GudLYhi7LIpIjbnKUQjXdlAGL1X78dR+/cduWX8K0ceXjjbzMAJWrv3HCodeW
Nq7DiHp3SskV1FWLK2JiDjNs9tnV/dL1qXHpTK3dP7jLs6gNpm5nt9uOnyhJcQrC3B7zIxC/r5Sf
cf+ehJdmfsKs98yWMSwLdKwCQQ59Bq8acPJ4WtoxrW/QOdkNaSyVn6gBTz2eDxK+aagxI//7UjI4
Ai8HKQ1FCKnBsqTWc/DRjCmpcHjJVq4V2QVukTOLAxcK84HZ5zbx1+aTReaZLwa6TJgY6aObTpKJ
wxGupAtGct6s8pj6+QPIS4nKDyrRYXWzZStsOqZLGsRH6WDrYPbBCJ/WWaKxrE0+/UlomkaQaYki
B5EmZOyr8/zV6qMaE7mOME0sdmXLnkNP2fjy8/tZVHZv+l/oHAh1SqOP4tHbFOYRmdfTFs7Vc5Oq
puNYVS6D7/AabM36zA3ZT5fBjoccStnc3F85Q0D6/jyGBnbOJKWgtjoOFjF5mRwfaUpppcDLAku1
L8YOqvqIFzHEb4MPLQ2tnEBqLdRuCPpZrX10Xl4nmnZb1WwPfyDXLt7AtPxCo2hTTad+TMuIufAG
WD4CrhXWDC6hltRUII/08TSPdL6njovbkpX8vignnvaR6/iSDTPfkof+jmBhLIW1c//b8Hq3hMsg
IA+J5cwJ2Wg2u6oXEmTsGdxgMjKmSRQ3IjRr+kkt3Kwxuz7M+oNrbFmWzbJ82hxZkMkWKspyBO7j
bxCgO9BwYcXqJO66YyQh0TMEimru6NcUlkXKuI2bkRP6DbIOMrXfkr+44/AywGPO2Wj4EaVmOiVC
ZkhxW+udGIMWSZjOsIKbvtey+9HpXPWjWCJyCL8yWRkEpOgsDusHSMNh+kVcJJn/MCeAgPRlksbF
PAef+Ldi8RIXxD3dUY4rFgqTodh5G4SJxj4TBnRxCMW0FHR9JTzXf5MWsF8zQ4Fj0DqWrlT503iE
m87zAqsqvcL7xbdCx7mueQFBg7OS/RaJ41AqdCsasF6je9rt6pJ959TmGFJg8x2MtAh+A3AI9qUJ
QkyTS+GlGqlpBamDnzD6yPU/NJ+QDAiXLhISG3xG9jdbDj4/9e5n++BC3bLuoL+mP7hAOBzvMC+D
kHsoYpVEgKdu7zmet+YQOSgGi/rzuVss/tcUG+QRfMwF/fCyuJoMszXQf+3BVllOmtBdgrnXkYMQ
lt+6bcXM4ehyhSVNyagvKB7WdWDilYLVjp/dGMPqTELdTkkjJGm9YTyGVXr6cbWWYGxEczv5VbG0
RPD45+DzdcGTfzN/EaJYw0WVhVnC9X3TIDEMPLPA+GvhewawyNAS4C4Z64wI648ifj6v0upSCyey
wTbND/9M5mv60/G/euoufesqEiNwIRQEX7Ve/02whFs9a1uLXnG44ysSE2yRLEZq+bhMqvu0EfcC
a1lmrI16SccTjbWJtbTSbpEBC8XxPydE6h8yM/N8hIV8dycGOlHutiUrKKeWA9XoIMIlJBFX9/lL
D93uKr1CgVho6m5XQDwslFag1SIrFJ9kS9EsxgehcAN7iSJhfZbtTyvJpCBSwEBTa22uWWiLTW+8
TPXnFwStlQirQxMFTwQaYNY0CluZb10B06lYhunMGuTalPbK+Bq55XmAPqCq43zHgEM+zaslCxvJ
9PJcRk6Zd2saYUzDbFUDlby8oyzjHHbkDVjVv9zT8idnSiKzcQ1ObQLQRuy1wYWyjnYMByXoU4Xy
QO9aRwCnxI/v+1GwfhWxsIza7x9nl5SkN1k3AM7eEMMHi0KiTrb0d0PBUqIFEOGVMCbHt4VepO7b
n9GHSrY1/FVXR302uhIjEH0Fqy+xBfgSCZeJRW/e1QMN15KwLQc6l2xX9YmiG2Wu2ekY7GIzGMJ+
UEedpFk3u9oCOGu/JI9p8+2oHqc4g/Ly9rJOhqb+XBVokPHi4RpBVf+X/e2k762Z5wW7rKO1J6OO
Y7Gj6rMBdtQ0psZW6nJXnaENoy25F6+HKjFcs4TCNj/z4u/EhhcQKvb/UjxEIrzv9TusXRPxo/D6
v0yOoPqxWL7rQ7Lis+343UHhV7VrmyMj9alorfxof2yQU6qi4Sn4BUS8KOfx8jH3WfR0QLmhXl2m
ro6ySSCo5xQ9iBWYEOczW9Y6A65384h2KnOxymKVciJ3rMZTI5dknMww+T854zj3pps5atxRzZUn
jaSkG00vHYuphKdrLowg2RlyU6dDg0gS8CdSaDvceV8LpfAJcXkGy8JGjOzSU91okjZ23coDlpir
tcb3OZzq6SntWcmNmNrF6Fy4KT6rfXoFa/alVTQH7U5LZH++JGv3gOJLeGVQOFSBmhYSTunnu1Ui
TSkZRH2ijbajrQceEPSNeI3Ot2ai50/IjQXsLW33zbI+0aWB6Ii037KL8iSjvbLbkPoNx/LQbpU0
Z/R9gPrXOMDVTW7yfK835xRKrXbEEfABw/US5xsdcmW0MWFtlZaPSmPSfUs+/9gdVVgG+DA29Stc
aseti0nuqeEiDDxktUYQJKKaHxofO2Db4P6Ybl6lyCIpSWx3THk/RZsBCBNjIpMwPKzZjLERx7z8
38YGQxBGGYm8a2Ghbv042jz72xJvdee6EnaLfarwITlrHEgLAYiyW2vZdXOcQgQEmxuZb566BuN4
KCngYBmR9kehZyXbjANyCuFxqjI5b5PauUZP7m9DFaPWdZjzOP22ozOfZbgWGDgU2tqM20aFAqUF
CV9AUWnFu5+ojgBeqUdsnEac+ounQ/cqz+BnGgbSSovOZVyMPpyEK/G+s9ndZls80TK1Is1GF3JU
cUR5O/5j8GgX8Wk9E4c1XI6xgswoYQXHyPCwOpsCg63e0kJOIvWWX27zp4zc8eWXLQViSYRTGfWN
BXiMg+Kxbdz7MPNtWDLd+G1OfS46M4wVOHnFPeTK37oor/MlybSZac3hMH4aaanuJeoih5SSPyDX
qvTwXhsKwwJY2IpCmj2TkrjqzGSWDkptdjCu3Te2/guV1dQaxrQp5MsS2nk8kxorOMjJd9AMJBPo
PKVryx3yWKSr/9a4DP/f8CJk7wLxgmvyPK7IQe0EoeWe7ZS6OrEo/BU+6lZah5e/wf+fnWLEId17
FNirKq6hpregGZAlq2nkqvm8fRWbCbJvIHwBm4UkR/ooi+wZeJU9IjAY3++ng2t1AZybdfJJJO5v
K6vzRzqWX9OxV18m6+90sgSZBb4o5t6Png5V5kN5dlQhcffMBx4RFO9nUyBWId6WsyyS8kUpfyJ2
sIfkLeR84Fmd6jIPUB7Rp0FbRclIM977lmHS5MexEsKIBsDy1aIzKsOaiKi/fJAfLtDsf3tOsaTo
m/FXFlyZ9ta9P4tFZCtob8RDyt3iK7zr00ZEppTQZWmB73BAbaexcq/NXJPOi1pSqR0nw1WUCGjO
QpRrvwTTp0Kvtdp6qV601jvb/ZNnkciIzfREQ3EkTQyfgQ3iRoo8oJQngJYslvJwvz3GqtrSQLST
qb0kXjKdarCYlgvUUf8KadlnW2dawhQA0N1apmDPW8RKpHtgddSEL+h5CyYiDJOQbmabgy8aTlv/
CWg84NFEkPHGwSnRDw9KvN0N5jgkTtSrM5q9QHSXaKEiC6wcGSYhx4CRSzdhTKdOLP2eCi5fwRck
+p3Rx4LEjyzQRa2OJul1VCIyFCy4DHxxSnTjH4AtDgn/rn302JEtrAGGXe8QwPjeWncwhBCFtHqw
0VFpufOFzUpAL1CUJ1FmpmLgDdo/u1M95gCPIliIMheLTs79T6P5vHGOTpE611tDqkxFJWWLQgGl
LwaOWOS2AhygUGKeKomHeMhMXpoqh1pmgRD/8kGfKmMi4EQsolQvSEGCaBtCWp6dclfqkVd51+TD
yCsR+P43xk/QH5Hxgq6hi2MUWbvPae6zA8ByF8t1BOmhCjDBcjbHJfvyTKrb32k6ysiRM0Sr70FM
NpMqkt5gpztCsGOHDeBo6cqEzN5nlcFjKb01G1gSLvAKvszIW18fKLvpcciN+g+YoYfBuNos17DY
1Od2qoIGCTiE1QMO55XewmnCI6BmBw7EPufNiB3DJ+GZE8Q2LpakYrG1+zrJKMFoR3aQcQhH2pka
DLzpNUFA5BPyxIcDzPXY86TJ3dyrTW/fMuvbAAQjI7ZjfsDnsoaVNRnV0LpDw5UCtYReV/svbcUy
Mxa8a1+xmslW4AEKYpBKKuy2JQGTH94yfEvobyPjlPkNugZQUytEiTLzKYFqUZzCPl85GXbxxyj1
nKEVY7vS7uaGgP8aNgQH0Ta7qnpkZ902ao9JY64DY+PqgmKHs3kiKoB3OBC3ODPDdJcC0AxPngb2
UXy4DKfSlKo0Befw4JStYejrxmqItI6iuTEvw09H4ssBwmrsB+war8Op68lzFS8LrA9AAXCWhBpE
oiRR44ED/6MCdzxFiyXPItcvsuQR17pGt7qMOtr2OLtNpTAgQXCK8emspmyFehiM/fPWRCMQ5Gvs
GZAy5/2o0WJ7b1bdBrLLTn8M/p2/9pqdEqDFjL508e+/IXkQuWeGSw1dRc7/0f1QKFalOm+kzYap
rlMMZqPPgkE6HsiaYxu4H5THbCRoIzbsa5HHziRPJd+gt4026yv5UW/sGIrzuCkrKF7WhDZ8XP1B
7J/CI4BWPsGVAa2Gv3aneVDyA1isk2UUjByabwqahf/G3+BOpQ9c7JRMWGqWhYFIsigL1LrMKVkH
qkq5g8GKmHktQlC1Phx9aWmaPPvXK3IYHVCnKn1V81mu0TAkjQFqns+k+8ePZ69nBO9439ghoHu9
9F0KMA7x3GdtKHdjuOhlAVm4WOLlF+tvBhpkrjIPPxpbOC+2LD9OKAt7+F645RTvbZRX44e18BTC
2dGe5IJz7ffXszk9h2hrQffioFnkRn2EtMcVFxMgxH2cyQGjOxtD8We4zjnzrfeLtTKQdYi9ul5V
0I0rVAepGUGOaMhmtkE0HQlDomhqD6aVpDTNz+zU+cRAFff3sau8O1pRswlxVSiamQR4ucCkNfYi
1W8EsN7Gt/tTxkdiDHorjB5G/rQNX4B6aS7p7DYCgLwXpOjWvvPyWsjrbqWlO2UxQmfxRmpfDmLx
y+NjbNY6+3PYpV+PKZPTAKZ+X7T/pR1y/KAvY5UVNgvO/QAXopMJDo05CRGzwDoFBd35ht06/bxJ
F6vFWkCIis5kQ9159fadbxGXvhH7xGNtVTL7ztnyciV4Z4xRBf/Ak+jIRNmj3i4qyCxrPd1zzUT7
aBu5Nokixl2yE+6F/8OdmorF4Fh4gieVEZKfQNebEdL4+ma5qvTeDeHmQItXf4mHtB3oYDWXHfcp
CFjHBCQkhFtCdoJ/Rug1y82o2b9lsor9WnNgqjUbswQwayT/O8PCeHT2QaPtm+Oy1UdV+b8GGGt9
H8+RpOtakui3P/E0FbzZiR2V9twQTWkwO56oOBApRd91ldrNPN9/rrUOdOmzjYRWElPxaKAF9oot
fCI2n2cZ7Zq3/a1hoCFnGiADuo22NxfkI1Mx3KNYh+XNRSGctmpVIujLFDtrg2qGehBbISdziwlW
Astjk9TnGaCAarze4FmvA/9qBp62MXWxELc1DaHsOFLQvYF+mIbt9tD2BhCAwz9dpgv13NR74sR3
/bd7xcS823NHV0rHnWvmzWlxaAsDaXImD6B1JYdOYcPbTy/S4VprdQy5x6+7Qt2TnVzVtWR4Yc9i
bgg7TbOhYWIqemR+VasXsRE5YY7/V+lLwJ6aEa9l0VKt7BSRBbPLwFMtodZxPhkv7hoog0RmdzTo
9tLxkIPmpWpF2wZYzB9VMmjvDBZ38JzWtUem2jLXAiQRM5CwLtXK21vcoGsF6fbRuuaZ7iA3jMJ2
qacqHdYdwtEwUm39nlvnfV+rqNLRY9Z9O2vWAsqSnoMBJZa2jp1/XxOoORR6vmT13L5gqlTLE67B
o4cCqyMkXuEMzOuNvBaAMdFKfJ3z781Jk1kYHnMkgEU3qU3FrfziuqDSBJfTBBeeH88deMrDKfhW
TDPLQRG7LxGjJeytSPEdzdPWNfpfwtypNRQUf1en8MEtBdBBLLw2enjJ7JQHWJPfcnFVeN7up0Xy
3FpoacxZYOeBTuH2PtSYZ0H+sXg0+b32raM3A/e8sEiDU2wOhTbxU4jEUZ98tcd+DIbioU7O+pvG
uFWrIEsbl0vkISSGtfG7yBNVF6NhVFoBGwLkw3+Qyb5l01LPPDLoxmnrpKqb7yT+1BdJ9ceWVea/
aI1AL/40MHPaPLB3tWnhtOPdDwFJyKZ2iejfjZS9/rScGIxvUdWKV08NfV079ipp6+4elisTPF0F
ye7Ade4x4RcPPYMhw5rsbdS6aVmpLNk8whw1dmc6iFAlShE8c6TM6llLutUfSwx1KJCbRJ6QG8nu
ukz3oBcEpMKYpbLHZKq9C/1NLkEuASapkFQSv6+9359v0ZbzUSFTsNpFur4bbwdmXwHRjLBoFGdu
bq2AYWzsqfzy//hdkOXodZJZ1Cik6rzZCv+GxH5OzAR+JoaZYPQ/8h5WiRWS3dXRK1UrOPHfOa06
6oO+fNycdqAK35RSVWtES3OFdvTwcsB1n76IXXWDEwaC5J4Qc3LqRVROpe2j4weFXG4V6GYPShfT
K92s1+Qbd7He2oMYTJAHn53h7W6augUzznRYi8E7qZu+o3rNusyjc2b0XjB+Mgjwnd8jPosHWo0w
jg76DUkhLxxwiBip1kajQxDAE4lg7vWPTuyefPGAfzPw8iDsgEsFYjK3yEb2g88IDmFhU1gaab9w
GR/XBd6MNJEQmFh+UT2lJWW6PxM1pFd0O6fAKh52EIFYHl7WnASvXUmpopyvVMAinsy/sKgLrCXQ
5BYW0d/Xn3l1JF8XPHkEtiQyPRrVWoJpCUfQfN190JTgHucEvsST6DwOM32s0Rh8qXTXpcwdRxNf
Dp9gTZMxiCIdivCQx2kKlkuw+1Mgc70Yro1CacekCBCbNOS0OB171Agxx5ztEmeogCZGj3jJNeU3
jhnxAr0z5mil2eQZqjDWNYBIibHs2Oxsd2LQh3yDOz0CtaF0jNkgQpRL+LmOj9GxmaZpbs037wAd
Mp2gu4te98p05R9KJVHVRbg/Kl4VBRARWFFs200AKp2/BcmaBVpNG/URLxr/d5FvstNaRyafzb8u
MucOCvi7GIEQpaKH2HfmyI1+QCC0vh8mR8lpWRJOOjn2hcNpFE/kdiDTfh+GzYpXVKhFEEu1bcNi
//oi+wJW+kf5Afw5Zh2z6YqJFklmKEK8P4c4kaKBYbh9RmXbbwJAnbavIhyj7nSFxrBSG5SepBAN
CWTizCva6KzDqBIS9bH3xof5MlAf0gAvWUmmiGZmYP/u38Ar1k5ZdupWjo8YG4bFWvClaSCnyGBS
mm5XD42PmU7thdEJeH0Rgec10ytmuKClqLHZZkrqZhEnv0YUQKH9K8QwR7GdLIQobW25Lxqkpja5
Mr3Xz7uvvIug6IbSArQNhoWj7AGpfcQMOgCR5GGSjCCX1z4JKXVnytUVKTzYOXzq2+sCpyLuLuxn
hUvWeYXWSIf5srUZVj4osFtB/W5r4U1WFvQRHyoxoq8doPoVqqn89SSD0ekH5MQvEJ0usfqShNKY
6WHTqi3xDB2BbwhnBbaWz/kQ8/C+a+4rJsihXtVbaYcR3pnUpYK7KPJQb5e0K/PK/Jhvb9ETtP+f
d2XNPAKM8H6yUN4ucRM4Inpa2zkp4Px4qkwTlqdiR/yez6MviZ+1eDasAHbBWTgOQxRsg0sJ7I+D
YBbYkQb+S6L+5JMrXhu5gHKpZZMJJr7z4canBUwRP/ANtlO+6qFmEt5vPpOH3mV242lJfRnJXfe8
L15Swa4WZ6TtmNQ6GSTxYn5b4Rhmh+w6ZkV7F9qjN5925kHhwHThf9GBS+JJF6CgsyZrHWihWHUh
kOJpUApjBOryKoGt/vyXJgznml+zxclYlcM++P1dlzOv9tkZkCJPxdx5PABV4P5/CEC6qGZ0gZkO
sYb3eq5dlXnPpk+fRrr0QYXclxG/rr/907DNSf809SqLAEQ55MMbl+6EfDbH2QXDYmyRd4Be6dY/
hTNpsIwZJuYlfLwNFrVuy7wprW65TBzgEfTDERZ5Sasd3o/+vjZtNiAjTdBrf0VWAN7LWsfPVQ2e
pj9lt9xgvh50xp3sjfZ/8phKkto+2SXH9/iQLRL8cKcZ2XXgtoDXlG794AiB12CMMDvntoQaU/YQ
2MKHQCwIhXGW7m0/6HkAiEwcuiGN1S/kj6b6G4Kw6rc19yjxoQwbDsowrZJqSdrWk/yw8kV8VHbH
ynJDEooE10g7vfNoWxnoeabD2lDOMkAT2w+hGozhVxzpV9QxMp5gc3OW5B/qxgHpW/4nRM/W1D01
JYo06Y94QNAfIGzT71TA5+gnHVutT3RFPPIrqUzk+9S6p7e0ggyy2Df5DO8wm2TY4aGF9My2WLpK
z3lhiQ/RxYlKs7ilpugSRooP9/zGl0TE+4k/ziGxJKyYzmdWLekn5jZoOHr73g0DO6zfeE4dgekK
CmhbSCShhs2+zxlxlZIPzk8of3ht+Qnf19NtACQaJaojMiU/3ntncIWnnm677iBa6K0iDPlHP1oj
7p/YfX1mWk6x2pnDVPmaLoYXuHKqcXnURqLFI0kIRg1U6sZcMEYaYDx8+LVWwo2yZ44KDNq4FadJ
j5laXN+uypghoq14kzNH6kX6HnHYM+bBd+r7TrzU8rme8bfGliIHDOITMl9JunAYJDhL5QHPhVVM
FAFS1K3t5yHGKuf7RlAszket3+ZQZn8NmOcPFWfT4FKbzW3+TBuu7qUh8Hkn7/1bV99qfJnRkNrv
PA1QdfDJPBZIKCL2Hcr6KbxhBMbDUbImoYVAtzK0ip9Tpa1fAQ37y8v16sI59Oh2rp0g+faSFEgO
JPUz+sP+zanljP9LcieGNTQjpjRhlMwm3KqPw/cXQTMxRxfpvB3PdNPUWb4OOhNn7ez1JWn8jnba
QST1dENal1Ci74b1QAnxYV1rZaVSjSEvo8GLLGT+V9TYAW+2jToJUKQM4prp0OUDE3Iv2BpBXr3A
ZA7P0OBTpvCT0h2utUpovsEEliU2RPb3nKkkMZs6Lzj3epLBYksPzzqo4oX8jCnlQxPi4TZkJRbe
Shb4jG9DqLRXPVKkGLXrWoMhN6OhPcf6kuEBzFu5T704+25RoovHHUbtKGLPOz7Gz/WK/dOHkVJM
YFmlYY1V2vZP3raQ79IUljQN/nBe+gcM+PMj70Ki9dhPe6yHxFUXmF94lVSeC8iUORRE0AY2ym1G
khOFhmubi3cw6sakTQNqepEwz+jtSYHRVhytaM+L22uUFMOfXcfc2+bzCW97DD+UGpJ/vgqEcxHv
DkBdu3QRMNgZm3QP9iGWXK31lPlC4VRToBkpw0r/DvGAOTS0i3SZOfiknpmj4Q3vs3NuhrogVhph
Vjz//VDKrV83SYpxBnlXx2ryHpEMDPSAbnOIYJHTNW4qLUIj8EyDPBd3qrw3KYzcJEb3Lj8DR16i
amM4MhHMl8UQMxWtF9nGRfWBN9Knb0AFV+t0F4rmZ5o1QojExD+2iwGsKumHYr2qeNtzKyQT8OKF
9MqVy3ro/NUDkOfy0hTb65paToXAkJLAr9yKsHaIN2bGb8D83uPsZPz4B11WInOBc5lhpPxJBd11
3nFSCG+rK1EXRYr4u1TpIsGjLUoknriwoYuS9LnmISA4ClEYwljIXst/xugri7uNKguUE0P7g0VB
fmHBA8ngaBUS+m+wocGB+uyjfgo7xw8bGYeyVpuqRWpuygwnGOF8JDBvQQQDfpVvUG7Seus+iHbk
WGOTQ9aLoAGa9hkSNSh3u8OBJTkxB/DvJ/7b/5fs/66e7wD2qk8AlMfETxJxHI75hCcX6KhxqM3x
EULK4EkX1VgnI8P16hYGvIBm0wCH4OU/dIdu/DxmMEo4X7CApFSimcuVaKqDCInhHchL7Ur5bfLC
V9ABYMZWuBHVUYIv9YlGpwVW2sRdxTwZ6zD3z27PQOtrAOmf8rHDgESUpaRxUyOF7VfJdn3Kxqa7
cuGT7f2Qs9VtnMqZJRW+96mbSnnUiM/sCTB5GwZGYniyD/JdpmsDhnv/AYD/cYmwIGrE9w8n02/V
BlH0+IaLQBfDNUcQUpBwv2l0woTwzpXR6VVT8GYa/AAH15IJrzerzX/CsWiS9K2JEImsRCYnhL37
UqlnSia15Wf7/Hc45/jWrpJItdk2r+OtNuIecLRjEx45ZM+0ctuzEm2pU5tbYBfAq4kNewMbLHRy
FNzi9CLA/34d+0khhWbFLr4ChCQ/dTfLPiJJm+fCrcEz8fs0ni2pzIP14SCQD/oVdyghRw42RgG9
E9dAgwQMqar9K6FqkGarunUbOUbe2pf4JNbsn1XHyjuUzVlpeTjC/q0K9Edmii1o0SPMZgbLlO2R
gl1j82n6oeYP28kW98n0/CjVPZkS4GA3tSxFepBjjuBDqd6MV+Iu4Lmtn3spH0aI7w070NPrfO0P
Elz4U+X4CUA3FtjBtkE4bDFvKvbLBHyQ1JC0xfos5qgkTUjlBihGNEw+ov22JyAOl5Rbp32gyVD2
SPzTcb2Nnnaz33Cv9B8sy0q1JjU6Ti2q9SNtROXax2tEnFi133MK0To/jIzyDBxO4xrv1Y7ZMFyh
kOW+xzOrWLdhCY3u7gFvH6dgabp+j+5BjmUqFcmQ6RZeoUN8k/wRQawPYdKHM8LXUBriLvNhMWq2
fDiONte9gqDP0qUJlBy17Faanw06x/Ekhw5S8rJ39y5zkOqyA7VowWKBHaV52MBA5U9v/R1hzqkP
3gf0hVzIVOz99FujwPto3ZLrdoU7Im7kOk/ZOamW+QH99Fti6HrOkN3ySR+XsHdLvFBIXL+k8ybN
Bm3K1kA0+O9UvW8xuR7+s2a9oQodj3GVMj2Yt781ZEXdrUntYaurcU2mov3Ta/R+14azYy2r9Nq9
ReAyGVHnC7oTZr27LBxMQpEtKlue0GgGmD91yUhBL5XBL5oHz6iPrHhENlOAvI6tIaDWyENf0si9
Zi00T2iBbgK1Pa7Z/6uCSm+2o4MFBYNeFr0DZBWCovRpm15TcSP6vNcGz3om93jaSrHbcvARTTdX
DjiYLPrH88kSBhHoUuIlgVIFnI/7V8KuGNlO2JuPDmW0foIYiUbFMF7G0WpnTcXVy747g+iMsW/I
lLh4rOuy3Hp1qIBT1sWgT6oIcWcVT7gk3s6vyB1cF6gHmS1/6Y5a5NXGkx01p17XBuacfnDfl0Gg
GFGoRjzNy2pZHygFWr4XwHGBoNfJgSCd1MA4smPIkXD76kIPF5/3Fk10WFRHh3fu4Y0EbmE/o0Ef
A8zbdU3fe71JOOLu8rNBTCIfAFiIlgSKEQDquX5WLoMrgwkNAUPk/wvvijNt6l1yMvLR80jQsI6B
xBfT7qxJr8D2oKFoj2xyj+9Mmsz5DbhpEry4a3TzEkhpLXM2NP9VPmimX+fIusU5a/il+sSA8+nD
+LpcwjnHEKZfBau3pW1xmifQ9g4kWmw5MVBpsZq4+05v7KTeRTHdvNAxRf27F6YbnnItjjLtVvlh
YSUvmnID6ectDMFKArsfUOgNBxozkxH6MdCOaPhbEoowBYHM3Bgn5DyZgfoReACfylpmTTUooJRP
s/Yha4xd6YHFDYDWnVgdUExiIKGDj8Wb2Gc6F9Ekjb19BfcufuQmu/UMbDsAlOSdhZYkTVlhiK2g
jJjmygTa1tUqRtnLEpg4Ev5QFFmq9l7CxJU7b4yCVeDqvaZ0hp7dUKZaQHiQQJAxjV6XYWmdfDWI
Pm12NOaGuUaXM0HSI5iYTG7jDSidjDEtmuBrnrUSXWSy/OP5BAgObF3Axk5vwOdC1T1MrYfYB3Dp
VabpLbybSC0tuJcb0Py5ws+fafcdB3AqrBUob2rYf1ZC4Zjvx+610w+9DNIkexKhb1/q9a0h0GpF
ylouk9qXgo1eJUZZKrt70ZIfS0DWkyrElhZpCLZ2OsZ7AJA8ftNdZ7ruRgYS83SZE2/7r7Aq41Ei
0QgIoVn81sBzAGDoLXlGG0ozKjtPuWQZU9CEmzZTXl+WiZ48B+vm7QR9m69jgla3rxmhbaupzTSD
Zb/s6K1PuwFgyZrQGsZM6gM3aLmybnG45p+F59Cz02QTbhFqCZco5uKpbya9F/FityGuoidMDVJo
wbiryYdEKVAbtzsDujwDmvGlTZuS+IHBsqORs8UolZ5NxrbVatJ6DCAcT3/fiSJe/lEo+xVDHJM9
A4gLCkojtIV0IWtIicgotaCKOaLvifXpSs8jiEoMOd94U1T1qf/DBYZxiiPlzPvx8z+qdckndHp7
BeRhwfYJehqzDgaSbIexSNkoqVV3raJm9zN/nSbYtwzTtYkGTwUmfl7Hmp35y/wkk0tYZHqJgpFK
Gjo6LvF5GxGPRdosyYfupSlKJ4mjwH/sr+mgFCOw9VDdenjaVIHFnpMAgVtlzI3Volg22e7W7Oom
aaSd2hmjNl5GE+TQODgMLXJ1GycuyyT7sQVTj1ScgM+JhxxS+1rHuhXoow1Q5gn+g6DmgZlfeG1w
28NA4P7ujOqU5ha+4mgNji3qVnPjAVMOCJutzDyGz62k+gdJeAqzAeeyiMe53LoAjPvDIL7GnzRF
R3HgIGzjvWnOrfGoa+yAVyQlsXg5HlqmLAXZ++o9Q7L5SYwaVvMGuDcTII5UMhEuchtxlAoN0ic1
CfaiiN5Y5uSeGGT9I3kcr1nc2KTcp3jPBnlqcv8jxUvqqxH8ok3eG0NJoOOG+FWev9KAovpeMU4S
DL2G1CX8UvAqGa5vlPdMX+1+yRQmHMASU8QDGB33bD17iXd0yo9hJ9LIni5cknJp89fzri1AyqDi
D9rle5eB/4yz6Dceqn8KTIU7OWPa3Hc3co8sjMulf9J8qpOF/rqwoHl0gJeB87Ro1S0/vGCL9C/o
Dx+lYjbxHDujWEbkjUVI0xBTI668wHJF9oYJwS15kYxDjTGVCkQv/vejvR+VHgmKkoZPsFym2JZ0
vlaLBYL2KgSPgxl6My+OBWJJO0y30eb+BvuhYNy9DelaIgNHr4FOzoiZ+zxyN2tcduMiaJJk/P6D
wrui1E2MVexy5vmmIyBHSVksA8PndZ0xKrl4Gspp5pqqvRDTF9/ip2L3EiiCzUh8VVRuV4rcGhRn
EPfsnZcqrm0xbIDDIYKEusYefevJVpNuR88D/mic7itXta1b0wSt85B/ZwlNnSHc3tk9XveZ0Xec
2pboC/rLmlcevIumkvK2EHBRWDWE22DFSwbDwZNoZ6ln89zGPpnkVIemPLLp8lkT/EwkH1ObaqkD
f4sO90mE3s0oflRw3iVzoc19JKP8TGFuYX+uMZFKt5sB0sztk0OwGZ3gQQfAkuc40LlQq16Cy3zg
DanVcmaZuoOWcrZNXkSWpFS5MgXh4vSqiwLOtnGEG2K6OlkUqPs64iOKsaF7r5xXsXbnUVzdC1JS
M3baNIizYCcsRYiXLjlvNB9sQyoVNDuc7wR7yjyLdtSl2q7EvNbvi9nuqhWwbn/F7aetFdz3Shoh
NULKqmP8iN0YG1PCy9tcGwnfdzS32+T5MfbOYexfgDjX0b9NQJYimsZuAkoQp3A5JHqtn7XHl9va
oxB+4Hq+toyKb2IvfhiY1GyRiAKKjEWgVr2dPQ0uwO0QkjZMhzLgcCe2SiahCN2BxQjL7Isg6nZ5
lWiV7zvg7nznUgRpabJfdcjZOkTORCyiMG7KBY4LTd87Y3vagEcGw/Z2krK1gGNA7TPrprBMgwTv
/PpqnXQe6m/kygyZc2DgfBSOaUuGF8hCTs6lCLWlxkPJKs5aMod2MaPbKxA+vqtvFw72ENLVtDt/
UrxWxQh3RTGq4sGeaq/P54zmOaFEtWbhEIbnR/0nobw/VUBHabucrDjnTh5Di6hCA0Mfc0TDpM28
dqkWBb5B/AdArM4n/VWANb39+A4pUrZmoq0IKuwYpZMhBt1pj1uUzxRifKvU0y0HMWfIb4xA34rt
7mzrAM8GAVeXI1ZU7nVzcVnMZ8tK7kaq38Ul0M0c59zs6SQD7lWWcOIkX09NNa8HhqRAPleWCsVM
/a4syPjYyNvg7MmvzjXra+aRkn2E0S10Q+5laa2eOyAKjSjCjnN/s65TNM4CfIvW+j8pJatoxsxf
BpG/Lc6RkvnD4Abhurot08IQ+9gVxHaX24HG+LQdV447dFPEJN0yy3hB0DNeAwofJ2/mGazxvZuq
bomcAzR1QlN/FVYJUlOAKFLoURCPn2pfn29xkl88SplOcmOw5bAY/UVcXAt8TUR3NUYq6H8H2+0T
qjzSJb9P8V8/RGKboowu4oG4zNdX0PKZBXVganNH74ZzPBwnSlK9IGYUgMIHh79DeQwlMITZPbvb
VgJuUZfYgmJTglRWZkN8j/WsSMSJkgIZ9tOPGcMGk81quj3iFaaOPzNmNKwl0ph24d6CqQaakLXk
4hcElyl3Tzx/RRCXL80x4e2cAmnqnJHrgM3XK6y9RmoD6B2f6YTWGSm0Ov1mPspunvIP4xScemqi
Spn3V7B5Tee6mYovLMoUERJ2ZRIQGyHxyh5tEmMEExhgviRH2/XOjeKRfgP+43HBTkoTStQqF13v
GlLy9t67iidFI1VpYZYbHdV6048n88uKfDvsOa2jpksZx5ALBAcPV7TVdS0fsaEdvQ8eLAPBAHOH
LFj7XwgYxAyDf0Ml5HvtS8M4qarEsMG4fcPJGyadGWMCoHUAQEzAx6pwwqHR1h9sCvs7QRef/It1
C0eloM4X9Q2lUIC31JrUGG8B41HyglJAElp2grddv0+oEd4eil5DHvFurFM92aVTCffbnysPEUu8
opjw2RZBYi2Ey5RAskM0I/2hwxDAH+eswK55kBBENvNyXqR/vxyhEHhSfjbehDUXWfNG5bfPJ5zL
Zk7RO1c2VcQXwA00dE+6E5PbfQkPQruxTc4IVRyq1UUM8E4lPZaw083lSQYDNQJVuWrVe+GwXXtX
oxL+eixMjv7E5czI/TvpulSbmXLpE5s7zmxDxqyWW25Fa875QEFGcfFgdZ6uo3BEcjJ5QoUjXkxF
Qy89LSj6G1es96aqj0Ys0Yfqce2pq1xTBTXT7cuY9yYxcVzw3dEl3jdxEOlbwJqJBBWLu9ZJPiug
KDkroQYOQOFPMOTrISgi4ZXVWQvPz5GHWvtamsJ7LkRwEazGFKEOzNDdMqxd+lVrPI8ovsMI8SO/
9l3vzBWnWpsXKPnmZylQi+vrak72f0fRgIIxZ8Pf2eEpsU97KQX0zJqu+0bCv+kJQIo/99V5aBpU
FQmZYWszOUSIrYofXMeArEMc7JghE1KKQuDWLc3+x5guNodRirqVoeUJnnUPduKNKNbJAkQaGq01
pqg0cIj/QqOGooGoq01+jam04s2uor60ZxVo2Wc64hfWayPKhADtQqzkyBeTbJKvqjJXZXJtAeiS
c+DYgLY0pdI/5/BTVjzaiKYNyyPk7cm1Sp8Se0p5DxijJJdfB7UFbOY67UlvvwTm1Mxhi5awSES6
/LvnuUQalGSuR6la9d0S7MOS3FqlshpBzHTSSyfne3tm6ZYNuji2PSmt+GEOkrhMmQUGOtps3D0O
iNM4wt72DmsQwJA54mjlnN3eJhdnGmwNgyR2KoX+UhadgOA7wpgx8kSNRFeeI8waqbu9H9YOq7ld
uXSXsS9kqfErzdZi92V++c3a6aYpHSvHHaGR/Nkywx39n3P2nS2JpRT2aT2UYU/9pDSKeFokhD81
BHbFFSruagG3GdTNpbdNfBv/NDh3vKXm0Q9CWSf0YKBcYeVBLggJMSAJEwvdaxhgwI+05WH67n4J
SQIKij5oC4v+6AmX7KdR74bK5vi27HdKrDB/BfuQN+3fMT5wllXdc7H4zSvB/1HRXE1b4JpUPa76
IFSl3npI+fNBqJo8wp30bOFDx+1Aww2uXpeT4PPqFe0DkDvTL1qWI78N0ttezZXF4gpAHyFr74hw
g0ZW5mbjLSPvectWUFV2VD0ZWbm/iDWlLp2I5SyFttr95qPs5Yd6W82aWkXnZjcEC8CSdnp7vNlv
TW+AWpwi2BV49/Aqr5FUJoq1QeVEPXikB+GvuB137fMhhDf2rYhO+fubzMf5yHSGHHL5zpZhROCV
k5nDY9jtEjJA+NU9gFDmywbSMvcJMzpc5ZGXK/HNCGgUZjftw3DlaIqnQA40v+kM5odzCILKIT1H
mvmBtmAjSsaCNv/SrejcPdCRHMH5WAB5OVUHRNiowTh1mENL5e2IUm1pfvVT8smBr8R+wCgkOi0A
+F6HM9R0N8pcCYH7tpLUjKjaEhSU1+sixCFtY3PZ6obZBPyEG3heAbvDmh0AcxqXQn/n9+dElUsZ
0hJczoWE7hkME7AUTRqFcJdE5TQVo72AnXDcttQ4TMLEdMrXsgpRSzANNZm7KeTzmy3WtY2Eclhj
a+hBbPHYIhL3hrdF/qLwBEo7Gk9vZu4dE4sifFF8O/jCw3CuUHkGmtv664Fd/IF1nra/9vhESv6r
6hlHujgCgh2DYZ3mhGLbWjtg3NJe2pJSVZgUWjaz8Yv5CFWxhTn1TvFoRbgyxsshf87hD1zMgGyh
ZKSP5SdfK46EfH9hwyxIp338G0N76AIJdPzBp44fD/wbVSDvxR+0+rm7VBSKRXECHDYmDrkEUmPn
DyHjtieYXXROtsgTfmJ8TCCF0vd7Oe3hX1NOZuWSoxDtaUuUK7w3thtGU7f/+o5+N0o3DAV+GwTU
64CKW6d8WJVu02a8Oa0Bw/v80NEH5vcGYqjXVnOx+gSwAlgbeY2XCjujOx02/ZVqjLoNcuu5z0ux
6uanAVWINFJljTCX9hdYsfZphIxNOWnYqiwqlz48qJ66XxTpUEMVT1FIQORBhvIQUPD3uqFwgz6l
2XyUF+cy33c3a/x+hhBHL14POsCOHbeyaVwlzFJAoIlmVrbH5Jjw91F2DmLp0AHZW1NbHv686MUn
Tu2Gr2Dl/QJzrYGnKAC8KC4uHS5Pemv9sSOC752LEoaixbMoDQkg6n/p1Cw4tb+58M4zd0NcIUtb
zPGHV6/4ngBjz9AKLaIxtTPf4/1vPHZZsS+z/8OMbcKFXHFU/ueX5igeioYjOTH1CIGwxyGpxjcg
KJsOSQTJY3RqsBJ87nmRwR6cegL3hngMGH3gsjYsfRdbAfT/NeMmAkbc7KDR1Il0ASa8sihqOd/M
OXDKAiwUJqaFLGTwfZInPxLZQoWavKkZ967kGANvVMWdiSSppxSCs5tS/g0O3phuGQ1EMmWwsMEE
gca1uz/W9N8MndY5QI9NQGqBIxErUF4TduB+4DSXpTasDWVbn+aExW0QYQnOI/1zCszQw0iRUYLu
7p5+msutlShtjCvyKGsI5RL06iACKIXKRmO4x7JqOqQHlvPX9vwlvP0scJki3fflG9i+fnUXtbOO
fGrjDUvR8nPb63K/TK12T+DZAYBs0KZ6d7ba7hGWEgsk5OGlbbNmr0SBGTkDjTVfpS0anwdFKs7g
QFs/E9Ov9j3Ny8fkHxHpbii1X+ohQN7xzAP0gu2rTCYLXBe/KRxy9eUViD3Yjd0WJneZ/1OP6cT6
HcsS/4d85CVNLnh8UtB4C4Yn5JSfnytSJN6zNRADwGvELjqjQAWKWKxHduxt/VRzKxFKeumYA71+
ZPqdTNG/9AtcFsm2IRr0Tx7nG1L3jyTES18ReMAKq7fyhAJXnik+zJ200KPrFL2PrbUnM5arQYHz
AcWg/7eEi6KtzYxiFws9cmCbDyDqUXy+TMqdO/TEWCoBs3Cc7ruPrrznKNn4hYEeFmNgxYEMlyWN
WXwIPP23tQOrtGxQgwy4HtUe/lUfig0tyeGcSP2itCU500/Yu9W7A6RG03vhV5pppSdZ3TeWaBR4
EUk+lFH8mOsH6yArj+mvS4Ul8UJMGtSVk9lKw7Hnjxr/rffB+EhFWdHmwDAsHltV/v0958IU5cWi
/MFPNy7ayRJ+FOEz+9RW6pvQbaXzmV9a21wztGSkuBiObeu4MPH9btoR55wzN/N0xlVoxL5vrs3T
oIpWGKwZgRsGgfK0XXPLOroeCQ9VRtztiA419A//iT9BY49cDL82IbSD1yP3UEj/Onl7FPO2M9dV
hvZNWtvnkviZ/rTsrcAhfaiRztqtC51rcMYH3cj9c9g9ljywnzrcCBCzOISL+v0ALl18CbMjRaDA
5hMqPwLJfOej1iJmEuPrNcr74jTABiCyNCLc81gsBi/h17o5kof/JLP+3sj+4+ZbfTadlt275/xb
R2Gu72bgHZowcW257/7+iarPFtb7dcKAiC0gdwWY8i06h5X+kByknUYL2ye3lRwFC+YF4dTIsfUV
VJVUeugne0D8WPqN8cw8ztvYk90QwD0oo8xtJ24KyajLVgU3kNleICM2VL/Ap/5d5CRaxl72IVK3
wPqlkor4qE+SupLN1W11vYpwlPfjukMg95pX7RB2scVzu+FTOw0BK/KEfFre2OFTnvAxnHWA+ko8
/6/JiiqXJQhxC2vqCLWiGCbReJDz42j4zDMOMZxJBrfTwwLHj+zXr4Pkk9Kc6D7iGotctDG2qRHu
iGSDa4vbvRRAhBQZsVR9F9MtHt/7PlDsfwu7Af+2e2UQknXvXYTJ+yHONk4qqGkoPiL7Wy4Kjzcj
wAPKIV4BnY8J/Y+ROvPvCXLnyENS7dOiXRT38HfubPPNbmHpbjTsijhK8ClYFbGKXIRyPkvbW0be
j9qfUH5Oc3qJ/p7yXGshEDfBh790WeYYv/k4KS5mxSmwPq1myjwVO0T1S1/mq+9bonOBmM8BU3Lx
Fh8e5QoeHyb4LZ0x7Y+iJh5Yy0DMn6ak+OJ4MTwPiEBLJsXnltSq67yPJM1IpaWGhEUGKTTiU+hI
fZIHwOT1+bIHmPjVDrs+fpe4jaXByxn9UbpwCKCfxBtP/tUDmpzLHSkZexhyrPdc2hYqXWdsFPSR
LhOAYgT6vsO0Y0DL7u28FnIBnqlPKlcsPuKyd1UndiyePPyzlsQZ1jVptvNe6++bRhXNoOoijmS9
LR5J4vVQM5Pf9uYG9NBBbSlxXyRVLqLVLyFmTDAsEzyW4+22MQ920I3L/OXr7GRClP3BVtsG+Udl
/Fe9wQcUzHadUXhdUmPqut6YjcLjP6ulpjbVlIjUCvtlFsASFUCOtRMWllNEGWThFU/TYQqWaNwd
CQ1zGnbCBncuG7qZZbIm4ETkwOnaktitPnh7MgEOV1YmYarxWPrFLjhJgczlIjNnmwyz9d/qU4su
uMEfFrmZcBR2mWRiJDieM7z7zx1b5QALVHpPs1U2xSVmGqoupLC1ti+9Y/vyyG/YE7wIJaAQvy4D
VVJc+NJJvufyHEqgA0ZplIn6avnBWyR1gCKC2nPtBgtw89bHjhDoBKmQZZ5NoLvuRURM8UHDwgF0
xRFHS/diXYDdgMrGKVsT0RqEjlCF91C0bLP8duPSX8RZn55U7LZtu9LGHXDsErUHpz17kFZxEhJT
L+vqsB/rK3fRm47twX2SRKgn6ZSHEqhDgujnUW3tGlKPvnX7nLgbNfTab1ySKCdJkf0FPjth532i
DlOnMJvvGclox9ECvf3ISUZBfV17EYew9XFZMRPBJ3Id0bJsdTKjK/0wKedO1t03LzEkYjTwNxJB
3BvPrGOYrM4ApWCOfD+kSBO8S0pSHkPL3wGayX1ggZY3pdKmQG+E7BNhyYFZkYTDGzk5cy39pWii
rQnt+oX7h4R0MLI205hlcXn455Xbs8uddtwYK09/qwcUX0r84Nn32HY5jcRY7Nz3Vxv+AtXksBmW
9s0x54r/FsC0upU9cB/nZ05XupWZ5L1pk5dtJp1fm02oObXYJZjanKD3vZqvzRCUez+xhGmFVVkd
qBdFyfzMiWbQbMdRsU8rowOszDCNKbbEt0/aXOjqSyfRvjIJhx+dzamb+eip5HLdpwgFpRbScC6n
tVcW3LM04cVYZ+asAaRVwSlgQDpoehFyauikogqXdPOlfZSDKG6MkaBCMiome6ZFsBLDEOMCBoqq
d5+KAKO0XjpsSxOnJQHk3+nI55IQiCtPP7ZzN//vAxCFPTZUiXeCLwn85TcnObCW5D8qZEW7CTgu
uLV9Vtuu8OdEXUeLO1uwf/CQwnPl2u0w+d+wYSEu2wKkPzmStLTLz0EYZ/JMGT6yP6fdf+xRMPbb
wEvq/8kDy/kvw+Jlt6lvKJSXLD9ilcb4SDWyATJFpH3WgPwWx9gA1E5GXuzbsb2h67Z08v71T/lj
tWzkfqQh9Zvhm2awzru4MqNUy0peEBkezgfudsWC69IQUwRt5veCVYd/vSnTU+5+Qjd4IawN6XW/
WCD28xY9Bu+x4uD80XMgGprWcbL14VRAN5zawEBicb5XpXrJec1zmMjWcZjlpo4tY3lZ/V9CfX6d
+s1Sv+Zp1En2I83VHyT9zA9hdLAbii9rtQCSn1MFFSYn/YNChgxgrpYvfvtXZ8ksdgBY1x+orNtO
AK6baHTjTJRnav4jCOkiLSXUtGuvVwUYwHiOaMEEyzNC+R41uPn2dSn04wxxAVaBir7TH2A29S0W
41zIZNz0coJ+9N85s5lyui9MG9OviYL0IsntAZOHlYiTUUubsv/+mt9mg8FSHmV3HEqXutkSzYen
iTRBs6EHGYBcOwhHFVAFy343qDBv2PLUR6yePoyLguwrjRu0kX4Z1XFof/lfeiIPUg1tUKS0DExw
2dH2RAB7HqlDpIaj1bsugwfuR20Wiyogbbbmna+cKWkez2PL2fRIqI7ZfFqFm/JJUCIzfzhDTt2o
3pXi3NLUDyYSs/7RUCP62NBoPELu9rDe0OYe3QyxMnPpj1lRvhKUCImFaptsge0Uyeijz7hfYI/T
dNQikDC9CZhQ/5vM+naG02i7VG4HE7PHfz0GmzmEy64UIcOopuyCO6vOBAtaPKhrmoYHJIfzLP6D
oRSCcus9Un/4OReMGebqIYzpuyv8pmS3A21bmUt0VoctQEbboJsUwl7NQUg6fuVR8R5DIa3026Ps
doT27qIkdaRjPiU84/qPNpaQB6kNvLPIafDMngknE7zvh7W/4mjkMKxu6VwPpiQvlSTBC7ClSqpK
cmfZAk+yKxhrGPuWnvqRfq7kEDXxWK9nyG/nnIU9xMZMukcdaaGvMigLaY+2WwYv018TxiWWckqA
iZUx1zzQ6tClO8/EPO+lKO2sdeq/gAYHo9ysfEtmv771SvPt24salE1eERucseGvrCHzTOdvjC5/
gs9ZKDYl4m2k/lhypRxVzMV0KEKnV+YVVGsrS6vKRMH8jdaE9aENl1de+cBnMtHZyAEvLh6ejGjx
HViZfwhqUkMa/dHf1ZGM2f1Q7r9BEyQEo+2d84QxpxHz7iaTxaSk7GqRHEyh1ezk/+VX1//Y0MIo
SdPHkZpsbcGCi0o91XdEe8PZNSWetqTaibaPdZNxdmx6GilefthUmuY45oW09hWa53jDwoCcUx7o
JDkOUN2MYQ81GzvU4Q9MQIHP7QrpVHAxZWg7ZSvExssGuKI2gIjTKrtyk3Z90Ixl+m2TeLxHjhDt
PzpBxfmJyClFVRkiqCBtdKth4l6Qgqdb4PBTap25v6prC7+XxVX3AD9fB2V2wsTZsUGM95YRh3Gt
B8DyVJRRIb9kWQrUNt4SmTLW1AU9u6MWos0/TXfN+maQjoDUINOthTKNzAQoPaIWDtZzH+MFavAP
saNOiM613Q3DzbQLg9wFv9cq23EX9/uONyXaBL6Zk8wqXArD+uwg2jt7IUebfWFVva7Yy4JKmSPf
BzNyWXlpYCmIfxTTi8FlNEOBfExwz9kDjptHW6Lxq7ShTXMVaXUZoqVKaKNkWAccQ7Ee8JqfpiS3
xFw6GM6YPVZFmE2ozhoY8i5jPqNVz5WqGbt7FKm+BgBZ16coE2rHDlmScvhgT/ZInPC+eXrEdfIE
T+VvDcexs8Ywn52BcmUlQisjOHRA6SFBcITJt3Wj/5SIVjziyIj2EzTuOvKkFG2SNbqq6I2jbnxa
BZqNzLyt8sKeiEGhE1gdwge5CdjypH/DuSn2vIIexyfcgvoHNirhaOXNHQrDunJHyUM/VJ3nivux
04hASu34pmceXHBRDO6JSf6mbMw0gck3Ng2ua1lcZ0b7GyAk4URX0KFIpM6U4LemqsZ82iOMt2yr
ZbhdFFyj3b17ZqkwpPo25kZyURuneORTIG/5m21uK4Th/5KtHDpDTQN8TuQRwCF0Z70tjqd/Bu5J
Fi0FI5kcwB5ok4j5STjyrz+1gxnTalQkTA6HM6PVqXS3Vnk01l+/RfeGX7Ge6tjBQsdBZkjX+7SR
RwiDRdklhZlfbJ0bUXdgk8ZKoEDD9g8ktZNLqn09yTCoZ5Kc63P7G6TBSmHg8iAh5irZCXbUPUhp
X7TxGQw1LW+cJ9vBndGkc7plumTenHW1dcI9bmsazQF6DDlbQVdrqlBrieKONa/ZvD7UZcb2qsH8
9Kns1mLedvXbNhaVbX4IBl41SMJLE6oj3ZXsRYhbY1DnpuRIcg25Oda7adF3Q1jRUeA/RkrsXoex
qnI0cEamzAe0kZusNTFXZZqGywsIOy8zogWbVeRLwmCce8tO+oPK8VHDp1kJ7lTShqsnVLFiHVZP
LbIdegYzCttboiVZm5wul6fITIsNW0zU0q+k2vcaKcujLWG1x+eojJ7bohXmHeSr0VTlDh8LQeib
B23Ts74CFdtjic3MjMzKL1WQVHOMo+2Gm/gnZRMAfxxKgm1T/XZjqt75go1wKaa7Q3f6JIUEzxOJ
JSAxq3F+LKb9P20z48Ne+BA/p4dDv7JN73y8dHPyzGYXJXMSteBIaWJaUfY9z7dK/s/krw5T0r/o
aiNmT0ljeAOMlNd25AbpCbihfcS4w1XLhm6qBAFTzs2CvwvCtQeZFNR1Ojxx5MAdYvcFLVV21jkD
nx76MBczrSI674LWFuW1d6dN0CpkpumBWZ6U/YHjtpSvHRndhcsv8cb4E9XlnVH09uWGiOHgtvuV
MZfKhadV222JpPjxg6IPNoH4o9gOzF7iFf/67zL6SNTzdQ+gLISnjWYAnVM9UKzlZbl+kwgTY5ht
WEj/m6EYpFUxWpCyQ0z+R6F/DXP3pTCmTQ4xafUV9zZpYmgDtNI9J54z3zwNcOTWVlQlUosbAfT/
ZSG1jq4fGZ4dDs47XFLYu6+2K+gChwATXtfxVfiSrpFkogYUTFg573fnKAzw1AJ6R2cPpfAMpLwl
D2GkGfZ5bHpx1abvFyGVkXonLsCOb1yV0QRNcJuS1/j+bEir727dXKXLOnCUAYDaxU3zLsPuygL6
jKNLbztrZS3w5gkYsIW/2yq8ZIL/xg2tLboj66KWcpU6yzN8CXod55C7aExDC9jU6cD31vbUWeVG
PGX9DHX2YzbEoHqh2fLXlWVehFEBZrUlXCCAUg7bFyERiYelN7iGFUtffQ1jg03c5v0Gxe61IL9t
rJ+ne9nldnuXKPcVmvx3A6B9caIJntbZE8yTmrc4WNpa292NhBl8K+VATWdPMGYPIXPH/ZPQo7BQ
2QwvWKk+v/neUc5lcbA6FrjWdF6TlB0uUfb/lU20zHDgRgOQuddSwGBBx0xs1Tclu4kE0R2IlpyV
SJPX0zjMAQ8g5CIv0efbGjvTUjo9anCJVaN9mtGMYr9/zM59PpU9FB7CFik37FAJ5S/HnnQYAKnG
dma/UkMbOglBeSGDb7R2YoJ7Y+krfYtG64A/QVymj1DMXaL98x3nQKUbrP/dc5wgC/OEKycFl6eg
pDqq0Rbu5jihBuSuoHjIdvLoyIxisbNj/c+wa3DDNp6Dmovks0mv+mkzH79VZs24iu6WIUfoc+1J
euRaHRx+ZuV1PCmbVwR16g7z8HMap5p06puvDCqniZTKRnFZRDkzszoVebLJ3du3+oO57VeeNixq
ApVQJz77vV4Mw3R3OVj0wxe58jqTkjgI3cD6nlKx/Wx71kMAzQmf7fpTH0/B13k6f7uolqqOWqeE
36HvsWnXZ1BYJEQh2OfIxDgJJmCNrvIM+DOuu7lHhAXSonKsvVac0j48u13qJyE0r8ttZy4Ylkmp
1kHw5ri3t6WB0XhGf0QJhW0r2k2biwJJIVACMndcxQeg3oDjn0KDhLqzDli/vBn8tnUHPdLgtqDz
AUJSwUS0r7YYpuFNtrwYGYEqK2EXdMTV2+ptJUUBIETDiDEc17k+Um6ci0OZQJS6kz7l2KZBWDb4
NQojzuZF5I+cRRR3HbP/ygCULVX56D+olUqspRn0Mge/KkLrgo2Vy0kbjbCIh3W0ZDd6lNeun38p
3S91csV8KppZbaXFVvLaQSuKHkI6sBA4Hq52RVElYPJVWf8eJoPnMlZ2gAXavEFfODNbh6ykvBJF
u+cAbiO7kI0r97nQyVeIZML/YNRhk6TdwgogDH342zOuTjZ/dFLab8ZPJPMIcD/2gqHC3lEyRuMS
aDr25SjCqJWpcENtpFur6OUE7DKvSEZE3G2d+QiOIX+1ht7+jov4Jp2wOecf7bRu6gELMqn/xkWa
CsjzRixXz8KDXaRsgWVRdF7G/gCffqYyb9c+1EQQBOrUMc98mAFVmkNTaJPlaRsHF0nmHn9ogD72
zQPwQtQ8FMh6+ZSTXXZRMKGz2cu+PGWAR5Q2yx2DL4rLEV1qhlU32F2ehSpFTdgc4PO+2ezYnZAv
ban93s5b4Yh9u9zwkW2WjJEh7E7uk88I3nxBqA10/vZGaSI5lRDYxMH13fq2EV7B4MWRmbMWZ31E
5F56nMlGjxV3TvQkv4lU2jou1fu7nAC59E3F1GTqh2OuQ9jo+gxxupsEfw9uoz746z37F9LobsxE
a3nUBrEy7FS+krJovqbw9n9vH1DGwQ7DepS85yfCeHbSG2IDW2VPKrXfbGIrnuUae08Gt38rCn9+
mwgaBw0gLX/7befd6D2r7IDdPgkrsLsO+goiSRUKKcp54C/8E0+G2V0WBgDHyqgAGSqq8czSO9kJ
9YFbvb9Nhj+Gi2XoTm/xjimNRGJ3BgaH6EWxCdNgirQU7oHC4mQO49peXIl3bFpX8KMFSBAVVdfA
uYf9/SOWGdAcIl+OkGWzuoerVNSSCQf0f+/XgJKjf2rIcodhhWL9LXKD7HlUmn75ADdBHwmAV3x3
2nhuxAFzKngZeNABgLIeCclw/yIuunet06DvLGWFNE50gaX3Eg9HFw/TQwz1gY5h+Lh4xKczchbV
MG7LZGNRsZJC5oYMB1YKc3O8noyOOBOzzTzLgouE4l5GIo0/seLbwUo4/+WNn5GKHbwh1cUHCRJ9
d4N6eTGoMyPe9Xijk/Pj17bbMJ8FqZOw32M47o6V0ernXH9IzVODy0Z8VLzcO3MJXa30QsMfvrcp
OzCKazc8Qx7ElZEydtBPm0nMwSqvGY7ZLUyXE8QjiRpxGF6rvlXKxFNQd1+XfPTTWnPGEndJl6vV
DfrdQTuyeRaBByGYQ8D8dLIvidnKYmGD+e0AzpGkf9AZV+fdXAVpjpZNQA7G/bkgCg98tJuU/3+i
/vSGQQ+lN7Wi+2VtVaRDov5Ss8sTLljPzr+jidWiwk+Ntf5Mnm3yFS0CYN20NYXoXAQkCKVeQYEg
QJB703VY5vR8DCis426yxRwGpbHnloBPAVM/wja5OcmvEEHZr9V0CDUtsKsn14awM9dRMa+wtnVN
CH/CMIGQV5IwfPWhw4ofWJ4LYDkHJ+tsEfX3W0il4ZEDrx/2BhQeqaKPH7PFWc/65HS/1M8v8gbJ
/WNGluQX1IKXPfAM9LZeNxugWt6HYmCcKwyHQlPcJnpVgFj6OJUxn6KQbEVawIJ7h2ey+93m+Op1
oB7PZv/Wt5c//LWSfksQj3981Zsz+OGiQQXP4wwzaIDSwpc7YVScJlbaucJXB2Aogz+5XXCm/4J/
EgyvlVeqhuF3JFOhbkev0/5+v7WwLYSYa96mDWLHonraQWBk7EkAMwpIiUaDRtQM4YV4rfoYO1DV
5LtON8jTXAsWuzluFYtSJlgO2VXyj4qXgQbjWBLI8j+XLhC+U/foVJW+GFn/QhhKaa7TR4kRv9xs
mAsom/ztZt5J+7C3F+BE8U07PCN7jYc3OW0bvmk2o3pTrp48GOKqowMhoUqdycPh/Dl+gGceqK99
rNvE16cO3eletM+bO2EbGglcfJEhGaxwAVbbTB0LpUrtnrqtNpHWJdhQ/Dh1JYAqP/iX8wkMTsef
xCsFpLvW7deaAI4Co1iHat5clM5MVm8LmKO/nrTX0yXS/BBK4ubN17rysFoD6TcWy6AQ3vL6s5L1
PxSdoAwGj8/RNtLq2RdnY+QyFig1FKI1bsd8luYEwVwVnyLnn/QrnDWH91IR1VCtRDmf804S7iwM
ni5b9Ggm8soRwYOE8Kg6pRTnm0/6fGIneSSedsX3v8gXdecsd4vqb93pT0tuIKF66vczQPMifq16
Q0yj/OuxpV2a7c69IhPLIY4Gpm2wPiS/SaBnaNlLXSX+IQXbKkl5fuqUdkh3KbUUYPB66IJmQbX0
Iv14fxO7uG7+le7NqTad9AeYR32AFmC6ApnI5Apaq3+CtgK+zRByX9oBFbSQdBJKc2LnZW9gQ8yc
HXX1UK0FhsYGwUn/e2vPK3n4sIfhC4SUVyAgBCiJjdmDC/vvqntXjnVQMzm4uQQ0QLwI0bHor8wu
Kwj80mM9jftF+n3sOlwoEZcqNaIyLaMrwCxTdbZzCmqmoGwXJEsR21ZQmozQbtJcIDqKsA+SK5Cb
t072Y0YSdvL96fuiFCnliy7GpmEthxoSHX7kMiKXiOa5AStjdSndc4ORP4mxRTahs3h9NrtMq9UY
79CYs3xjc0PjrTXo7UFT/XqYa8bxQ2CjwGKI1ZMqhaVNnXdwZR+vRXcIDkNgq+psHzK9pJZNf2lu
eY4woHISqG8+MHlmj7x3ewit3izqj+OI5UFardVqSWxEm+6XRqhNskCV8/5jpYe/LEcS9H1F+bA6
hlMVCn2hgtq+8XK7I1V3+vGX7EIiKQj2heEbsO81TCFvi3TqvmmDsjbyaOvpLBv5pSVITfcLmz85
/hYvc3SG4xvZV49S/4yVvdKI0vCLpMsmrE0DcV3UjarT/n8d+XU4A9peCtDIC1j++pPeBJgN2+AE
LDqPbUufpLS6HXhCt8KaGWC9pAyEopPClyQ/JoANKDjywZYcpp5OFtVcO25zOZ4lzYIFxq7vh+yE
MvfUMHy2z/6lh+1lZNnIwCQgwO+Nw4mq/7hdqvkkvT0ONNyCEjCjtzSwPLgW+IV19lUQAcsjEbp+
NmmpUoAF+btaHzdQ1A7X19o4oTZxYN57VmuRW2aMW64ep5DrTXRfyc9wm50MQ/3Aac8R+Hj3jyBV
oHw9dYFBgpeiKCBGjyZckfJYYIzAVuPtKNnZ9zO/qfERAlTUtnL5QMrC75ht18/K0gYA8KQvhDWU
qgxeXISQJvRW8VaVyXOd7hMJf7IPpig7DP25e3EISlo7HVpyLrvtkS8tnJ75KqsMjFKyEO5xGyGT
ueip18LaVAFtsKhrp+Yu3dERxk19meB0zHA93Yl4tPmSh3H8PTUQYmc8PrmKMkPRMDvHxMmJs8Hc
/PdRx86FLLH+lIrbzRV7kvr7ltUMxaD4LvRj1XNswz7T4wIIHpXyJK5Tq8DmODM6lxLBqvuJcc6b
8lE9VKjF2lCHWbggtOBVLaNzrxo+iO7v+VwY8wcN4UiiHiBi5LuEuNkgkwJUSuGRgIPcNYn0KSgX
9OwJNLdZImH71s04Tiw2qy+zWoh4tuGW9mDorKEwHtB/9wTO5VeoOr+DBO9THpX26xULUY4IDtk8
ZdMSq+eiTm3XCcCf1B3nAm9pDkMw3M278ExQ/ndW9zkDrqWeuJ00NGPORLzY7xubpFFeTLwQgqdl
AepAjjbxaOR7xfYTovR+GtTpYivJGqWlum+14s870KwFrUpU7YG1YSJqxbXqWTS26sKmGbW+ndvD
+GcgybcmBDQq2AkQOaAnK5O2l/VUXSVWDDGOCROgateTmwphQV2GZYo2JSdpwjC9HoYZn7Ivc38C
xPHiDReirewYjQRo5gu0nFkPAjVcyGWREgAQq4S1hQLWiABzLKZqbqFFQKjy3TNkhEcxwLtD0ron
ygDuQ3vfQk4CPL08Ql9Xdj5yGVTBeXJWbFq1MC/ReCcDwV6g5pUMLYtVSKAZDi0BTIrNxrlrIyPe
mCZLuZ3QpB+2A5ybvIgNzO36qC4aF3q5x4pVqmnNCmN2AxVNs0xWiRnMiBD0kD94cpkY+puEgGNa
dAq1GFp0xVJAljhQQEPeA5g6Z1I2r3c4dpuzPJIjb7sCLwvnQJ/kFoD1dCKHuJrNj7hWBvmeviox
N3oI2svcAj2vWHuZNeumM5Puzgp4yFibGU76To905lG7wgLTWitDXhUnKdhY6mzOfYavJt8lfvR3
+XQHYgovahL/tZf/whRkyz7LpsvYGMWKOGmeyxq9YbivMTjGYen/v99iLMn+rjP13ecAQvAdwNBM
p1+YjOx7e5A2pAOOfP+TqXqxtssJqUbNr/IrqNEmD9KauzW03EBhRsJ/SR2k9vUnWY9yJsKYynfV
ijsrg3c7bKntm7cUJACEd52Khp6BaHORvfnc9q2P5PSWFd0zY+v3GNr3Aa0xLv6tG9AZSzPDLWSI
Xi/n98uQNXZQrfaV1mOISeni0VHkBLv+wQWLy4IE3qQ/EzYoSS4QImVoqeQRocrIw4V3icEwolm9
8abdCGMzT6u1HBNZxW0pIksgvErTyXrS1i+M94kcH3UM8SEa3SvJtbAfl37bifHFgt6uHeNXe75O
rtwRtlswgHZcJneYiILzyBOO3DLvo//GhBRUvDBFNA1TL0/Uz6iIMVQGkTpVIbKcmnduKtkREN+m
QSfDyk5QQ14dwD6z9PZHPL+J17v3IbuhR7dstvT1Fuhewk+BAGFcwxJlwhuEgr/twWVqrd6Xw2I6
lfM/ZnPrizeL87fMX7XgUq7+tB7/paaxc26Rb7zZGn/JM3phUuH8Wwjnckwtiy6m19hZw3nFoW9/
AYzYbiM/ghJHfp5gO58r93nWBqcmjskvIAHFWPmzR6+AtxID9N0at6AOPk+gKRampe+TwSEA8kS7
JCyehdKFC4cMql8ymuJ9ZApyoT2IdHLfnCXusGnlGF5w3J+uEvfy/ORW2pr/3i13QMdO7BDHxguV
PwFvHzMyHL88MPPjZHsWvkKZnipbz7sRYhNC1pxj8B4/Q2VTVgJZ5zvy+PRALFOIwBegXoGjh82m
CEMecjd0sjsUb3N/acKsZkBxWHoAWaUHb85D+cihCjtiMYXUIDTvGtiPoc+3CpiEOFYx6NBjPI7P
TYk0jIQM/Njm55QqBKJCmTQo8Ys97YxNRKRCovVgT7nXyc/PfwQP54O1HWb1qSzWSKIo7dak0Zvo
K9TA5ihGe1bQhJwfuC82yRH3Cnh3A6Q4xKbDW77Tx8Rb2k6PYvIqDjcZUcQ24tDG3CEqbgRx+gcM
Q2pfbqNrcbVabjkjao5PtKEsC82pdrLwaN7d4rIsq00lLr6/P+5iGTuzvmN+PPA+56jJuEpdsRO1
WCX1oz1U6M9cMNvY4bxmiRV5VgVZIpQjK/6E3Ydve0AS4bJA5sOAu6iZ3N1pgH4oFzt/yycZGDYF
Ug4xlYSA2zHJ1IxQ/pX6yZRQhmcXHRS7Rna2EEDd95klDyxHMjKxu1WmxuuEz0JAdh0NT324DxVj
cscPbjflhl4cuzNQvoZdxxoYKylhdGCPlPHRy77j+eLgwh7I/hM7CnIiiZoRnGUv1sgKR4YzxfG9
4UwuobEOvna8BznYJDPJ3T8ykMey5Ks+I/bbJ4CSaxHlMC6S0aqoLVOst+AlGN1yeR4YWoX5HdQ5
kVPZ3jkzWfnef5au4j0xIpIv//yOtwQLV7z0zELRKoUnafhliiTDzo/HxujqjMiQk8drp8LouD6h
4UwC+C4PoTGsWfMWslZiSMnlZxPSw9zQovqEFBzQgZTkijgR2gWa/SLec7gpAgF7jbaQU59kpcDB
FeeGqv61vYigH/2aLyJbha6cU/rn5JyQf79fGdODXPQe/v8daNxyqraKMaLkHfyOSOM/m2yWODt+
mdRPQsPfaWJRM/U3GbfDDEPVqaF2V3fUEbuqvog+B9vnmUO5RXvWnFWFi7jaZ0zhMLKkZfG0AkR0
PMMPNmSVkji652cbqtPFBEkgUfWMyqKdZN92+OhoS+1492v+R7aBYhT6Dy9axAppYjn7XEun/j/R
69X+Hg51gx/0Gjk09/vIDdyN33mRBPWUS/NK+J8u+wZCjnrErdG0tYkL0i+L4oD1Fhpv8TU86eZo
B4LDx4NMtCizXicMvWO7ZZTHnmLFs/jsjp8Bagx2ks1vpCgJIwfvGtI25/1TUZkYyDTdNnnTtT1Z
a3dov0ZG4rXQIRlgnCrhrgOklYpfDOUClftOltNqAhJTNvccqL+d1w8D6/EXuI5tdc64YNpcEgV9
sYW7yY/y8INbYEzzC9Sd9AgRvXSzYu0dJ5fd4GHE9rvt6lVvNGz0Mh+0U5fIqPcJcO24mFlqmRI5
CAN3Fn/8e7118FWQRVEMwkeX5z7uvD/HkVePZFIDtvpSdGy0mYpdYRRBvb2PjWWToe+awtjXxUT3
VHpH8S9azrQz4+ly/nX2CKH9qpoPdRrVvdWRyp+QNnB3n36TfvwLJ1SZH1eV6R2UTLZg1AsHvoWg
xsl0lxpU/3iuFouqAFuak+QChlXq/FjHygvQ6bHEke9TyGlordzetfDJFNt5NS+aRj8XWJSwCo9V
pFhcEBYbdTscIz+lmzpqv8VdSK2rSTKPzAUqwmSg0uTTqbZmmGFIN1Vzfx3ciyBCVDwZahKQDSwT
/qX6UXUut2uxuRoEo1Kxu4xTMtufJzVaRlBHkCu3ikFqRH5DTM/tM8trSKh/QIIpGQoihdWYjUIk
dgXjS4x5Ae7Mxy5hap71wir6rNYbSTq3nxEPz1ihmiWiLgSfrukuOFoKrSXT2vSf+6FGgog9H+O+
ByaDmJRrnjNhc3+bZXI8KcxlbswJwKaibY3axVOov6qqVWQExDpF1BTD8lUDQU9rMIq9Th/WVgSj
EPfx3M4F5MqJZTZCzbXw6ADhBb2QsNRfyrwYupERloJjTLiVlcJZOoJfCD4VCttqeV+e7PYuVnje
nvmQdEjQTf3AX/0eF1flJBvR7AAQssuYHMmYR+mX4vPROcb5qKaC4kO4vO3PwOvXRm8QpTKrVvBU
w7Xeq7m+VXiwkOqhlImkdXqnkUPP03yG/1BaVmHVV2b6rRW2ocQPgtDjRY1vEpdzSCSyvoy7TZb5
lo/T5uehnKbgYkMiKXsMOdYPVwm/xFNvoTECQqBxEMVIqo46saEWgnOPJYpO84C2VEJtG/PZmiX+
FDGj5pzUr1MSj4zEErWVYiw865AG9Q8lKB981ZS5VvUabbZZW/zPlCGCaRxCWEqwnF0PGAeZCmHS
XdOSg2O/pHdhnnnEuzjrfNyB+J5WND1Fqfg8m74+4GnHcEx0hx08wrZhoUiv/0kNxM+Wl3zhasuv
Qi9TqIGMeafqtTVFzpZ7hQxQlfa1WqFuX3sCmTIN4aSaH5XhOph0z4DOUQ+k608uu+pBD8+CUi/R
YYw1rCC+a+LLX6YECRuqi8XnkTxbfkLVYRu8KHN9Y0Ht4RZ1nl7jbuWbbo0fGl0xe+NiIKCj1okC
deXNjtD68oQMNWWzvS5bfUUG/kQ8y80DsoWsFhcCvBLKdrIoShLmVSEGL6tYQ79F/vdOIKA28MQ8
2K3JHVwT7vgCXCTYo/N4wDbhktZSlEvQ5+rKXC09hI2jHKWKExBadKwm4DDLSyK42vCoHdnrCIEs
HvBrbuX8/uHxBa8GDSD9fe19vUCb8xuVQnJ7FzAhFm0WKh/n67gsPsU0jM4+EYDJaB4/qKrUM8Ki
ZBz98BJ5W8Z4S0srCSuAqYXtibBw3ED8yerGtcEKxUV/j9HD0pIT4Hc7ecKiGab/9L07HTOPE56r
yNcg+M1hVmbjrUcysRxK9kHnUgBX9INwrZrpvFLPWbKNQQkwaYN21t/cOCiKlEIRYSAjMct8kUxH
6hJzgyKLKSoIWgct/T7h7mYKFXBgv3naCmRiOQrKtqN3f1o6FXBqieNFOjHfG/rbzcxYDcGXbRAd
odYVTdB92zbib0YuUax8Ns0yVWovuzFlwuiBqU/QuWC84JTNVCbjahg0EXCFPSt1I1mp61jiIR+h
GHKS7DXbQxB6xoTQ7VEaRDfGaUyH3f7VungD28SY6rHfT/5T0NsS22ZFA7/f1V2kH42ypMI/iSPb
tlqrMDulzcPrr+TsNiqoWrfgwzBXD9u/6vb73AlstrZhjx8qA+EEhpHb2C+3tRlp77CCRW074iWF
dYf3EJ9ZNpyIzBmUKiLcuZDl2zSrss4vT+CCKT/BsaDCMOvTz1CJRvjNGnMzkz8lq9VeRV+URgNR
ejYPTZQjspOVd512JI1RrXL4Hjl91CfWNYQPIYc6xbakmiZRir5CWaggdB5kMMKnuhjkGNHbIjmn
bas4/ecx+Y0NqYp8BwnXN4VW0EWMZIrLtymFSqo1LFcVxme+bwXTcbnhvM7xuiIvcuemO8nAAKo6
TCQMrDQBSTP1G8JgvIWu4L682yxrKlI3UVrjEFpS1uQH1IBeLMLm0IlBx13m/6qYTRDeNQUm9Kwe
aAd6/bG/+Zx0tmF7ceEPBRrPST8aep+RSN7vH1gypeEq/44UunoclHm+SLhePq+p41K2Qx4VpGNT
BVMhtbdULtdH6UmDXSr2B1X9jW2HBQoVctJNavi213R3JqLGyxiA4+O7M2kyZD3awOuSsYp+1Yr/
jvkCBRBgg4lQZHmNVTvHbJoYdLwo5SmWc1LSKebfrl94O+86eLbiSGejWUOvIRcH9sO8O46BlNCG
h/m3iMnQgVdbwBPp7Le+e2y/wBEbHZsNZfn1FoQHKeTCf6n6OQuRSnpTN+o0PPrd7qdr/5sYjajA
8YnPNOz1drGIsulv61o1lRipWdjeTeOYfujA1RrjC74ofMcZlgJcRlUjVBXKaUJmoib/kUu9KCVV
g0omJkNlEoC2Dw6iRBZmx6rsnLh2ZHVAr0Bb7mDNnF+xQBnsup8WPrqNod2zsIxLUd/tG7juPttT
xFVrMf2HZ3qGysvxaENnRG4xnY5BkEkmRkMVAXjhseSER93j+erxWo2ICfk7dcP+f52RiC7TLj5X
e3sZxnY6/DDWe/+ayIdBXZaaoyNHARgnxfSNqgWSGaprhz6YedroaSLyXRdD6YA1LNGkm6oOiS4m
V6xp9isFRSDOxO7PtzrfM5PYs02PGfaU7Zi0Crz7oqrqTSXMH6MmFcLZ574EYakV3hB2q+JyuNoh
B5l1s0O910jPRRvzE22C+uL+wZv1MFFum2Ux93ZMNFrbry8saViPQXPSNu7DOiBzUAgucKidRMtg
fUxO18B9rSJcB0AXu7ZyYu8TcEaiorO8OZfB1GdWIlxku0/OgKTnJmMX+7zdsDxNdEN02TNJ+cGf
W6CPDUFDR1rqarOQQowLPzKBfrsVdzA60bM0V49hBdIFnUBizMyZ8BS6tqp1UlsTbcYwYXEZlTL9
roqM+9tUQETlsdZ2JGT7oiJIXWi6yCmQbSGXliJFMiIKhu4cpWuLMjTO9Chh74FDZasQFfIF+Df5
DDtPiiO2XbCCtbOFzKEP/yaJsdOj1hIxdw0CO4q1AjRNdcFCDOzMLV9vAinuoAo4RNimT75Sty+2
na5qsbCsLaWcUhCAHrEyQ41q7lobOiRIwiHN+vvVZubARjBRdikq++q5e6a7M4BgvhwyLPy+XEs4
hPCRHTO8ttGgu3rsRvl+A7230JU33YhxI1x1TcuTNkUx8HZ5OToXT68EJ+DCjjI3FRHMQzkoqhAY
SioCtk2g9cCCwZMRUq6tFTcSwJLNdh41iha6HdWtgxT6kjIVinFX7zCalQMFRB9vftPmpn29uTob
U1LFHtYn3PoIlVRz8PYDPeMtV4SUlzNfprZPqy1F0c5UJ3RKyFki1fuWrxzkgXpmUqlT32oBQSJq
9S97ZIdzXbF5s9iz4JOOD3hKqBr6XSNXbWZhOCFWi1rROMTc/Ew82Tz7WmK3saJHvT5zzg1G9720
YFzyhx/i7ySEgc8mym0okCboM0YiWhng7cAiWmQ0ZEpYvoZ+BBBmsYIRdEx1lAVBuXP/Vqckk1RL
t6Y9h+bvpIMqAraTRpdehOgquFTMjqDfuOiDtOqtLh34+PGHwlmoEWhRF0QDtsAUz2S/3dk8BZuj
V0dPnrRTHWJPDSNdRMUuI7xt28AQ9YWM4pcw1FJTl3rN69pv0Izme8zVG9c/xpO8mzgtP+mBahn8
HfyyIvEEhjKWmMv2gHwjCqFhJua2k15y7OAVnadC5plzGNl1PbqRwLAtWLial7ZSOydGwsty0u1w
d5n7+4/NLz5EKLOWaD9rWanSQIIgG1x/bNyk1HaHCGlci34zMlMUfkOhUKf+o8nn6UZ+jcCRuQo1
zQ2uyulCoBApRkvyyNLQPANiq7WIyd2U2pWLakhY4hDqxgN1fZX2MgwQe1AicDA8JYHvQt1UagED
/ZdWLh2R3v069z4JQE5qH3BF8cplggNCR7NOcw+uubuKihovyP6d6TXTY7I2o+TNH7Qsx0XozW0E
l91SZuofnV6SHNWUxH8CQ/X115zCYQB72ten8kHzN1L2ZvwkiVQL4O4cn6fI65Yqn9mzPPfSGKHv
R9niWysLKEgDu+M/ONosHfTof1KyVHq6eqeEKy/RP+GcfHdN2rtGC6+/O+ZRoompSCNr3mYC/76J
T1yfD8+InDMOD92BQ3XnW8PDP64Bkd8FCHo5YQ8BOdEvB92AjfxEH9tMp8PR1LAataJ2RhrLu33x
ob+o2/in9UF+/QlIU54U7uK6r7S9V88KbDBINHMPsrHXQCJrA5vwaLmiM3kv26VukWtPBDlilbHQ
Oi191j7bdj1t6zVKRqwrVUG7Zr95+lqx77HMOom6L2woIMOHAjn/XnMmRvAEQrqP8RHbc5rZdOSY
gup+g1d71zzBYx8Um81GwsLCkG1cU2B9/+gcFjTWvkbT13Q1bRP/filJK1d6IHM5ZI9JuMuy4tnL
yPVGBDOAxFOo+15bYvqtOahvmJNqPyhSmk8lOJIf5VwHkKuKlAmlue6MkazxF7Bi/OSLmddhL4aB
u7uNW0fWH0dAPwsvmW4iVfRWokO1tL5NtJG8WZMfFjAOVlxTQG63Jm7GM92ciNoxi0KDzkZHDQs+
fecedZ7pV8n85qKDRe7HpvIJAj4fcUtOWvQeab/gzKtL4VgXxJEsxxcI0g6J+AX5PameI9AybJjw
BsL6oVuWZgJ9kEDWYw85jWRuFEQujgGD+TjZXetw6sxXbJN3Wz3/79oZw5Rt+MRPrgexecwmragt
WngmNqX6dH5o2BwinnEmF1XwUSy7+koueWcSIg+lpzgZiPxlxLn9jKhLzPElx2Pwty87UZjUQmK5
LgGbIg5p2yg0lebWubh4s/wUAx3diEtAH8kbr54b+0SZ3gLkAmb4qP3JSapqra98i5L4mqoP+Rtv
qN/9R3jj2R2yn6GjHpGEgmmOGCpKesAaOdEl0XA3oE9FgcIMFNzc65yaQjGeWlizqwjKCzYEX4py
KIzXfqpGAJEKChsXaOdQnHXjhduSaSvk2n4rRxAWYoGVJIuSewyQqSeH8NhuDIHSemm8Usmw7pb8
BalJiPJmWck+vslEhKSzA0kZOWuE4MMAGN8BOnqR7vpFEI/oOUBguL3gh/NK6MPXaYNFxJlHcBa8
akzN5wGkhn+t2ayyr1X9gu7Gc032j04X4zOwhi2VUTMOvflnM6siDDqILVLJJ37vul++mLETtO6S
efEz8dTRQBJjiwZjts78ijcBFiWa06TErpuGaRxDahfJZqsqBmdh+2mjkTdr6SZgqwBI+lnDCa1e
/7WGsK+TtTooUsoSZNeVk0bq6YLvKPBeazL/fG6TVB1TM+2xMr5jzj/fyl+LKDnXH8a0YDrnYZS5
RoY27vmoBPRoqcL8o6qhdKhMEAyBLUTM9Lseq0g5hUekDHpdZ168BIOE4YKcqnxiyJ3ZVdphQP0e
RTg30/G94gpiUqmKpwS3jmHE8afo/ZZxzk1gnqE8++Mnb1qcPfWZQ0htM3Qt94VXmrbzl1qlhPKj
xkoqZoFHPu0DMPPnWs5Il/q+TiH+n+HzdOWPYY4Src3grRUpNqsNhPhx4Isw+zZOyA5HPQ5eeBsn
f6DIeiHukUhV7oRo5pMOtzpnqq5ynueiU2uGMsEQPplrhYr8Rsbwrx5S9Ky65Yx3V2hJiYHqTZfJ
fI0+Gig9cKd6g9gXuMh0c0eoChJpA3F+eWLpyV2RGNOT8lMzeKqZ1+n7CpWnWA3i7dHqxBiT7nxA
/BSO3dMovicOP0N1rYq+NE1O4Jq3WIxG2sTkuM9Jb+7fl9+N3lOyraK+sIbD+Kqf4dM9GF+YTfYp
QklY0nUOfInkqrdQtc7VcFBXgBgN04OgNyE9Lkf8qWtLDwHsiDuNg+WfeR2RrWmWWaF/+WuzPmB3
uZvnjm8lpDwx4Va/WNW1bo70xCQWLat9TnXBjkDHGahmIoKXqipxDY4v9OaXdX/3rBRcRS42qbmD
haNSHJtTzHrXsHo91DYZdmP8oQdz4hmcFQGK2LcRDqC7HZlmKvmGs8WQ9ripfUDpd4CthkgBEn97
Pw9nooRItU9AsTiwkxDC/WAUtXm3G1Yi2g/HW4bwEZCk3RhXPq7fmMC6Nze79WYa4gOr2YDufGEA
an8NVB/Kp+5R9on0rvXpm3RGOTaVU5FwG0ubSp5OXoni/l8yK0IYJi0xDx3CiYstVVdL+HgMA5AY
vEqCrrPRHg/woTeGhW2wbESOarfVIaBnXZYpm9T1nkb6Yu093RlVxPMd7xbl9ACQREZnLCa9jlEy
+5h7mWWjUDUa07aGQGrOEnk8GnBx55hH7uhN42GFxCB8mDRTfhchhrCdx7xCLSUPZppCVP7Nyix4
VQhpyVAWdYCFsx6aVB6QFz3T2l7fzUSl0+bNCe+PbnGWZlZ9FIAYkVGSdSgNwoGKuMBV5sbune8h
KoKvlhBU87GlZcn/laqoQubIvdYvR7LLX9fZjfxY7dbm6AHwslW9m63yVKqZOLjMdKTqms/K3YAd
J1J8IsTr7AtTK6gy0w3HBPCcsrAlY2tgHofv19/syUqtz7rcSSNlux5t27we8MaEh1DixXG8Wt+e
1nYgKFmZAUSiqrYWHXKruKqPGzMnV/F3/UWvo4N5dqJvIEhB7xlJjWhZjZ/KXer/zur7mDiDr82t
aMhVju9rGBDQqSbme39D9nxAUPT5IPNtyCF1gPN/iDZHBA+2bMSACtJ94dPiKpoEsix2esE2RTei
5iYD2Ri1EW+ga/thjXUbpgI0tgwRHcOEn8W4zjPbymtStoOsmPYMH4hbsqtJj96/isvh2MjzE+ug
PgUTUQd8auRTnt6D/8mwiTDH4TXkXavuPEcMptGe4HLgnEh+APf/a/lYrrdZB8LDLlsMy3eIWYeT
NYrsuOckZbATI1bdWieEQcF/nWy0uLiCTqU7GXn45J1SYbjYWWoeaGR8SN9ff5mK6tncrAJQsaC8
ZJhRJtFUw8jnZH2oemKJD08jgIt6RwIN1JPiaEVhsvdbvGetuOYZUYcbBEtAS8fPOW5+qi6iDToe
91aUudVuIyz5k/ESLAinADCgvC9Qf8tWXff5Rf7n3JsjVBTxAvJY9dYLUJ6SIVKIHBH/iNsJswDF
Ude7rgybL4UB/r6GrYe4WBCFW0Yu5PeXOKuH/XkuvqDlIe6DSXWmuDZh0xKzyEzPkobOd3PwzIjq
wRZWhdbt3mblFgal8lKVUJAzkXPC8j8SuTDTsSZ4kRurTqdEt9LlIkUtYDD+5uiSAvaEqOTRa9DG
tafkcTMMwhYKHNtBBCOFocbTOjeGS1boniiEn7ngzpHmJrGSSduht+EINhYBHOATCTMswo3soAYw
IxCWb4ianIDx+J+18Ecu72wBgB2erv51R0gIdUOxL/O0ES3eXIvRKsa2qVZKTyQw/bRIBOZvMJhB
tNzAvIn+U2Fq1i/THgQH7jmCWmPkjs6IYo7UzK9M86DXBGKpoKlxjMTKosVG9AU/oNcHuIFpEt9T
W9FdCpqieJlU3lbd3RpqgAiBdPUHrMDbizEqD8TadE1iBr0BJKUrJInU1sYSDjCE6XTSZP8Squ2Y
CA3cbS31DQVQI4orQtNDmFNnpmnoxga91VOjLEl6e3lYNlF9I/0xKWfaNUTY05CnjWLwpG+dtotq
Y8+R37PsBKD3ncEXWXZNEMVY7aicvVRyumwG3UbbdwsLiB8bSXLqyNZB3bcI7thTQRjlVG06nHts
If+1hvwteBAZa6zQCVaAKz5uDxPT8bSPKjDXSgtY2lRiCOKNYDx33Ye2LD+1irfLGB1G4V4Fspei
wERDHUifXiSJsb/fs+QoJXiAo+Qz/cs8xap7re61SaVPP2AD9XnR2MGA0zC1zXSXFwUahRky/gAh
ABhKGbQ0RNYlihw5hf3ZbM2LRzCafOoSo4Z2yioXjF3g1iWrisI5iu7/4J7G2RC0gcb+9CosZWfw
ZOeTx1pF47OrjFYSOnmzXFKXqKSJHupSMU1A/HqHzDlW9mK4+/3k1Uvwi9bHwDvG55y/Ajhj8Uzh
2Uu2a0prEcngdpsLmFUf4+fz/XXh3EqXzAvRQFIDzzEFakQ4xMEyZd+HfsiwiIgFUBXxaJ2Fj2/9
g9DVsn48fba9/5zfvgzhDxOXiMH3vawzaTDYLc/GRDHNdIDxk+Hw9pjwPrHlpW9TtlupZWBu8XZr
GQnL6q4zxWF+Dydf26LmRP6nvabTko3TMVlBnkXubozW+v/wmPUEtGI7xv1t2S1gBb7Q8ywTnq0/
Usu4U0GtMvXSN0ywKkOfCq2iY5/AHIo7LPw/ClfmHM1fMNfZwRxQf135SQX9lROXA6+uYlNk2RI8
xSu/3JeBKdpmIA5yPDyg3gJ4l1lCcG9GsX5cuE/PXeCZKKr8FvScV4+sDh6PXsDIlyfvMqVN9pOp
uQJqWKVsKHHQZHnhzT9/2gZrxNBGxNBJCdj7nGs73QGgGOML7qIVMTY4ZX1Mfq1rc/cpS1ORdnGU
qgFoXjfzNN9RK1da+2oBC8VDET1na6x8w3vJ18EzCn2jN6C0XK7/6t5ahdDxv5fffzbzm2/OuMG/
WSc2QLgkQKA1lPD4aSe+nEkgMiJofu430cnoByrA4DFVNMdbhyM+MOiGQDrO1WtqM7aohAgALTwt
e5uUFtZbj2Ri3PMj0SNKJzhBavDR3ONrj8u2kggZEtO559IMlVMpkMz3++D4HRTwxViiIEQqgd+4
uYISTffCEyBVb0I2dz9oJwBk46pwUrvrbGZz87eH7p6dj4qHO9AmNO9MDOQ3gUB5A+l9W2eBl+Ui
3nLpOF1YTnRKC7qusT/GAsZ/P7oUBYm1Yj0jsUXzK3Bd7TrIK5aED+s2E/4PYvG6LVbVRa1u5Cgg
RjSIUUgvCyBEhjBU/dBZk7Zr49xm4kCyyIHoItU+XOsf11SNT8LkolIBUvvkKewbG2tKOnMzndoK
TF39UXqgGpdDWW1B6wAbyf6be7+pNUFBWX0Xp56F6oLFaZsS7fkzRG+hs4UPQhvv5U3DIXpUMluv
KQzbHZIsfSr5vhzqwhl2wuTQ73dhHwmm30A+6MTmbQOQ3q+dloxzH/Xx7TRbDtyWFGCuwrgx06Bn
U+ybTz+a3z4ivBBRqWv8MSHHfiEdaPMVmblLgJSO2IjMzygnYBqoIwlT0NBlyF1T+Ygsc3u5SYZy
fx0nkEN82MYMxu1Owyz+slw7MR0q2j3Kz0lJMkdkAmGuCDWJsHzQonjunE9FawXlS5Y9GwviSRfX
zLmoIjMN3JAR+sWs0DTSaXjT0YDt73J0M5EU1prN+eejWMZk+LTEa0lvzJLLQuDaWHU7XrlNtguG
/LMhq9U+N2kabFXMvBnVQ3SZbLXVkx5/xKe799J5AHfE+NNNwoaEEIwuSP/hYaMQUMlOABGNnh4G
xCFvQi014YTsloCBoHdOGIfIAKLBUDtKd1i2kMMnW73cGdcB7uQrhOtLJzZwmTJb+B5bp0NvH6S9
Rg5hClAQweU9GUyZz+c7jfwgg7g8spdGo01mTQzKOkg+Imv5vRSYNH7R3Rkh9/PM9ARnS6dxeYwL
1Kx6BfLOqUsnqQK8ZEZtfmJ6IM25zqvmzYZ3IRBUQz/L4ShCB+K+H1KuB1p+xlldH5UjUDaStMrn
OWMd+UsqracQxr/1CVnODNZ++HoMltDxSjdfFXC6z//UZKfKsV17Q4BeCZuXBn/JFxwrIikfloTY
KKcGZoI+bcFVn2iYwx4a9nnJa8/4gpHEVTjiaNy941ywVKXeZayqddLcYiddFkTl0Gvif1tymFVS
VWUK/5JbbcGN+RiegBDDoq9hdWPrYt4oTRGKfoY74bvFtdMz3fszyDHzg9/B4hHNuh1VPAYPtcRb
A90D8r1ukb69o0A3nPpVQen/pxXONOPcr+UGLNpefGCQPoRd/8DBzvdvc/0dCE+uKb0t3cvqY6+r
cMHGS/f5KTQyz+lQCPrRREhlV7z5rnBBWlyX06Hg6BdFXgMFFTcvcYXOAXi2aYjGeTHMR92xC98R
QuE0Gn47bC4uB4iBXHDk4FLiedU8bPn5AdTqeqNXsCO3lQ6x0I1DHtJlAx7aaILUF20Nu0NT4USW
Db8SGBMs2WCoUBv22EfC3HkSXX2SLU+Pz5XKeJA1OBUUKDRf8oLdqgwmQY661qfbummkZXaDNSFK
5wqAG7BIAbxWFAXOiUheY6QdNAugbiX+XbszTUSAb0ftPhkLuRFwqpqO2vyvYlaMXKAbU3TfHjsJ
YmaZYpajvI5NGNTbGM81b5631JwG5RAH7poibTupNvVQTQWQnI4QZZQXPk7i7Tq8DjdwvL9cjxlB
zA07CLcRdrsX/D6M8IHaK8BTSAcJRF2+sQED6AtXP4ZXi0abIQ+ez9JLYVLOSBi6L3SJwNP7bWhv
B96esJBpBfAVUE7HBLTXrB87CwHKzbsiWH9Qx76OWsyhg02FHBXmqSM3d/HIz16w4XBNyh0QWPbe
enL7sPkK280y+Lb86umxiWUmB1cGV+6qPtUG85q/VC1jS16wdix1KEj+bcT8NWWK8PZRJvubDp+P
bCNAW1UDuFf9cPYcLlMqhJix35WvaVJ+XXBH4WP16HT+hKgoFuwKg1kvtJIOwgDwBjL+aD8r2nx7
erSZ/bKgPCMF70HgrvceHmR7UM75ZGwShyRruL4Yuyse2Hz2HOl8zT0QFMLIpp/jS2uD/U/4IQob
VgBm5D24wkXG12QKknjhK35Rgkox/PgXpHGRrZGQkTMu4luVjfpF6iyT/Ma5zB7g0u3KkdmVJIyN
LEDgsJ0yqmRDz9O5aJWqyymWRswfTsD5Jm+4lbDJUxHtBFEj5yTtakqE8sSPdeK2KuyFekgbhjPH
gWTbaUgC8rHm5HLTGEIdMXv3mnm0JFdm5P5ZIsX3zpQXyuINKIVPexPf0DHA95qmCc+lyKkfnPxQ
h9nhKCdOc4dIZ4Gu5owGP930V2tE9lvpOO48OmDp32BOEySU870lEG8nFyU0xYwTe8u38ZK+ddjl
tnDNotoVEVV7NFQZKyPaH4WVlcCzHfpZqYjwAiN/H3KlapK63bKNP6jHrTdSWaU0SeLqWvrTgKZs
xjCZyzQdGo1kjd+lMeFym8gZjsQllKxrShAKbll7vi9e7kg+fyp44kwiJKeW5mlyI/NiY3U+6ZJa
7yDTwXG8C8/fZNqg30EGsSCXLikXfecA3k6iIdHA7ygSyg2vIAaGMjzrIjJ39Nq0U4dAilcWITDJ
/MuR0AXqK3uqc/40qQg0UVLOAOgWOMMqHtJutS79O+FSqqqEthiQburbity5smh/A2/8Yq2uvHYl
dT0UeERSJNjNkX7jk/rXN4/d+o7YSlhzLvCLuwmYwz5o0KGHegySbA7D/lhJ0sWKuZyytfGZEbEB
LPABev0CS1Bgg01ss/aLIoABVy9R5kYcw/lywk2rFOLJKfW9uAQ7Kg7NDZ5xQBYPnp/8/SSrS4pP
ZXP/4suvMYGApJg+KXTONVsZMk0yqzJ6o0yUV6a88inGRSegr84nwaHqVQVFuZnKlSc3bYtP/G2L
QNFWC/diUSD7hKNjaIIyGkgpVtqM0IflneEL0D7Zsve6U49MPzYlALiczbfQD9fWuRcefVkS/Cqk
SWqeqVHvHiU/FyUFhd/2YJBZGHFS3+AIqXCuaHYcFdcFLQcbC5+9hFdFsBTh6J9FM6G2oIv1+nv7
vud3Bhug7GtZoIMOfJI/Y1RFAuD2c3tVf7+/XyD2sHg9QQtufuhSQqaytabzRzgBNRgL6PpmQDio
3Y15DPFQfiAdaZ+rpnYPM1jHETl5xqCsz4cxKaEaoTcyR9HQrxfTRarwwTFFlsgUrpLeIFFdM7TT
avSVQAJXwyMJodtVT4l54w9j7oYC6kh225dvJiEglifjBjIzVrrxyjlaFCydogO41Xfbtq3itOLG
vSkK4nA0tXh+yhIOk3s2U+EDjNdCsyXcvFkBbM9D4rWkzn8w6Y+SLF9BL0QuO9uWHemwINh/NoFz
InLA4GttpOffe9D9EFlJ/H+8nr1XCniXL1rzSZBmx7xYNyvTYQxUw9md7fihAZdzXKCBQXRn8ZEI
JVwK8Db+Wg41eFmhANdRrQDBzYoyDgzeGxpijZpPwUf6F10PMYAarNcdGkJDBj+SOikrbds6w9fV
0VzYkA8zWACiId/ZAYPQzkt6i4gQHkmP47HImvAZ6cOzKIwPm5ludkBgSU9F34ogl5brfIx+SWbX
FmPp0vzm7gerbLXsyEBYnuFt114lBRaLmzL2A6a7f+ZbUgCb3pLh70q1Y9qY6Dw0nvKuYMX/U9qZ
YMKfopcis8SHi65EeGz2T6KRKHAQeLU4DIpt+Z5lVaqAFIL9B67SJgtUnPAX43S7zCYtLNypUGUt
ISelPOpyF1mbq2VruiWnU28+7Tvsb9piCL2VsnMNXeM1ZXztf6MytcT0aYS+laDRY/PlFNq8KU+N
8HA5H3AwPCabhWh3DXlKtsbuCPOxLx9OXDxz2dn48vB/OUXNAC0s3LMliRMbIjLYOwQGQfJqNhSx
JsuUwy3wu31eRNs0TU9crP9lF+Ctu4/5nJDha3CsKxCFryT0d0al1QTHp9atFf26eBK/JhKCmwCQ
VUSIkaYXtiRODFmioWWk99ZgT8ZaaZ34DuIkoXOiT7gfmuqhQ5UmoszfWaNVflT4da62C6Vz9JB1
5EgEVXtK4ShZJJF+4mlVmyorCUAc7HCiVgZM4Vyf46pq5AnWkB2uuyktn2MfMoyPuaMU54V+AeQd
uKXVWDhOeQ1id64FUH/RSuM3Kzz9gg8Z0XThwkjYxfDEcbE7Gwmrla9Fg6UnF645zQtJQ7kB+zIV
1ynfNhOeufDcyc+90TgPCMFX8Dk4scSgwTa26F3Ln6My6axs1mLuiHmzjeSD8oxeKgWIwvG9rmpu
oo7WKWIfVk7Whx7dwNVszCA2qdVAhl3qLuckHmr0GaG0wWftR0SbyvNDd6sIwLzkkWHRfasY5yja
Nn/O9vXZ82X8XYtWkvO6n3V3Sd2aUi6QlSLEYBGCd86kZB8SEf3eUBc7nvROZnD8xOkPOsilZMI7
ijH8p5wXteJ5Jcc2e3ZxnglVBPfBjWKI0gVbi+NYLwxABuVbNbxEJ2asFT3ITmgo9PT/AEx3nwBu
Ia1N+9nC/NhKGJbhNMo3SpUrV3PnRWMO45b/0O7JHX+IVDnZfLntqHu0xJzYYrt6i9izMgFDJJXw
NuCkL69u20owh9hTU0FjudeSf28c/xALDPsE0hoMOKnKWT4cn9aMSBa3JhEpMJ+7kUL8+SgkkMfz
6dZKJkUqiXz8l9II/TdMtXgp858se0RyNgTLG9IjO+AMOhhAPCHiPv7HFudhmc1c4B+S/lY7UuYy
SHc6sZyC7CTypUasZnTdt6pSrlhZMMi0U7WoR3DYh3flz2fNgOSo++KK9yuPfdPZ4VHLFNyFAv8N
OQwwpeH2bIKR/X8AasJf5f7rV+ZcjrecVeZwcxiX/Q68wvd2AIO2rAk9DO3JSFiJn1R/TEjtq3N9
i2bYUQMJt1ye3YimCGJdqLaxtAQEQsCZfLT7TFYkJrjQ8JljqD0zGb7pQ1I82CooFQl3EzO699CV
bnzNg2LuZi6Gl5DC3Uk6a75w8YvFV2Q3cgpd/t47+UVSXwd8D5AB8hIzUmzBD64i2WZX1OJBOUnW
5mNWzXWQqu3J1cdVp9E+ZQ++ZkhpG8t4K4e+/1QqF2ZR2uy2Xe8GXO3go0tIrdSwR62Ieu7oc+r/
Cul78ZoaZ8KUt46802wWsCgFxiT5LG68EL657YHNcuq0mMoiw9fylbb8eKT+aITTiQnnPvLP7ZBw
fY5AJ8p2mQtBKxrtjW3K/lUTQOMjvCju9sUFc5+5+E50FqIL1JDCH7Tf4BMLiLdkl3FostQQESPx
j3angjcsQ6TjWNPYQwhk8B5oDovOidXiFXLAZmgLKuDuNwG3RomQmUfN8KXFHieMwZF5GFPtJRgA
EvIR6/J5q2S8CRFBTwFQkbjS6beGx7qd9tU1RqY3noKNzoFRFea2GziaXi5lGeFDGbxYkrzrvMVO
AbZwnOK7veYFiFStR+vTqXL0f0NT/c8kanl14w1arGTjOEZISUbH+xx/Y5vPXx9yAmjd86wLr11e
6w7QKXolMPUTDu5TiERiDFMYF5b1fAmwVZT9XwDuF/1L647tKm21Zh4gFD15LxOnVIMS3zJoHhHF
tRZNiKwUpw/V92gkm5ayL2sF6EG2HWw5lfq4co1Mug/9Ab0RYMqLEdSSW3Wfk3/2kpiu9oG3OHMF
Ex1v6eWBcniiIHq+facDZyzqkylsOhbh90dyRORO+6KSDuLtUbsrGF56cRybP+JzR7nSZGVer0ui
IpPalHgIuGc3HcrF8dRqXE54+ZaYNqpWSFjwEQJY3GKgF+e6EWfq41JmqsfTXPZbd0HMva096pU6
8k1AVMbjZZvgg6ja4MSw0Tv4VnnzFNH0r9fB1mfRVOXJkjfe6omacG7qdongTcwtPDnR8e1cROXr
Ya+NRXHFnigsKTRvAKL2AMRUsMtRGtjYLioqGUTByuwRfkyIYyHbhMI2huHejr/lGsbJ6Z5xDYMi
hRmCIXRAXOmfwOmaSZV6yEGcR8eJ2T7HlLpgW7OBt2cjXXAirPw5Czw3gx/In3OPgwki6udbqjOO
D2WQfmdccoTbv4IZuUoCkyJ9rYsYBK2MH6qyT3G6Gg5//CU1st180mogb55EpGNPHGlJ3FrCDi7v
MVgekmYY6ty8XtyaABEuR54u5dyVLbtcLmSfl4P/po1bFvN2Dior1n5aU3Ch+HSDgsrvGm1Y+p7B
boUN1GUCrWWJNYiuro/NLwC6BAQk1oJmhPw1DvYhi6zTjCAAtJnT1i/KhXG6dmdQ5le6g16u/Ire
HFbr+x3x7hjiaDA26ktqqfsXa2BBoy9SBTFR8fOjWwulouUeQE/de/NwmUpLf9B5Lg9VeT02yfPz
/LKrnORboLbVknfO5xZhEZIR2WnvRWJ3eCrEKqYGwXqB/7IJhbGoIoUlcrCLrhRISNKQcXw99rXN
eFXdtAtMqp4kYUjU1kvHv3mcq5oJtoM8aJLbSPE5vt26ht5+Hg14DHAk90V2oJ7Gw94Th4TjcjIz
6WXYIzgkHhFVcwMqJQ7xPcoD4pOen2ZYD0gj8gsxC5TRLkfMQbHZuS6LO4bR9JkM+NMZq3vcEWb9
7Swq5CJL1EMkCdof75ZZfKzTkgsleYDLpgZ8B/N49AMmKYkT3fFomoBLq65fyoPzK8gPqMPBlfSM
e321LJejD+ku78DgKNLD8muBaLbEHAvb2H0EaN1+BWntHnypJ7/oM7tYk2jtSp1s9nj132Bsu46G
hGgEOJKatfWb7M+29gzjm+YYP1Ldgpx4pSXL7VGtl3D4fQVUdYypnw+WZtJF999VJGt/fUPJHIB2
fXYuK3TccejqA7MDBIReMPuSu4im9h/xd2kCoRYlEagy/W9bJMmZKiQSKebgLDehEQivIq22Nnta
JnnGrJ16QZx/zwV8H1ZuauFGrvuHC7tihjNHOdLCEBh6E/nGb3jqjABUTaBPy9+jLm6WGLLy2U/O
0AXtI82OpsZhZIpJgmFA6ZVrBoRsTqaKyvwM+dyy9xKX3auOChxexsPHAKTYvZ+SWcltrvPYnXvb
jCsxJXRli8lrFlmRvEr/x7CkWMGGmNpDWO1Q27lkrBLQEKYx9jlU4xG+WrImNHUiNUgiw4wNM53w
tK1f749GwhwIG1o4o5LYpNfqyGvvJqyJ+B+vj1uNlb7pA27jvuxhk5C6S0UMdkiETJvvUknQnLha
79RU3HjaJZ/1nIj5JnidNnggWMQI2EDG8Ikd+0Q/mRrD8SpwQiBcka+WAd2eShRXictuBB/IwBl1
I0bQGJJwTHfGKu7ewM7RWbSLquDOshNMACHTVxiB5YALzgfW+OmUzTT67mw+dMEgGUZovzf5w75Q
spwIyrtDvj/MqXmWyIBeWYge2QOGih0U7cM916NgDuvuJ7N5agmgp+YJsVUQfGGy2+iMbYAZn3Kq
dGZAJRPKo4aSzADdBt0+9PEYJAe2RLbA4biVAPemDZRyu73UcRCmRSaiy27lVI9aV+bpjr+P/2WH
qEbk7Gf6LZUrQ6DiiTgkKfkgJk4DJpR5m6FBU7HTM+M0IH8hpZdRpxp9zErQWwcPq2N+4FsCluVU
CfYX7/lGZizLI+zGXzRyFJ0SKTOlSkKbkuSOjv5AktaxP4do7i/a1GrSFbXpt6OVm8C4vjnGku+h
H7nMHElaW9HDQcyWtrfe03Gsh5J+BtRDNJHVQjGWm5PC/upDEMiXzfPoKV2XEsf8kqNq5+s2+xtB
ePg43xo570FNnYrQb9SfvXM/cGIvLibx/2e3eyTDka4gjjo/60gS+Smzs19aUIZpF5hdNaTRtq6J
c7qK7Zw1Cb/X37jNgyl/DwsdDt+FulChW0ynN9RHef8rE8SS1a0yRa+bH/mJ7MqI2Uuf9ZRMEsox
zdTbqRQ3XQpLSx8s4ddrRX3VbgrREGAWCzcVQtDZ6IVNRrKPik5KDl0wDLnfgai0mZThQ54lLb4a
lfVkPnOkQ9MG1+Y9E1LInCzQa741DG8n2yewF/vfncRzJtzuRr93pWCp+JIlr73sIN7nIPcItoTU
noga/kebpsEwcHtsoDo0DNySn8uEIBHHKtLvOVuUxezDTNSG143wOSMg6ayMvJGEs/Wq0nuJLh2m
5Us+ePciVmBzoQwKPOGHvzrmQOqatRoK7fJwLbDlx1qUDf/fB8q6/wOgcRXI+klOobreI4mlrleL
qeplshLlLQVBk3P4O2bJ7Cq9oLyGTyvCSIulmTbSCSlwS35eTId8Kdm5gz8Li5vNK1WG51OQrY/F
GF2q7BoSFlvgBywmHWUvuQHzEiehTY+EbH1ggvkbLnWY2AOi0IDUwNu/o5X75UCSm9HrdQEBGbdK
ZYocCEiNJDFTWKAiHPmysbiMy99CvQ2UWYRbf+fhqYcJGI7i9+gKreAJZ7AuKAs2ZfB2vRc29ZmY
xkIPb8pONV4EB12M0eo3fGCoZbCvj1AJVkv7OoI2A7qu5hwYweiMTcvjN/N+DDdZL9IOSpRn+7a9
tdRlCPQ5jfwGzSlwGtQvtICMPaV0f2851qoAxytJ/7vFTdofzcek0x/1CAYq8lh/PZuV4L4Vk2Ds
EfpAFIeiTBLlN2S4aoca3BEDU+EmxzSXo011e3JS9ufXFY2N8tLBIl80k75T1aM0ROlzLNVHT7rl
PRCtKU7tmnvmIyJ6SdaHMPp9C/JNTV+fpApZWYDNsSIftjyQIQG0T72WAKZ6WYuRm0sbaHZ9rWXN
xjWrlHG3FRvdtJM1vNXDYV+4mMuUsbJLJRoGDsDAD2FQZd1qJEZc9ESR0qquUIctsmdP+hkmETJU
fxFNn9xUFxEazg3dX1tH3gR2eVF231zVKaKww9Bl8mTPNUzyc8ebE6FJrx9iZ+KTnsWXcJr5Yt6/
NVTqkTjmSFSAVnMP73XG2uiS3LJAermOfKFzZfOKk2dxIqc4NGaFc1QlvemQIfmYE0i3H4KE9NWt
jnK1sj6uWsnmt0oI2AivKKDprCxBBQKl5c+SLeQHqTPBTBOiaR21sjaxyuKDmux1XhCzFc07hKyW
3lSpP5z8H8ljNohgZwYxj93gGvaW+dgjGEwuCRuYRSkKBRkKlOzorrFwyW2DV3yHn0O0J8l18x/d
6veACCnmCaJFa/eYrLSSgx9aE33kVOp10lnLEhelJEXqdXOhKpG7pNNdVyn4G3ze0w0NQScsGbpt
fkCoY05ujTd1NxZh2CXpk3mxoL3XIj/ZlbidtGfbBHUMjIyducMD2W783svb2whzvXYKEYqB+9G5
hSsKXpkvckmXvv9tr9i0JWVeTvIyHw1XbTyv9AKPmPCI1isKifCpaRnq78NUhY53t9edggPFARgY
Me/vYwq2Sj7ROzp/DEJ3RzT6UMcqQs2p0a7ygga+6ZDxgFuk49KcsTZyhptGUcztjBijEwfuufm3
2rnwM1H7I49N2YJTsPpHtXmPZKalKl3I4ZERZxwef3ZQdEFOOPfNYAyJQB2j43U4JHk/zn50CXjb
0GKfRVcAqMdJw6ft2vUpFJ46/R2LlN5DNVk0XNBSMC+fq/YNaQM88cn3Gj2JtNtckJMUFiHGD57n
F8p04RooDgJle3dsLeo79Rlsj4q65XherHqZ7aYsL9pQUxH0jnUb2ngGAhbaxEx0bbr1gNh19eET
2VUStgFW+Rt6c3RdJmNVHckohTgzrV9qnRx95zSESWrzM6ve4VlwG1uX6ccWR1delC2uuCqtFBnd
+RHUNWSpfxyMf8ohD4dahhO42EqPzt2V8OvOnsP43M0bDA/DGNpxBwCXFsMPoz+WmFl7GfYmhCwG
w5OfNQoDp29etGqYASMPuB8W7TCkk+ak4Hjt8gUqSfRnUlvjtasoqfrxHEt22z+kGW5jfE7Ba5bW
rhu5Fd/kjFlGBV9s6T/pE7Ld54u/RSM+mGA1cCdRLBnwZlD+q4gYtohuJVV27XLV1QrVcpDkuLW9
AyiZooPR0M7TLSJeXk+7XKk7tzCiTImLC8JMvvlz2kNd1KO4FVtESw7BV+DCH1NWx6xvCfZO+gi4
Jz05ccDB5tV4tic59ghy2t5sxr9YRUameJ+JujGH6Bd0p8+cS53Ltgv+3drNp+U5yVsyRtKoE8lf
SKHsDLheakrO0R1Nz5ZhdwhUWeuwMiuLUexNMK2BdDctZcAUmyHw/t7AvLx69zlGfbXSEFzfHQcC
H8ITxM8AI4MLvH6jwK3PZKLx9PKv5IkPQ/hm3XXko958kGUx9EFzDJ+l7U8zI29b8MXVARbF31y1
ysvpsNHfFA2Nwu77XES4NOyAzs6enqnkKiniW4JiAzaSmYmEfHgWp9dNwFGjq9CTVBvVtVcB/HxS
KqSVcJ1iUXwECMzUFeHBp8vghX8B4AOlK2WePu8rrXcR7FIazcMrqkN3RkxjNhwd/3XL3WWGg+mx
jd2P8/W0GV4ITvGVFP1K+KCqie36GhwVDlRTb9MEuCZUJoQ4Ogtz4c22efkZH3SpRxEvIJiMPCf6
Iemc9rEmKCyd35mq/7eIaLFl5HqAZ+E2EWyAsiu+i4jk9dbawOpR4p2vQI0ORlGJuTK3hfQviePe
uQzfIvPSEGVuyZrsaD5mlXP082cA1BcdEHv5Rseo9cvIvcBflkiEu0UHxHq/2HX+jxDTNXxSQQ2L
HEAxvyzc2XqTS8JO5PugbPx0c0mC+AxPZfRsaDJ/ahjGv7Faz/MUapqLuLoyFQNmABzlzM1NoUgI
NGjoka9g6bbPnt4z/FbRUcQ+t5tuo9mZPH87vWrFBS8cysp/w72bxOuTth+p0zJLMyNRF3mr+ZQ/
MT6A0BtdKa15nc/uyOAYxPGzn8IU2PncTAsJ1mjV87zuBlY8TZHcxWjhNaGrV7DTnULXHDiFWbJN
sc+IRdL7cj5fkHb9bCwuovjjTsDFebsh4NiMJGlaRrW4k1Kr7jYuGm594IGk1EIAQpXOv1wZTyPp
As8ZNZRGzJ8vca7yuGyXWasdZPZNQu+RXHLzJmTHbcsMUPT1J9Zt40qWEXpo7yK4PU1VZ3MnC+66
7afBNh5oLLcAvEy6hwkoSG9CG9mNkKE0hElqashY9lImCPbXPkBQNp96fSs0oZmXduVTDtP+IocX
epthwg1MsjjYX5ZvakFnobn3oJxxuiigkqJV6myvDtF5iXkxpbAsu+iJBRtQWWcaQvlRIbJtGj+N
veocvlP5AZctttmhsFzH7dlD77VbOcb3v/HiiVqbaUOvQRKrkZyHHqZkcidlFPhxiCtFEgtjIbnI
23mWJDmEWp1BhfmwdbtOxyd3TNYbe+PBTGL5JdZi42OBpah1cuaeB1721ugQCZ0q05agLPA8UkDm
l8GVSMBubGOp86pOZ/04MYEthfkfaipKCTezrT0O4LR06nqIpkCaGTrDwRUd239s+0gWnn4k5T4/
JvlHdfUrXUGJq0myisIumx/baB8KClrzIne6fVtPKgPdAQ6Fyn7l7nhpotQooV7NMoLUtPjnYCb9
7TaG9iru5IksvsO1KyAwg/xIp7hLscQtP71sgD3cx7WcBl4Et80qwexxBvWSvGUHKIuXjOszGq0q
9OYCR3fQVKQ3LnVuwJZN9imoO/tbCASJTpKOq5fB+Z9Qb5FmU/Rrsz+U7ViRix4B1nbO3+VMQ4OA
Fp99hWy47rE83/wb3sT9koN1vZkvY/pH6ZX3G2OnUQFFYBNphvlMdTZopG6oByheD2qWlfXfOaF4
1LMZjfLt2hyGLJrDAKzrGXa1cFN2rOdcXy5xp9zRDE2LD8AthQTbwTZuImtlj8Zd3q2yeW1PgpL2
8jY+3rJmfiGfwaHZrDmQMU0q9a+uILuemzIiS1wQ4hjudXAXlqKFeEIFUetT4/d/vOxoSX8EPW1j
OTR7bVf1aWKDvc1yB4QNGjYq54whX8Dw7sVLsNF0d/X+mgMSA6faAs+dSgxrYClGWPaoOQx6Z4o0
2HsEtujl6flxjasYBeO1hMEBcszYRcZMxTMPyY/xuWQTEm+9WXL/WSIw03g1y3YcdfaI551HXsNp
GF4IHQniSJHLYQHtQxjcZ+gPJUO5BybNPiWSmUWFPcjHMtKPmLw2uivDkDA7B9ro1INpKkYAu0jX
sroSTK36+fH4mJnh38RkqjuH48Qm1fvGmLJBUxYWt7cBjbEf3QgNbG9VDaTfhd2Dwo3VaKKV0iN8
zX+3P01DRK0pBRrrJShg3yurUPNhiKIQt9fjnKEwB1gppFLyS+Uaba+4A7xyhsYHdAtCOtfooOXr
R1tHX9Jp0WkIuHwB8shDCjpIANpZNly13RZCVVdqFsyb5AQvc0h/6GQLa90qDHqhZ5oQlmfECjjD
c8BkHuEOGRLa4hZA/myDxtEgogEILt29txJyVDtF/p10dzb+y0SFr9xtjERwRVYYmByHZ5C34ptF
CUBD1adkgtkGNxt1Vfd899r0SF4BaBm2OyuARI4zTzFFPld59RTqtwEnPBKcnuJn9Bqw6LUKq9Wq
t5VwWmnh/XVpElkTKzTKykrKs0CG1Hznh5z12iVxsgPmdo/SzepNrf9x0gs/+ueCNXpwtrIPW0Gi
5cvse+q/F4pzmXEx20dqElHf5PXktuWwN0l9w3bXntmk60aD3MWnGubisRO7Yzbh+frra5VqynbQ
/mQbHVBPjhpsoyQS2k+LAW2TjyIUNwxc5xyCE639XfxxXALDlHC7XpUkUFYbuZP4ph2au50uQxa0
c7ygQk6slyNuiqsGQYrMd+fgOgX/Ye6yGpbgsL/dxYxf7Zc765YCr3a0/zBasRy+4mbXT6HG2XhU
InebXKtNoEzF1+kLEKl7kV1iM2FXeCvW/1dyPAeo3+Z6AzP/mUAUqx0e2xt2aectVlT4ijAF4yxY
XHM2mZmiigKoNLceT18r0qi3YMF2monTwvk5nKOqhQ59KN2HtQIqgldEVparN12rEuTHxbjQA1lu
bg09k9yAtDSDcJNM55cCfZT8mltnVApNDOCDKGFXnZizVFYDBzI1XJXs8eQMtMn7AE9MlsyVu8do
fl5Jta4qU+XwhVHum84gp4VGGxjpub8x//0u8mNpUEShQh/3WK4fmVvlPey/nNsU8TMAa85ZQt6a
OMGJB3u5oEHCxuwk4QXfyVnCzouQJcsROBVx0CMv5RXYeP5Jf22qgm7/PpxktSfgOXuoBhVa+3AM
nMVtAxkDJS1B4pRrhRDoz4imWiJxnv86ZVnB0eYsmZa4l6dcMZHnEEUqSb8w4CTezcI2bEKPEwpq
Cekr4ljv9/3+ugzJmQD6T1LqFQ6JFX3yQ53yIangPm0Tt1sQyP/Blh1xFGJmZ+OtAq+1dZPvmIxw
fyDljz+EE3cs9/SQ0B4wuJp9hYmoRuIMh2HUmTJuKuVChfP1P2WV4elvALcR5lwz3T99lGKR1rtY
yOoQByklt3M1F2gZnXva2OFkd2xS3XVyHj5KnuXphetdLLaGT40ICjCSPOif0MbORkGTDSzNayK4
pPS3N8KVn56l3EAXsTPXpvoC5sSZ+tbq30RNBF0gngPsHY3qJOLOUQ+iIr8AE5pBWyhhDTFufdDc
8I664G7x3hd6XS3C5jNVSZi2mgUT4agQG6Zoh9HE8pqksuivFrOLespfyH11iKglDjg44anY6QwE
UW6m9EKWVN7iOiXJduYBsTX4+HinngouyoUrwMz9ySaawQ3bvas7R6J0O343RflEgQZijrBegord
MIgOX6nq8XurWOBICKYURul/Tt0qhIMAH+hp7XVmJxRCMATyJsHZRSpGYqNJnnyPI1Db1JeXQ35x
5zWE4VXaOnIzk8mlupdy6QzfuUp5D0gTj3Il1ctjabBWip9XReNWjuVFMHaSZ+XyciTSNeKMqWH1
ujGGH1Fy8mLqvRKDxhfRbXZaFrmmQtp7s2xWDpZD/pJ1Oz41bNTeXG6yWwMpMquq4rvEsQbfa9df
gR6wdyEpvzuIdMsFPAUBz3z4XggtgUdWaNxnygG38OjPkxue77Fil8uu13RE1n35YGFuxm7SE4O+
UVG4eo5w3cYj++GL0VWtN6Wdsim4Bx51inIiFWe2IQdarPVmLQoBe9B2G3dx2BcJgII1tkAlwvB1
Q/+EHi5S4GjH7YpM+y1Md5w2v6MbIvWX/QGHuVHNSBTNAMVHTZrz5m5WKTDu6GJhDz2TQNIQvYbM
kQsmVCrGt0AXl98/s/VkNQu1rGTVqXEKPU1OTtPXCDutGBnGhmiKqQPRM3/2YgP6A6jNmX1gh2fX
BzhkWaeSGAOoJzHk/nP47d4C/FiflWLwOtL7pVa8EmWSJxfjK/ehxjMCkmgzPQ7JoxjYw8lOARZN
gI/eSQSBVGp5D1JNvtyfLlhRCZPdvHff4rmAyHnQkoTjkKPt7TUCcRFENcMRT1j0ygBQRaS9J8L1
WOgwzzQgvES8zkTz/G27cAo34am0SE5Tfnr1JmqAe8nPSbOrgaRrdggkgtUSUDprjNs6VS5e4DbC
5TszoPJT9SN+sF+3FbnZegIR7LikVO5Led8FVjxAD4rzziwxsRb09fGQa+EjGo2tBjln7bpKBeOx
fBrSS7msba/vWPGSqKZwzNIPqVR2pL9P8Qmu9cDluN2H7tLQYHHRXGSKUrfkPnahYkiZOWXR49X0
l4He8CitKmRvYsGKl372d1NmUPGKTe4Q/8HHqaFPFroEj2uCYMFUPt7ARxvRdzpsPANS6nJ+xMm1
RzR1y8BWymhLPqqVYPKucWYIxl4BmixqsydnHdy1izKWLIU57Wr0I+BJPKQXlA/dIEdtlEZEW9Mu
G/gadwyqWFKPuiG9najpORY4Ym9rvXAzFj8XzMWWNs1VaGRqPwoVQ/DcAehUy/wJWy/14U6rnY5y
wJXm1MMRe1cmb42AV4HS2ZoezwMFhJJwob8TnV9Alkif+edh3gvkL4Pcb1ne7skrq+BEtSYdFNu9
kfZD2jsbLhDMUZXqJ4JIAbLSvwKbzhNn0nubgnq1hwB6+Jvi6uHNrpYkMXXFmfGntd3dquw6hfOQ
O3B1UbdDR5OYMfJdhvEx2vsj0/RfCBRtgkIi7KyonlCmG19PhUrBJ633MrNArlqKSQvri9asyliM
MMoDy9og5pxHUDTgPWEoRFoTo/p9O1WpBmYEOKdkUzba7NartqbVZbcqJYMLIu5258qofEEgcUqH
+R6umCAPemJFT9TWYF1BsgTVcegSLUniB04IuFjBmQnLlN4TrwFn7+nVw2tUAD97X+PVTTJHs0IO
qBh+Al75wVJejMMEm9BBUzL/9ku4Dt9d5wTjiWeROBXC1YC5LMnQqXWLQWXXIwOvqTsYjMa1Ykkq
J4AEndwtOHlpOkMftGHincA0Xc6Ay74Rm31fMKa2VU96Nj4ToDrkTrieVsjxjIPiPKVClWo7nCul
TckInd5bv0+icO1hPLeuLjXXi/TKK8xnsmXyU5xNEwnhzgFRRW+hMLK25oxpezSFExDBx0mNITqm
pQMucopqw7Da+4dtEAmVLPKTZzkKCZJXLWCce+EeWF0wCDQM9m5FqfzyBAhLpDwoGGmnKUmeYu8x
zfsn+MYDho1+Qnj4fWUup42SUsaTB7zRYKSOnuUvKpr+9iaWksf85OHaJiw9szeSjnn2sEe74U18
lmQz7f/JIfw62DeDhVXZjYVzjOs62vy7pLzLXvoucrcEINolUDa5vpncHA4fym2PhO0ss5TbU3CI
mAV1Bu4UiC2J2L6cwQRduEgUyu46R907PQ+Z9reisgB6Ej9CcybFJp6Fhvk4e00Xue9rY8aCoBpN
vDk49V99Ze7u7nhVVlANxmnSedc+bnhYoJCsuWQ4+5oWHMJKzZSKN+j87nVludaHwbs3lIN+TrpH
Gm8ZKFyXMcF3U0+t6wsowXzRGMYJwJzFBe4KsWV69lQGVA/vaWRI8FJIHPoboFT4M/bLSBgP21Pk
QPxOv+FD8JH5m96h9rxffCJT/25lsL0qajw0kGoVTvY0GDCV+cPlpdK1MrhLTbmi5IIwDL9Q6BcG
kmZuQf482Ev8lTbZxdArSo5YLw/uJRwL1+kVGa7e15cgvVB7lb3NVJbUCg/Cs8FBjAoZmB4P2s9T
Hm2hSmJgNSzSPWauGEGw9A/UdBQw7aFEeVaxCJaAGC7EdFiHidX2aRPNN4O3JCaWlX5vBs3p8iTZ
Hmw7gxt+Q4edvK9ToJCYggTG1/A9aXvJ5hpIwK9e1Ksitej5GNpvnOdal1sh/Q7/w2GhzQX3lDS8
uTMmIya9H1NUrYtK46hZ67hTBTKxFnFTiKoUvUZ2B2+SYNndmhYB9UNg9/HN6geB0kRiql2RbAwK
OiWC6Wchd04pPoCbqIk0AyJEZge9UZho0Bxzggw7SSG1obMuTMhWh/KS3D77yyyyRtj7x71r3jQL
Gb2XVHAN++eKeOz426KTx/XXcQMHTQ74TMEDcdu4/KmqDFtuy/2AnHRUi6whT0IZZkiaPsulBmHg
MvALiUFxqAkRwqtsELhrgFg0XVo4CKZHBZzWUKhHAfcDnUPxGxo88nut5qZCbkezcr5CRvjU+pt4
aIGaI+obwBWpm6moFT4QZE+1GA86A/QZCJu2KZeI2uqP1L61f7cV81s34DovW/UC9xDwZ+4pA4os
ec9l4/FTcNB/+rPxFd+2Vr2B13vQOenIpFXfrB/fd+hsnKRQXWTsNJsmYVMvxe+JlTNYDOrKowPX
Yk1Ay0KvTAYXX4z62L5mu+yaEi6ItTsx4DmIaI0JYQZvMvErv3IiQ6U12SUQ2WIfYE1pSAOFbZY9
L1XZfxXP0f7ZtQcvUqbhxopljiY1DuJGBuUTHRAQRb7vfgCP+CTlLSIH23/z+JtM7rKpfstwPWzf
2fDijgVGQL58B8V/YcxT61Q3CcDFYMCaQbWsd7/gM4ZO2sD6sy8k5lQSWPfXpgoEqhVOhmr5+6dm
XSHncNJIE7Yas9JYHBbaMewjTv7IekNlOUh4gaw0mFUH7Ki4ZwEZ5FpelnB2Mf743c8gi73Yl/xt
q7z3C1x9VGojQdvU1ylJNnRTX/ZL7xFl2RdYMmsTFvmhG7q4pG0AjabdozpJF5fnMa6p9/3t4CS9
JwLrKNWfsdv7BdoZ97kmP8uYeormnOZRt/DW9D7SYqsYP9T/203d898zgs5WKJk1FshP2LiqwGwL
vXBt2UuQlazqlSpTVt0xWJAt1kue6I1b1A0K65j1lq4U4Sgq2EczeYvjSXJ6duBFRtP7cFDhOs0L
pU/VYEdKprpovZYrV2SsGphViDfsgL6L7r90VeZjnJmqnZm9+TOvK5LsKzAaBkU0jviwRks6B5S3
rOuAKz2XFwsvvIkWo3NM/au388spJgl8evqNRlXb53KmRzCK5zdppfc8tM822BIu5UHCBymW/oqD
hHQNsAW9BQjHV3KFI+fNfxDCNaIXPwRFVbEGb9JQfQmj5sZilL9DkLBldEU/+iqRqQSjGqwRO9+I
dK1Typ9NT2J81HFtmEGD+IvNWgqlRZi1fLZ8rW9LjKhIp7iV2VjIwIVOOB3h5gMBUiMsRKvPJuhU
R1YqLQNldv2ooPI+X8zUswX77wpK2xa8UaeGbYS2D29acEX/NL5GFt8tFQBAKu779YDbH4/LTZmc
Dx24JR385jhvUWEHnIrcE60cxd5TEUZxD5xZNkqzIiffm67sPY35GDXr0hQWrVt1AH7h5LvZ5rpn
JBm5cr9wSwZT/EbnrN+bG3QFI4PGGmNxjvpp6+RGRZ4BleVY5DjR/gnokYk4DWV6ryRLzPXomJfH
ALWxCJ6Y3ObWV5+rtoC1tAZ3ZfWOZhB/ffwmLXfon6xJKDD6FwnHmaTd59y/NEMPiEDYo+18Mmmu
C++fziUHjZoCXJHf1iUhVhxW+eeYKn6FGzKmNU2ayAioWXEQAWyrxah6zKEVKoSf7TocsH7JZqui
1jnucx2iOTEk3fFnv71pKavLedPC5/x65+wSpVq6r9R1IoovCF+ewNDrVgzyRYP+nSOj6TcZO3zZ
u3+HJmj7yUuM2oV5qbBdtdzqvWA5z72NB/yKNCoegzNdl/BQimY7BaA8bS6teLqwyvrGnIbCY1Fq
QZ7JZ0JtptMU/vUtyl+doilhHZRZXBFqdAFRajr4ojRoO5a9VnLZCovBUOuT5IDIXybyx6cLh/RB
VCHCyNSlResYI5C5Ked99ae3mGL5i/SxkJe1BoOhW0XD/sNzZiYtQFQNpKxARLUb3607QedqpiqV
RNbwrd4sCv5wMX9Wn9dIQIJfA1vbB2GGOsqcKzYbERvDGL9/Wdbre77mcRbRYKxarlcpNE5L/mWH
Qf0s/dkipEu6tQ2C0BzthCx+RLlWJUmZFlBQCwg2sbJ87bAtVqPjDBCFB/Jg0oHCcV4Oom4w0l2B
ODgJgnfy5NikFQnAIhMqmNX4lAveVuvH3skiwVoCWx0RC/DUOR70LIncVPbmg67bmmY9iE7qi+OQ
RSn94L6nFDqpbBdyWlWe1zlVGtw1kC8AxGhc+8dl8JwF8C0tzk+ofD6b6G/gMVkJxS/fqVDC5cE6
EQEOYGOqk1IrZfn+wUHbSl8HvTjxACzHjMfzzJXfmhKv76YeQRvytoz7eMFI93iYDJCOCtwqH5nY
+FKj+vdqk+VxEu2GECsLGqnfWfswvRDYjLN5vmBzd8WO0KfQBX+oSpx61++qLOtSdkAvKAW82VkG
OsEoLZLtPRrj5OVxnGmkq7pXPq/D2wQTLZsqcAHy6VBfZyyNaopYwY6zptEjM4g3vzytjMlrtIPI
+Z/wJ8c8JSmnIrUv7FXxs0SM3mxD56JjkkxtShu7Ev/OwqD+CC1f4fXOrTeItX9228h3BaI3ETgE
dBlEEbsd27U1mVPxPMyoxVn5FeT6P/NJm+0DP1hsFie09xFbduCGS4G6y1he3z+EP/g+frB9RG8l
JL59lz+HBlWELYlZ9cPXQkdQ/dexwBzZqRdZ0Qhqf6pQAUpgJd5dsT8WKZrCSQSj6qr4ozg3aESc
LzDqHxQY/eKeiG2nJ7h7/TauJsUE9Gd2uo/bb0rtGUj+O4crvoBoOvSs0iz2/zfBCGSIvDIpY7l5
QGHqEET7UyOUtBaYOwRyrfMWIxm03JS6c0sHWbzOEPmztL/++3Fq2nf1WaEZq2R9wpN8oOMsv259
g3j8uORCLwVSMjAJaNTmvc/6FFDYp8ePAxWzxWGrKV0LFiYITKgysRvDSziVLoWErlU5mVh/t9Er
nmxh+5oTAuXXEjqXEO5c5PbntFjFI9Rriu6gQVZhd6zXm+UUb8YvIP9pU0nQh1jaNLMkwpcCMj6C
IFpjMUqD/NqCxdGY1hWEj08ksZA0YhN2J5Lq858n835pniRXt/IjbZsO8GrSCQ/ukVrDfuW/PMiS
wwG0qT1kwa93mud/qDwFBvtp8R3cdiXwgo3BPtTcc0JP5BxYSMQFTEVbg9bD13hWnQqg8Dbt+JJG
SMLoAFektc4HjbBCzKlPG7u2GmChWEQ+3DXY23oDR9wPSCT3qR1geFBbpRbt3By/PIiqEOt6C4pa
fkRJMUohU/U85DF+FMuIyiMjB/mV5qz6MFKFAkwyzkAopn3Zir3/NVlqOTSWiFh3VMJ4xL6w/snC
wCFNODQvSnCrWm9BvEmmtDl9RrSL2wmT3jSalUA7LCg90AY8fT9vnU/MoNO4rjiU8yZtWBrKUs75
ej8TOqSwDfiVLyDZmT5B7zMsy5R12DvLT0WWrOBSXB5qBHT5lARD2vNPEOetHEQYqlLlWydPhQ5j
Lwj1zc1qs3xEzZFwfJtr5SKcyvHBd63ZG8uDyFYaMywf1AQF7bxmWx4a8bBUieIhpwGRDaMW0qFQ
QiwYKoemmdWWRqSlcUeb89NNogtpnPEDG9zUQQTsKEc0wWt79xQvC5KqkXoZEJMRm3HOJu7ggkHp
atQaWOb5IExpfkUYihlA+8N9/CeFgDsVVT6sSj4n+pHGiTL7D2kE8QlPtBItcnAdzL8w3KVYffCD
tHXIv6T5zBgwyIqsr5YPIpKYX8DPZgsQ1eHEfCggQA+DvPELPv5/tp8wo5k6mzkKQlt7nuuBgphB
O9Gz0RIimIICSN4HyP3t2IUTmW/Epnnj5GG+i88a1kvVwC1X3inrSQOGjvnvxrdUnP5aPivEciSI
TTilBmoGl/j5D9GhgjEGXrYopekQ58SRPgFo2Wo8Yx8qMu5cBgZD3oHzWG5ps9OzfEj3OCV4dcrv
so8S4E0yIrKkqo/xk0wKpzrou6n2ch3IEcahZqTPserP5RYqU2q6WrAkMfwEows9r99iWdEdoJ4W
WI1eMXE/aFZ8ZHX8pvuj2ldmziguyj2U9a1QgzLQqH9LWnOUcS8pclLNetUEa2TE7Eucoxoy2UAA
22uVPMQHqJUdOuApFfKxKgrStIpX+env+3Iv7ubh884x98Ps14pKqiSIc9Ney1gpHGvKaNAAiVG5
WA/WnK2KcxdX+GnJiMwnJ0Xg2d3rubPdVnq84lVBp25dsDHsxYZEvsXw++SlsZYxQJ/OLfHB3w3I
92vlRifn4U1eh9AIIxrHWMKl31MNVDL/y1aLWNR7xeHyiLxXNr2LNXIBYDfhaYXKQ0pcYQuPi+3m
EeqWxfir6AH/qHk7XEpNXwg0QKlhUjeEcWR2cRsKaa49MsRsbFTBRJnE/yiiSFW0JkHt5xxVNH8s
guRID/gW60JrnFJLzddEXY3bdjavsFENUmBjf8BwOaKTES1QZMkw1DGWwy2/wkMnaT2eEwFm2UhB
5HMILg05qL8wnwDOE9Qvk108lZoJ7nSU/KclzNKXxsNGuN7tXcMLM28YB7kX47sEPpnMXx7L/YHF
qfGYKyrWsdzxK97NOAhXkABtjIYz3eE2unGiYzq04pYH5Z8u6KNr6r5Wnjv5Hk5KqT8lcfZVqs94
ypOiContHQ6sQ7Td4bvZA10T5SXlKWH5U5z1V+IE4OYSAyXnGUUpW1q8S3StD0jQY3ValF4ZhO7c
cgeNmuSlg2XanLkN0UeqnN+YGRRz7ZvfiyAQl/8E2/d0ef59XindCCkjy2nKyqNurTPk2LSEMRzy
L5gPeKESy564pQ8M5CZbxISuf7ul6QYczTCG5AwJNbMOsurd8C2sF63MUfmhfKk7Q5NOM3SJFLw/
0HfLqC+U7G/0lP2PlrFFVZdgZOQbD92jpCwitnmw9GE1tLra6RX1ORB+HJTNRsE7PgJA65fN8TUE
WQXOypbqVG3AmvRRnQUe2YcgVsNPZInMr7YkOg6J1Sq1rsP7L3i+3cjrJcYdK5ZGi9t8lhrcMid+
nj2kIdPJChEhRuOjpVk44oKhrlaM0Jtw3WHrteL0NF8YytWUmd8R28+8hhKyJ5yNZJGOgW73qlVa
1tI2tqLz3dMEfgK+w7QbP9BTgwztmNxhNnJGkIfHCa/sEmG92MunWzl1U99Ef3h8AM3jzJ0ny8jf
LhW2oXrZI9TP73pZZhL7ex6i+h53FU/Ne4ih8zxwilKTkpee666q3F1dqkcAYAAcgVPfp4wEbNXR
5POA+TsEaEbrZd4JzAxojjLINLQ2KFZPrqfQhboj4uV2KfBGm1EsDQPSCrGE7srqcBd2J7J/jRkD
MjM/+xZ4SfCCzraM+6FqsLXb5+0GhgTUrypMgy9/qmJfPzHBD5LqOzCCnvHOVyytz7O9XGizKsPS
y29PiIshbjjeZ2VQS/0nQ7sNpyq6GtHcgu9juE+M4CAv53VAcnsUKYRtB9o2KEufXs0gTLRxqDmT
84eqpuOMhRzkSIBaQ8VwPXW6XHYP7u3p9CfqAXhQFuVWpvUByNn94uWXQK9wESwGhbvzsprPpL7i
z5DRdF8eggxZ2JwWIWCbREiWkOK4oS0F0DZMVeWmqhmeBzOo6iKUdMBt6AEL0sCgc1f5FpdByKC5
jaTaL7ovVNEhgwt1paIqFinWoEXK988aQtj0XO2Nvrfuz621m21H6Fb1g00IYvp18Be/GOwqJYz0
WWJMC3BTXj+WHlNB0CdcPlq0Az3CwjcOR/A0wZ+eGNFzYy62APweek1+aTDaB2bC35yHNN4Ex2Ev
0abEpHrKRcGdfyTbbBt8fRysaIDUljwFoNbQv6IfBRddu/9jQzp/YDB/p6ePbw1CpF2GDV5JP3zp
eIK3uI1TosqERagHhi4SVYRUd9NEt7miGN5n1E+nQq3nlIrIuhLyP4T200QFxMHP0B5jfR+on9K1
kis2qPD/Vs7ZTj5reqyI0dj1L7tK9/pzEszIKOw89FTD4NjR0ThHmVms7/WFkJ3VDwQA1iPqiUk7
3lngGSYRIUvaQQfTwc5RrR2VOa9BEAoNdeD64uboASZwOUdvuKZzyiA/7RUj9BeY32Lj7Y9f4iZH
QGFVwbh1zujJYzdR3rMapIjYCaR4/j+rEO8c70J0Gt65qSl2Ffp/l4ipwfL+ENgo5twD4chNdpd+
O47uWtJWvhaS1HiKi2NzsrS1W1GZfHgxniJP2UDliqxMu5RZnTlz/llaIdrDDJZ6UtpPHgY40aI9
029qkdIstW5preF3CnX6MzdlaAAlHnvsGpTR11JhQWclzbEuVSzAkERyFUIjPQybIX3QXXkaMAg0
QqJ5bjUBJcSCWIUpLyuBSD5JCl3XX04Q2cOqTLVLoNMybjKkGMXVT76zEOdOp5agp/cD2CecENgE
wBnuFDKGv5GZVREUUNQwubyiWegW3JI3fxgVGRzKzKLfPBUZ9Yq122a1NSbZylZoktdmdETS1Ki1
sIRvIMXAqwQiOpIWoK/oXcchbOuGltNYWX3+n2MAtShJYtp8VQol4+M7QSB5nOpco7RGbXKVHjqp
L30yx7M8UIq73vgFZVm3um0+HfnhSFXXbCU1shuKePKEsiJxWQIBCv8lA9vmJB9J/LufhQ96EIk5
bKYhIrdwv4LsXr9YHMrWYJhL0zwB0zPr5/Yj1F/sREeq+bhJFYHwoYCOsuz9arp6b4hQOTJ65pyp
nECtBWHSlqH5YDSzpMFXlapvmIr7fLH6gM3vIq4XL0nn6MnEFQu4STMLTvMxBlVnbe2Hd3MrkFwc
LjRj5UZYCXFychgDipH2HfzvRqzPCjE2LD8bYT+s65DWXxEP7X01f6Eaq+zPb/GvCHnFgWl0jDU4
cXqC0uPNgs0yRiHSBIt3vAdUdXhyY8ywAdP4KkW7x3OJaFfE6Cgxgowwp7znyOY6Ai/ZWD8mvfLc
/OhpKJrL3UczMeiRUowl0pX+YCdJ3q28MJGvw06+HiGiDtHGYZ8XcAQYig2HjOoDfWOlxtRLdhS3
YXwQp0n9CPltOYgvTIASRm4FpopuCu2J59aDkNZK7GQK/1K12cGTR8inPmx4IzlAWJIf85b0i88y
n5VSZU4gntCElixolTDvGfIHtmgjR5BeGU7cV0vVKFOYI4WlWboCBWFbQAg3nMo8cqANDMtnXF9c
fDLoGgmqemTH3imwLkzar4s4gGwYRNwkKAg1AZ9bd7RPhfpLPZa5kx1QKh9896Bm3w+8g/x6vKy1
vWcjxWJgt6d4siFD0pwCkxWrqqC/mqgSgNVPZYQ0NaXhISB+pIS5OiAI+7vcrhCvV9c3HbaHqx+L
qaVaj0OFHKWfBZxYxE0MZJ4onW4OmjcZiKXknuyN6eq98RnqYDQQ+ho77UBpBU4f1+t08ZyuVwgR
UPEEFDg2yuQz6ECEkdPylAKxJCFSHJy3J/a7eKS3dmfpYFQGBXGt8FkP1914ZIHh7sFw8eSNfajp
yvc4rfNTSuOmStlCK2DyqROXROGj41YCZg6uW5utaQ+FfNZkIqo7GfCS/4AOZxaAyjmJtdLVTlpH
lxc1W0PL/i9vC1FFUUhuFBwC+Gt3NUxQ5WV2quIpYMwFe/4Ker1Cf9AoDBq7hmcbv6ZjltXf1sp3
uonMISH1yhj3gAttRpLX2VxYx7wrXv0sKn+W47onqO4qELajLzyR4Qc/m1Gj4RU/7xnkQNxxZap9
n78k1YrkbVvqo4HXpTOFGwzP0cfKX1LNCDMun4rNfDU+d+g0dYA5OQhmnxrjr/H4irnm2aqOcNWu
27tiaDhJgUjsh9uDzVpdgMOH6pt8cyMTkuqrLiqZpu708lnO7/WTO9+QW3ijQeNUvvk9KPSL3O8p
mswdSaQHhH7NxM66jCEbviDqCJlouJjk/YI736vQiKzLYgCYMdhKQMf05OmbdV7Q+0m7PJcPrYLd
naaGpkPOrk4Q2ZNE98FYU2x7+JZu3NJBlRnwupk4SnTUUNzWsDFZcRLZVb+6sWQ4JrXw0qYhtQux
MfvVeQkllLnvjsL305johLhkwF46NO0daPFxT3/jgyMtpLpKlP0QsJPPT4hR6h0yWz7a/uDUn3AW
IG64pTfeGxNDJWYJWoGM2X0cjKFe0MLQOvb2hqcQNG0vKFsnhTNtibM8Hy29thQKQEslChoAzYGt
Fgmnm1nByZ7Sa/pUaTWbawc6q6RuR/7H2aZesRdPhK2vz1wdC4iY6GlaA1TqxBLQctCitF12i05F
AGGt3vJ+tpAHdlG4jD32XHaX70HbgovoIWJu/EC/bpKor6Unz+nglDuEz9KJFPjVuYKMdoFN2Xlk
zYJhxq9LeLx4Dz2d7LH/Fbys2sw24o7pHEh1yzZWaRiVwftowECtYxcgFagsECVAxLZCVeuyLRfq
wopDd496bOS+ZASp4AE3ZbPZngPZbRNO5jPBxAglJkDkYpbDC8MjVm6QlYaJagmOm+OFRj5CUIcV
TJLoVrP9HLLI1ee7YL0WZZ2ihm+D6f/PCo9jJpNKF3o3j14l/+OmPSXLDcxTKNBTbW3DABHSGvxa
gWcdQdtCYOdL5JR9/yec0YqW7RWvRnYe9FhHsj/7xNE4/d6PVMWOafXeiezKqpMy2FFHiKKDhWHO
l9MBAC+QI/DoCit1e6V26j6VbHow14MBlKxjKktUfIS73DNXE6Au9BntR2uZgUvGFq95dQ/jBJIp
vCtUFt5NAflazblwXTbsG6ETaLlaJ2sDwnhCQ70E+aycRTwCVl/mUdOobUo9P/7zgEBsTlRyL6jz
r+eQf9av0rkYOXzo4C4EzKs4r0sD171wLBkYzDu+at3PWFXG/fMvMyk6Zh9q9IHRCuVwGLvfaKZI
4GwN+h07Na8vXd0myiB6MWNY/2fVr846biI0+q7xLhLGxqZGE4gbO1Z0IrxYqrWxpUzRFU6FxQlT
4L/hCcuspPp1ez+xG/ZWZ9wRpzYp1l+HxA6DTKvSGbXPJPWItMqbqYJ2/0pVReJsZvB66/3c9Efd
N/bqpULWmOvY/gr6U1UPEi/hILZ7vGTr3J8lnmTV76yuljuiJN25AKOMgnMJn2qymn7lyGBW8vU2
5b6x2OwOnytasgC8aMOOGX944yyx/GsevBw1HjtFPK+KPE6+GJFbstFJq3KHLGVahv5jSF58+y+S
6V3uFZzrAepAjLSbRGNFJM5Pa3R65Vkg+sAHGTOJCo5cR/xkWpFToxAaY6J9Dell+7H/46W0LSs2
ADT/EA+3W6ttB1/G2+Y5iLCtyWS24V9ce29Ur01qDjHd+wBtpElMyzys2rgcnTbrwVv5RaU/wq5h
airqr73uYCspShnA9wtM1OrVFTQIsILtt1Nqeu2pCu8yWCF/w3ZwDIUxlKE4pRU2YJCeAn7PI378
ksUHivS2KPxL2OyVTIZ8kbv1tZR8kTUd5Ii8YKA1pv+LmbV2jJKmn+jmE1LAAIlESf2smdh0Tl2i
eTKpJpRuQeeMdxjdDFbhyDVVhCboMTXBNnF4qY8PpOIGz/M30ocIyPkr4V0PKqk5wZLF5rFQG9N6
E6bf4Keg+QOrMTwduZUtVyLAB6Lo79xg922g7+2yoG+gs90J8tN5dTVPuHtJp1xSX2YC0dDVrzxE
5Ngb9We8TFBKl9RNLGFYv0qS5a+TXYO8tqRjQCCzg0mF5GOt/IiuPaDLF4H6p6QbqqbcWzFeAKFF
1ipmc2Ko+FeYC+xbGQ3WB32U/0oKYiQhgWtyUnMm1StEkkKbR0TgCyicEqNJvJl+RFQCByA1+S8Y
FzNl1X6RCHgHF2J8cjRqQyzOY4vYRrxR6nf4YpwoB5N7oRfvOSwZY8i5RP82CK6OzPj2VV4iUB8N
sfKGx50XmsgIC2beMg3B1ZsL/Y1hhIaaauRdZ2dFmT4QSYFoFqWd9XaQDFxeK2C8L6DFAXNXPhQx
Y0mb/YAcHac75F0zRpLeP+dMDMspi2YIR3wbMCL+Ee/og15MkDVAbjzRuoxIQrVq0Dht+MbavE23
o95fN0g1Ze9pZVkigmqC0uXsutI1FH7kqvHPOVubxtqCff5cXwTPX5aY4st3PsMdV0Fh7FQ60Ttw
/8hpmM+ukRMO96RYZsoZhW9FIdLNltaqPvAAWsOkt8LUTkR+EdCYmLrZFaQP2sNZR1NqfKHeKRsJ
vXNfXpfsQCDOHGbe5+U1biDxwB8UPqAigs29IZyguTL1Z0uYbXMN5UZMbQW+amk2OsaQwMbpcCDa
Asmp/8DOvKFB0XyQ6NpaZyOCVAE23SXV47Rkriy+4qu5FQaJD0TEQXGMIWmqBBTy3VQJP3cJ1SJY
yQaNtUSUU1CSGLVgcYrAYB5/4j11sfZ+Xnhj9QfM40V7PL4lLr/19LuA7F78TiUBmil0Utjk31Mf
/ELyQ/Tk51Y+9CAKlgXnK7O3GB1YZkBEjRPlnyUONPYkU23ZOsmy5WE2hBy3HVZxjbo37lyaLgt1
4GOY1K/ApTQgTMfn/NkjGZ5OGgQxNZVdrQX8K0aHHOUbjnQJyOUaemJFzp1xqb6mEe2ZLecWE09M
43RsvUGJU2x15ryX3ZOi2/97lh8LCRoMn0JwJzmNgTcO6obM5+WgBDmSKjU2r5lMjyHI+TGpynBD
AbuHZwYFMVkuikUy5l1WIvbo3zBhzvlOr3/thdjDylEXlpL34PgdeyyjiRqespUZy0Lj08hU9efo
oGr1Vi5WytcEj9up6nHqcEEy/JTUoOOaZkWtxrbJkzuh/7CdXOmB+O57mWKNnXGgZO0J5vrEOqSe
gqHFcnroA4m+L4DySC6MCcz7ttVHF9E9jdV17aGwgaZd4TB0oNNLxnyb61BhO5keeGHBBROhlpEb
05BuUfST17zYne60ay2vrOuIcL/XJjwnmMkBcmCuzo5tGFVw/VHRS0KfRiJ06BtYYP3TKZ0nsy9R
MjlyCeiBqj8DIwEdtl0qt4K64h5612XKgqki8gtUCsEct2nU1+GV4t2cnVy3dAUvogfb3nAwZBw1
OffgsAKXGiNFQAo6nrrkAMQv0DDMJXccIeeBR+B714jWKksTe+AEiYMWMuIq9Q5jCo+LRioetKrE
h5oN49cAk4FZOVr9VfLJsGMCEsktmBlxQ8Fj0Y40++dVzR/0mAbZlKGqNujfxtrVtBb8xKuontD3
e6FZZfuYYQwbZA/lbhqetF/QedpjW3X6UGLGw3aqs4U5CWZ8r5j6J1jjQqsvTs6UNCH81FO9t0an
QTqgZ+3AbqV+N0wKIr/f1pzXf+//kFT5R2lykiyAWyuTd3j1XA8uAudktPIuCrXF8Q40stg9wO12
8m3mPE4RzVHCX6djnIoB27al4WHZ8izugbVlu7ZKE6uFUlxdFp3VR2y2XgXPiTCz1bSRhNgHoJR1
E9efqag2SdvOSTkQpyhlupGuu+HVTNtLFz5fwD+WRC7yQYk1AfH8AVPlQEsR+b93Hc048LoxabV/
GsuURMc2aoVc8q+bkrTclP2XQCpEWgVIrBUHxpm94y6JYd1VepQViQBOuZ2UxB+cHf2Z9UEWORp+
KpiQjpfcUGddKfMq34V8k764i9qzyFhscr6OhtonHrBgGmTKXauL87A6aGNVnpSG4KkDrWeDeoRj
N0lvoRJ19FK/YOpSI176c77QyBv+1ku/U0EvgiwSFjrzFl+UnaLftO7nIAUOHom0clR0PEj2LvmS
icRqFgojXMIZFGx2N80LV2Hm+FmSdcEZkAGM7x5kgOCIs034RyBDiAmPr7VW5hGGNOU51PeoU4VI
zYJtcVCpcPDn1k5D/2p88kyWcmwSrwfDWYjuaEGgAwnqBHCPVMVO+6mj6J4k+sm73FrXwLjDjLCh
YuI0kx1fsU7bmhNL7enalRc8PAztQmxYdMPinrneyvZZCBQsuTC965/ebXsg+ck+AHkcI9sF6w+g
Lcwmo3FBkheY8zlbvNZqofm2VVe6id+0Ly7eNZYeSA1scPskQ0GEhDlq6ATrT8cp7uW7Tj41ugVC
TaLIs7OINYz2hDxLM5RRnG5aXtWXUuA7DBxWHRzB074v/AbMYuLzxvuitVm7LoEHApIN03pjd4oG
CkPkEthP4pIiqq8V/pQ0XzJY/afeV+EuMo1eEt7cbR8LQiMYdRgkXXh7Do6nFBYMp6/OZDKCuPxg
NPHd0/U5X2m1aa+fKqONG9i1XiqUh0pwLr6+mwbYw7c0osKjX8mv0/EnsMb2FqIWcM2pDuuhFnMg
maf8qePjBnzctkJlPvZMLwEMM6fjOBmuv7UXquBqT7Mk8r+JrtqvbTu7d/VnIRiz/zrA/JKzM698
mfOVc+La8IJbPmo+0vHteYW9o68yVF0GxrD3IinaFvNak45SF1CyCE8ch+qxXImDhhgaKU70+Ghc
Eeew5EnwZnd0OB06k+sanGXqajJG/974XccQtYLpn+/WEmWoQGrnFTThGgeMnwZjz5032enPo8Gg
Yihy0tec3Vv5yiCYh8Kh6xuRmPhUl0adYkOzpbo8chgMBeG9HAAmbSY3WG9mDEirmdrIqtkEhvtu
zvlDA7AN62WUCqyAMnJgMzPcVz4ZxW4h4F50ErCENMdxWiutwFvTeVdrMJ4uJYJXZB32s3UfyCn3
p7FJd9JAfECxnFjH4eiqUzjg2XLQbTdIauP7FFTCYv+Ied4bvFfzIeQd/ppaKVSYqVeHjCV4D92U
dGFpnsR3pCyjzUxrcHa6yyA5c0pmDI/yOuY0nEoTQMfBHlIMWwKMk3uafdMZUOG8LIszGqa0mAFk
8Cj+ZOzi/Q1fb4+X3ChSuzw2v8BgIagbewm0+spjQskhpNK3nfqSDv52N1eSLX5krioY3ESDsesk
VX/b+YRI0KSqWWyxEv2YtxXuu9eL7o5s2Okeeh/lkOgDG854RxjEnCd03tfXuga+0zmY2fOQkTwz
5sTCG9W9bjENUh8gQpGZK9CzxlqoubGgf/by1tUdAIRUWWRYoZtXhjk+rxY54gGcXx95K9xTW2Rq
QJvmV3WvKNsR2kqC9NB3+7xrrjMlCZASvO8p9dkw/gxW+8b/gcVVpW5KezT7iCTm0z5t5yrLUn6j
FNruMdlcxInsxrYx7/Q4Tuhbhk9tuTFHOzs5xafFnI+5gL8yOhtp688AeCNM/HAgfgEQg+zOj8g9
Hsl2A1V3sa2W3VtQx30d81r4LqueBghDtkerIlNR8Uq2ybSk1YpaS+NXepgJXi3mf+NbBinMMv9I
wIp7Yb7XOusxyaZEKzqBwd6nS6iUpFcuO8f+0eY/KYiz6LP1ha90F6F7/loipoSm2pfdvT7vwCSR
X6sNhd5PVbTQTQsYvYZprDk0OIB9NLE7GubJ9XwEU1omrEaiac40RR6q+Ckfw2NRxuK6BRlXNtk5
qn5nrz6F2tmXLqSEkNhsUOMf2uz5G8Zu4NxiRUMjEwAQe7DuSYXRsS2GUBQ71gSoZWM4BItTCSLQ
F/nsoypAR4Wy0VS5Loy5Tp6/Oa4sOGowCeR+1Epf4rCp9h8Y9rqjg9erwEAFy4M9Sd3APQS4rSI6
HZX2Cmmzwc3lWcmS3AHVWLSUOqEXR52JrgBsAMdcG7qPNEKxsXmYbqv7U70fuDtpZWSogNrm/uu5
/UAQN4/lOtwVyGyQK7SXivsq5Zck4x0RyblWk0z+qLK72G7Da4y6WKu0q9RSvJPK4y9rkzz3yJkb
qKRHdwo2/J5kyImYxJk7HnwNVHtgRkpUKvHQ0fIYakVytZDinlEE/sX6XO3LWaEc4woMsUo9RjMZ
5LhQKRSFLW7r2ezJ0vBvtlbiCf2HyvDWYmb5DkB7voPb7fbcyhAFlombNnJEoTRpxq8ZRLRBWKZ2
7M5RiihbG+ABSSInOAXd6vuvS8kC1bXJ2a1zBDbTifuMlaLl9gVCBWiBPLsCj+bQE5i5AVWndSL6
NgL1rCdWUUEEA8nrpRrshE7FIEQMBnZDEWhDmb+45doYr58EM8rAdYzSgnRe+1uPYOoMsOcINP9J
SKjbWJ7PwIeghDiiMG9tFybR85TFKns5H2yO3rTkK9GiYPLfJ+Eq0l8WGrR7RTsrnhR0+vCqv9Tk
yvVGv1zIR4VKdSppW1/9VT0xvQr+MdLu+bPFkEDVDZDPzfNRaJIquE+qiQylDXaDtr8oq9HmdN3v
5cW3yjehagYFIzdFORGxM59CDMQXUKa9lF9LbFd1tYz8VocP89wRHrMQHQIrIuU8QaEaQCLIkjh7
XFa4+I9K49vuZBXlznH0dxfSCP0NMzgD5VsC81lnVHBWPIGfy/Pbzl0JST7xb1LSiXdQX6SeCc0W
owUp35i2zsydCyqxZUgHVTRoKzKkqBaxgTCMD/UAtU9hb1XR0nkI0lzi/VNoIU4zwNXoSnlxXEgn
E6+S1WL8FmqXkpYChTz2QQpYuhRQpqCgrvPLcv5OXmwLAhXqqzcqrsMVYWvg82Rkfd17KU6RpdWi
ZbjuO8rcJKAlW5+4kFJI8E6/+iQHZWKc+8G36daZ+3M5E95JFO4VuZG70ZEOYiRWwI8jwU3Psrgk
nhubKapwpLj85jHO3M6rhm754bgVxb798XwASUuplGwtQ92U5inWuOKTDqQHyLNoIJ2wS4+GOQJ9
M5OqddUrPm1Tl0OiTeH//VWNF/kGvY/AT3XSf+l62hjF+co37MUJ232IeDUodqVMAf4feLfEk4Nq
mhbACuRsYjoIoi00fPVA+hGk/1aWlILi1PLACoTEpCQNkIQui2nv8tmrJQzxQisXoQDUw9r4Ibp/
m0x1XPt5xr0OrmltxtXkEbEb3VWVEPNqf+oUm0xPHmk7BuDmqC8ampAFoNUPRmAhhWHTfrV5VCoh
aEtUN6+FBqr8I9VNBM13Jmsl1g1HVjYzr7eqgdHBB/92VOQk+0Y+Z3L8LGavNl6JSZgvl5lnj7oa
yVLnXKhOjkMb4LRPGW0ihHhxur5NvVYRScM3DApd3vBhc8JxrC2mlsmqQf1D45MpoNTKJt1bwRpF
PLkR/BTp6GjAtGq7HqJw0SMgina8UZL/H4HOIdJR/b46EmGGGYHqnGhb7P5uj5XL29U9jIAFUlJI
Rfh742lSQM01erm4KvZ8n1mrDQON5FOZy8U98GSnNB0PVKOfaV1bK5CZQoRMiXBgELtz0e3hcZzh
NRUu8VSO3KKVvsXrrNFZkew4px/vFX6gd3rp99/Zpna66mkm6PMWeLQO4pgaUdrFO3079kxklZow
HJBICD1C20zhEakdoNh98mtL397GS6yoHxjWu0Q3FiJRLGe0RjCXkOI6smMesRyk4dsUzR83Ds9g
aeDdVfW4nRnfjwDtz+pFPq5xCSMnF9R30/4mVQno7UP0ozJklIonzDHiSs4+ZCGLzyjnp9nAKIjQ
zcC059m2dOaAHYxW0UYiLbAc2ZejLiE2XVUdruiG9DwRTVRneovomk0hR1vft0XTrqLBt7xAHuZF
5aCjSlc5ViR9pN3cFS4+qaLY0J6WC8KsmP/YXkryVU9/ZnkmUQ7aG3o5zxkjUWcCS5w13vsejJYh
N2WCIvT2/rvU/vudWTuaZK0mfBjXP4V/1Z1FNALAC2LdVsAB1FWNqQapuMeVCfEYQYm6lUAraYdC
dWd8nIrUePgAbDeCcB+MHOUexEhNfb2frhFUnjQBchcLU6bfq7qyETYOQ65lprOAc9SKI2PUdkMq
FZ0gojTgDefW0T5Wu6hgXQNlkpflsvQ86S1J8vz/wFe1CFda5KAM7/q3uVTxGJgXUamk/d4qVoqN
uCNuNHvEDQVM2DCiR+AtHU4+7lpTNJ2FcJ3N89JP7ietf7VfB8CRQoO3zNI8hEQwXoHujvE0dWMa
ot33YZkr4YRWil1jl9kCdWCXrlOKKp6IhxgykelUyP3i4QecmzS268Wbfcz0GSIscetEtmB1A9lH
8CAAIIWTwvl1kvlWuEhTBicDPY13+0SEgyRty0jZ6AdtMXhcj9QTNabWgBII6O1I+HUfLUokJuE6
EbLsZWk/P/B5Q7DVJD6E6uVkI3GGkEc7ZwhOLTKQYfZmCBuQT2DcOE7/rKylrHtqkKSXff8NXk3d
lPb04gJtlenzVIFAPi+m8tbo8hltO5DfO2zXA9/D8KLQaewVFZCb/PORQzeVh4wq4C5j6xI8maMC
bwCyOHFV3h8Sk7Eg89l3in2pZYqhOMYg/QgeC7BAxNUQkTEgbNS3dEVhYH5l+1wIEUbu/quC9XSP
m877KsStnNSyBTxx/i/XRucwMi+qSl2vGffktuAD9HNacMICU3/lKZSilPwMxDyKtIBvCGiFzROX
3LYt+g8v7V/DWI/AQJ+YCSKDHgXmZQ6MONfeeffwilOKnBd1umP23k0ikvS3m0b44fOh2Cb224az
Q6iE6JGIBZT8JkJed12LzEZ4EjjGtccdxZYMHTLlONGORkAmJ0jw6Y/bZS1JfrypTqxQ5uemZNy9
X0HcvDpIM+fFkp/UH3/Gb6NZARkUTGw7gjjxe96aywBwHUROvwfaRe2qT16G1Kd9hqsTvtinjNlU
DGKxTlU1siRwVUFXnR/31kXi73WwP6vRKMOUlE8r+m/DRu+WIt6J+aQCstLsUmuiTiLYHUs9KCfS
LZQDFxa15uYW7yGy2hq7xWJLd9qLRBYU3M7Rk10bV4vJMVr0l3JuAmGpcjkanL+f/ybvMB/6LAX1
kEi/71GrqE7VWtrDVDWnxqPDqxckmy+tuwmo9AFL28w6pI1CTMlaBmncT9uaK+DRSN/z7BDKLrus
+X9rBU26BHahzV3GmaO6F68raDA9ESqc5ZpiRtog/+4JOSkdZnAIy5/8/BFYJDEESgyVL5s7f71I
79Mwg4/kuQ8lo3Pjqyco0r8r2wGvvCsnv6Uq8MJOmqi4TXD9Nq3Xe/gjanKVb2IGZRJbbkVimZcg
lP1AP5dnkKB6zFGI6u/3bE7OPurt7Q6zmpC/j058fc3nAC1Lf57pi+4hBkmDvLhb5D2KLlh39VnC
qkw5woGsdePFt8VlfnRWXlM1lSc/ht7vklQPFh93IaEQE204D6dxUxKVR3FXm3B0aLeSQkQj/Loc
AUpTCRUMJiE61gqichGtR+tXZMxVeNDa/o8NssJBf02DFTR5qiiZxQElTfcrufBRq3y2A+RNJGfG
N4gIV+QzwMRpNpCM60s2+4BsNA9Oyphy1Q0H1ztshntIQaDUbIouHJTVgX03X0W7fQAbmLp0mc7N
LemPlD1Pa8oRMd8ahTlRAiSZfKn/k8bPd4nk3RYkjArjmuP3fLyDA9WBUaDvrx0T5b0Vzv7vDPfM
0gMpVRPgcWR6hVmnY9CAkDe58EUy541/QmLmBXaWpzs6ijZ65TLeNbWhVMmkIURBkDR2kiRlLsWO
m3ghgrmZ6s6imc8RfBlgGWllVeZpKMApBwIqFVzte5X888bTIOH6tdzExDEK2HdEoVMsDRwCwtEu
hi9wdJB2vuHDgsKtp7L+n+5lwJcqOGu4eXG8V0N2gFeWBx3jZEDuzhgHorf3Y2RBwQh7T8kkvnof
LM6KTbZXtKttnhrcSmF/hUWptkpwXAC2BdItV8RHoC1s2Tc7dWi0GQcp0yTtXkcrseJ2LTuXZj07
BdTPEPszNXU2h+QoeLZo2x2hwjKJpzIyZZRQRBwduM550Ly2QPPZSG0Qm7FnJW2QBevuwXrezwWb
vtykodD/nvV3Emok5LLGe3rdyBkOetyVXraqDcvNI8b3cU2KGNBmyst1j3I/ULoemj8tF8hbTV5f
p1LXOTUaaPd0MHAliDeSoSKrHUjW03BwdEIAv0Rrv4n0wKE5sl+IeRtww0CJUQT0l0zl1/+3AWym
lJhEBFpcI2micRQDVHmKy6KIX6ODQ2TS9aA5JhQ8exd77IJcXVPOMl2PYd2Vb1r6AX4+DtRoMc1o
Uhpxb9IqlHPbOAb0lVFTWYI+72Ao9LHfLYQGUoTdBD/1Oc0SmhI3O/Fr+xNrDvhM09lfyKizQVcQ
hZtfMivC3LLgiYPNo4ufYW1hKlXhJ1/wB05e3maLtkurnKlSa9w9l0qPPx1ClZhYzQey6NRspGwJ
dc752DvaJ6zzoVg50iSNcX+cun3+p55OiP3NYBGSqzHrnG8+WbaxZiHQpQLmf2XaCAjCST0WBg5A
qBmOgvMebJooqrQIqKob8d4DsiODB456jYmpX7fbfMQaHHIBBVKHg2smLFQQrB/jCwwhRiYi3caT
jitMH0QZlRNJkLRA8XWBdWOyLitHufKf0zuFn7tg2Rup2S/r0Kg+ySYFTP2MSdwp/emF5tNplTsl
17miMR+/pK/wBgq/no3Wy03t0sqeMBuUHJyewbTjLbPoC8+hbYn/0WP3/GItpUQfNcaqiMDs1LM5
8Bv+MBv7IpmJ5f0nImR4Fnm5un6fusjvChTnwVT2RS2qnWdux/0a3zUZsZ/1ko62vngjIed9YesX
KMTEc3Qt5k/jgLW37RmhNHplsXfgjM2DNYr89zYG6r2b89pPco1TlwUk6utrsib1gATJcgbDE3l1
qzS/HopFIKifm13j9vI4pn2eYj9Tb3/NTZBhj6sUT645vsSsdSIGZLP0n1XRnFaR8U4ZdMjkvyBx
4DVmQPPncEGE1pn91VX1MkfDexc8jnpzu3hJsV+0/h3BFuJbe2gbG7mMWRX+tB0pi/mDjU02h1DE
8MrF5GlemASIjZA5Q2O6fYssaQXYo2di1WTpHHs59oOTS55OVUTqqefSqPYtNv1Jy+412BWyWIJ+
Sss+zG1tzVSm65Qdeja99JVEfPio7wgWDgY+yddcqHDscO0L5BHgtGXIDIs+J8rLq1Ez+AC+lGRN
14KwVWE7ZeJooq2ixdok5Z4pJEoqwFDKkPEOt8uJ4qv90pw5EDeOznL5T3Btg4j6VWydaZtCf/Y6
DQ6v6fq+1PmjgZUPT2tgrrAseyzgavU5Xa/w5XS0fPNcuIvpXOUsTR1FtTDgu48t0PCzCtlQdlTF
fiXakqc0TRHJp0/KX65c+YtOCBqHCqqXVABHF2gbPPyHrNlBWMRPI1+xOQoBg3fkHWGDStt0DvpZ
a+osbQZ3Z8AQ4ft7ie6Gc713H0IGnVlUXWWepH3j/yj1hxhzWkKmIf7NrXukTZvar3xJM6KCEDhB
Saa4RKXM0AV5bnxuq5a/hZEhy/XpPET5NmdeDDDOvLfMMR+WBJ9K687TiJrgre4AS9SkCh0ddekj
uZECxK6IDCID6UyUgwYMZGtkbtluyw5hy4PW+yfw+YzkqvbCTsTjvuZJU4xFPDcyBqNw0HxmF2fo
tONEajiz3TxIzjw5I1JepQTNos45/ip2nJmjtBb98s1o6YKkSadoXXO93AQlZ548KZR59ZStIjz7
JoQvPAknBuNAF13ZbTwGASADUJhAb8/7r5K4mWyxiXGIvu2pA0NFj79wDqa23qyh1p973CewywrB
I8eXHthLvxxD2SA74x6nfJTGRvktv5uK/t6qyMR9JzS3d7ka2p9BAN1bxSSPO1I7MlSBEVRTVA4z
QbF+z5d4aj1BIgCa7mmVfchpNZRgpmLNsPYgEzMsHJt7GkMuE5Z2wFiJj2nyw5lJBLilwf8Uzq+0
RzP/tHNgvS9vOLzj3nP6lcY5VA+roYXgKnt7On2jZg/lWE9cy5PgldHqzGyp3VQ4rhIIenArPf2t
Nzr5HBFWk8OBfEy0r7P3XXiMoiQG0U3yQFfpmwJmgCYALcC0qOL41IVYofseiIaUmXrGSFcgUDy0
7tqRuRlxRNsRDZ00g/mUC1wRfqqd3RAytTYtNfWOGJBtQGUa2/IkE5kib8TWYDHI0VvYX18luEpY
ODoYyr+xbbIt4h8UCwefS4razmBX2RZ1goEjL9XSq51Y+9j7OzB8VWyNKjeucJ3B2Jh/5GOSihXp
JlV23RhoeESUS4mFP8ifX3lIkKE5tlm6oJ+4ynJkBT/PqTQLIWTbMDsogeMjlqkn08vkg3HGGW3y
w0gkUfVz2uHqjdDHVyBhHn8wLZSBffcNSkyR8M+hJKLtSnIOcEDb59Jj223qPGYESRhXuXidNUSn
Djop/9J/Y5bNpIP/SNlmWONGF8R3PXIXdvMhda5M9OTwOelGaqxSOBdk/8l5F/QFOsPfo/o/xODg
uXHPZYtlQU17Tb2q0IuInIw1ZVh3h0FmtbCaJKzcKpniFsxMWwXRpZ5IT+T3fUWQj6JCVW8w37zj
3poxSx5mhq3YM4TW8KvnPa1PI5NB/PMJ35vywO1DgjyU8lmWr3+R1rK4mX1fi0wXAqh7A+/00T5l
G+jIYKjQ4TmcOFPF8VWOl42UcxpQzW3ZL5GpRQhHcZHwIAL2JHF5kFradtOMKIUZgksafIwaXUYy
frxSXFF1w4vl3qCoVf3at0I1Hfe62ofhYhMWp+yOKefzP6deJz7oY7K7dY3xszK6wutrER+VAG4z
vEm7Jyxd3aOHkR51f7RQUELMI0Sd5jCYIZX/WqUAaC7IBaIRzPRTz9JYdONGm/q3qbxs0hJdLHMr
bb49dUpxWsFNNR35Ve7QtjfVz+s7cFa4KpkE0rDWaUXVaO+HRDOUivN+sg0dYgw1lE3U9WVvCgty
sTFCsxqstVH2faLDs0d4q1C9TRS2AoQTqEBf0TNygHOPzkdxW8aqDskRx47chnefUL6xMF/t8wy0
80+ESZ8lzUst34s3dklJqxQC8vy6rwd/4iR3orLEPByqzVbe2z1gUdmM3wAXPumqfIV/QVEfHD5E
0goF+YkSXyyrsXkp7CEsQJ9HsWEioNJOdXIHlXVUN21IvnXmPADFnOruyUZi0Xheiq0bSfVSfTcG
X5yqMPCs70t1BEOdf+5saCJ91gWaGqJBlMVCUEyXdnhcoS4s7UZ7xmeaFysBrFl/nJVAy6gpyAeA
vru3jv5qISJAd/dL37lVBwSF7hiqM1yB2zXcVxlQlgf5iiq6aLlS6vABv12CtPoVwHK4DH5tRe63
7xePo2LCTQ3i/fwcb5xa1erPvLnNcJdr24JyyrYItyRHIdOZB7FmrtdDJWX/9/mmr3ZC7aPUjJ0f
gkViYFlEr+t3tEK+1g0w0Qi27eDV4XveZMe9qF3OWZRQ2tp6JbFkccUpQFX4UfgpD0oxUj5Q3RTf
TRGk402Hi76H9uT6NuO+RNPdCOh8OSBmHDtlHYJ9UTWqAfHW1lVXoo74vKnf1PlQjtPWhtW8unSI
ibMB8DIiX3XifiYvDCDESycxXKdDgurlgsYU7x/duIR41za6ssjpH8hRY8vSdIqM4t2RD9M5vmL1
MlIvjTKNyQWj2r7T4eHU/bVAozFW7kwRv9GGmllGZOvPl6GomkqIDKc5IoHx9zoWdDfyyE6xx69I
RRZWMaSL8bHaBNBUNKBJ3Q39K076+rv/191j0N626POVmzsFF9VaHD9a3KIM1u8apwkCvcdKlL/B
X7GjsZaX8KFZjEv/41lL3zpxHkxAYn7UvXMeoAUK+/UuIkoswQSRJus0R9AP35/sZ80zG0sRdzth
/iF+nExzRfv/zRgLi/sEM48zAfS1vF8WOc7GT0qdVuXAYBsrBYNiChawNYgzvvAI7A96ibv2lp9O
9quRo9MUblJtqPiTvfDyqLuHTE0YHjcanEuGtMIOT6wvb1LKjXZ051yg/dn6JCi88DIxbcvSWQY0
tH2E5XHUyzFU3tehN7mUKDxn33DKs4HU48DjQUCiPQtHvVjxmSkKNJaq0V4gaKHbKD/IU7+zNRqU
1Ho4twxTlx0EyTBNjOfT54OUnhsU6OFRIl/z2+GW1zQIJQhXOP5CdQgjA0VY+a2Ck11mnBY6kq79
d6VdrETvD5lj/u+dmkc7iqqLFt4YJT38GVzDqj78FOBKqfBtcPSMSDwSBfbpmq1Xh3g96BBIwra4
MCgqpM4WWpGaoXzFfLrJNUUSnjx/lIQ3miBMDS557ZuvE6DyZE3HZondOltJYUaBWBOgLFgs37Mv
N8E5Age+dT6iXwxzIj6fyB1q68Ywkezy18cTt7xceX8n149n7mcQGcv22HMNeoKwuzaERtdzsXbI
bXnBt+Iw01eiW227vISTNmxR9Ds8GgUc3QLOZJDVrenU0AQDcaP6rPmYbkFw7YmJfQNFBDLGC7eW
nDO4TWqeWhZQPrLbpkCXpL2hP9o3Yd1mHQ6LgVGB9H+8DfUvF1Ihhvl8cpOlNgBvuU3a60/s1oyB
MwsqPZJ17SCO/GLNctZK5lTVgfuBRK7QdcZRpIVgLuJmNselEz2jHABLnhFmAf7yYSgyyu/tyhw4
XDZj8+lO0lL9mlet7Rbr6Y6SXZrMGH3nEZVVGe9KiznvMN1p2L36KEC6otxkqmYtVpVxIie6GJ3V
GiDLvzNKm3SKOqJG7hPRGN84wn29Qk9A/tifY7qJALWR4vJKUh4QzyTtw895eHPmlCYxBLmrGc1R
9cngUiUwids9cEaDNyW0G0KTM3yI4G9ELZkHyWHlS7m5HUbT5lVInA453iBi3OADbQfldyCR4jYp
OaBvyVwvgCNBDrkjjU6UySHhsoYwVLPCiz+LK3rViWX2cJTIzWQcGQOGhCcfuC6ADZ9E/BXs6st0
zm6jBdNEDsoGETCczBUHEnHTFQX7UWcULsFYM75AhB8Y8IFI3ae/fa5BuIMK/+BYc51XV3VpMiJB
BjfGuYkzoprczvlWzNqBpQTVS0vVMWqsUWVDg+8wFg+z6ToEGCAIqfO4h3SwSJCwf4XKgCcNVBnu
Y3o9X/PZ3scmDdzYNZINs3VcWVgPDBzKAUh+adNx77LLatOMdCYLwV6Vg3UzVmrajuQLwpAJRtBk
d3JKAGSdd84f54BgkNY6judTK5piq1iZF2g5QB+mk305cNLgtoEDlkeVzIZfH/69zEcZwmOseJkJ
C2p9GxEdqJGtAaM/SH3vy+hThMGJk3gBGPRjNShp7miX8D5p5EjquKLm9BkMw88HdOQNE16XQxPY
ddT/PM08q2mVgjv3In8Oo3SoH0yqfR3j7P4X1+d6P+Inl4d2DDMGxOiCK2BmJIiPBmeImVQYUna8
Ix7VYElviXrE3wgdsiKqcceIIL+0pqX91EqDuewhdRTdIGUHX8unsoASl4lDEErUGs5W+TNIGBO2
jyhGZyFUgVG54miHX/80cyIFQTC2fPqZDVw4XpKCYUVeUK2Gr79RpFC2kgdA5+8jTXBuVkPoJvMy
3CLREg3jghTeaNsbIWZ0SnuAmcOBX6EI36Wr73WS6faCFADypITmtbBRkO7dpjmay0mPRTG5CiBa
wOAZhCHaK3KPC4hXJf565YbEzCjQktDnkUZm6hn7/Bi5X9ATWXYrUPITIuDPSV83ehC6mB8BeOnu
7SO07V3ozNFSKclaMXtLvSsWOT5aOrzF7Y6NKeT4oIxMR1iwe9J1DVYA+WL9DZq4LK2umlOq6kuJ
pKzQ5VWX4ZuEIJX93rsep6x2BfqctlWQsR932bWFHR8HR0Z3jRrJz6fgKbgTHNVIRYbLtubNe1D1
QDzwYftfTmdJcZVI1HZw93HO3alGGG/ymkj13GbwkkF8lQDZXbdr1FUtD3X/M7wZFwRSwh64/e1k
7UEcfIbdG0N1kNN8OX0j7l+H4cyX/uIFIJW/Ly5kYgXvc2SXWOz/c85o54cd6YW0cZVVR97UxHOj
GfClgH+w5S2lh+2DNaLTeKgmcYjXAJYLbLOGbdyNs7UlAmRbtU9F6jupb+bC8nJ3v5AZ0gp6QBiy
msVcJzHumYX269Cv6wenlMYRpeVRUvjrqjMEmhlCA1ZxSJXYk9ZDtDYOpIkuNZTkGBCdrCro+9SY
HMmWIPW863PWC69LWn3alvFIknrCe4nRVYPeLy3YnEBYOY8zoXm5Hzz0QXQ0rbeHKBMXigQxEd8K
1zfudaE0wBQS8GxerU5G3HNljPTnYPFEDHkhvYycpTqjNqhHUmWgqvUx8ESs0HVd4elQNbtBTnj6
LrAEuTQ/4xTegpvzJVx4NCLtrZxpV/nfsn3oS2APG5ttSGZIACgkTW7ECXGGwQ8VuffYjFgf0UA8
YpenbHanzdOG1EPrUUt8BKPkrBSzDUVhLXqOslbE95BBYdv4K8dqonctsXPo/31zFl5aJoCZn6DT
uqbGuKIAs6m/gIrDoj6MSf9pRgoADjDAHwQwuZdI8KtAkhR5iCLWH0lHAbXOUOtsR43TNhHau9jf
Gs2jP3V9+10p5eVjXrJm0Fg4+pbVTk1FS1SEzO74UOhdBY3LuR5hjOshUWBr67zXRklDM4HejUrf
MFXD1IzhoxOCW43ZAz2j4d/BdRsKnVMk3+UKKuq2jbI4DOG3anF92MuQXK0Hd0DMEtrjeIrAul+0
YqDxekPSbt18Hq3+DuxGi3r6Mb3u10SyYbTDI6LqpuADjE4n9DIAvGURdN3MDKcbOZuXMlT6KIGw
h4I37qq+xYrdODvDQA6L/Jvc4UQWO+bwsursTsbo+XCtK53biwOeSOiZmnqcfMWeMMW9Pj66UWwc
H9oJFn+fK1pKccV8C4UO9HbT4O6wx4JRxT0fNespKocaHz2jNjU80UhFpEWAWOPlRIBj3awcKZoc
A8kQvHY7XG1XAseiJgnTUe+7SwGtgubbcxJeLvxchzflj9Sl7mKcUnQfIeR441KTDLzpLf1opLGk
+BwlW2zsOq4Bs0N6ZmAjfW8nzx9NDwk0HPnoaoEQ/vec4QVBGEP2GaCyIWIvZS5QcjQEoaOPi0SC
HbnZLV1mfjpippfTIOGxmueB1c0rrU9Htjj766DrLRPVmIirIyHARdt4cQ7/VI2oi8XbcOthky/E
2ZsQ+GL+FxVsTMJafP6pZoJgUiLW3QykZxXBXjGVnqYgkkC266wGURMPUjIxhKgC5jAFJbIQO5bE
P2pNi4jPnKwfPOshO4plHBCwrAzvXIWLqH1SbwXIV8rnKXWYxQ5YqZkjatsYCm4Ir4JzQeJ4Z7Qw
4s2AHw6S+ym2ZYFAVtqCZkGKgLl31R/625szeTSH5mtUe97rdmBIs/WLx8wWkOnzxM9B5tvzQbeL
AhKqxch7RLOeS7z7P6s9dvUQSpA+xdpwexu5igHQY7YwNDIr8EOt2RMRA09mZ9i4C3G3rgn0deco
sxdwjwY1c2z8Fwewwf/JRwC4kmak9R1J0w2hCOyWooC0+LYFmYr7pEEF5ycmd5BXYhdeZTnqaqh8
2mktu8E13fev7SrOwLENW+qTGzxQ7rUwnjkIA8lzOLvM99egkIeQi5axLgIxliB391opYs6l9Mn/
6XWliFCrRGnQAvI6ZlyvoBc173/PFG+hKh6nijz0NVhwraiOazLJv2fDwb6GmL2OrbchDef63E/Z
GcsSMszgaqa62GESNtTw5EjCNR0hMQYpizcjMe6Xr4tAQMxqYFsW4WkhZJ8KAnIOuoZfM+oNWIcK
iPYWL4h2icPAvcsy9rd/ZqsJzsrHqJ5Z8oVCUPr15PF1+jXCQfU+no1oA25JxYHEphbqzyk0tTI8
EPQ4m2dMKdXiMOj3Tjcih5A1Jfg6I5Olv6LsWytqmJHNO8kMpWJPN4VO1UW527gnL4sA45UCxZvB
qFhehX9QG2JqH0Cey2HwVNOW5nSz5kzHKTorAkiunYSIzw1sADbOhYSh4666cbt4vw3K51msj2Jf
+ZFKK+HUY5+seuB7AeVLi3MQKKtx55rjSy8SeQnZexxtxibZim8aziZQJbVCKbzJsfZJgSO6q7HZ
Dy6wLK8huueLgZz85Sca6zNnSILyJ4L7MT+4hqfjGHEv8tO3EOiJUdtiyw5gGnIwlBjQQ2V0cnLO
muH/GZ/JgxZ0eCSXUsp/OmBpYR3MarpUo1lkxJJmAZq7h/JUUig9p8js47Bhqa9tGxlXAgWcb+61
dVMCxg5DrJkuZo1+/2LhiX+VTGXYfgY/2e4euZ2HlvA3VcnAVthUBxj7pTDNqWdZk3mwVl3HQQK8
ErNTTbA1nUwKD6e79z8UUYUg8a6Ai7pA++I0qi2smn9Lf95FKdDU/I85jl+hDbgya6ba7YoX+RIa
gyGdXowNFSVNnm1dezHkA96vf+uuHP2HorBfTkpcsNOzXSNQkiIB1yVm9y8Uz/88ujWYdEDdt+1E
gDmmA/V9ZYGafchBB1LXhwfe2d7an86t6HPZTjeXezzuxi9l9PrsgvQNxhCa7s/38IIW4xzHzcyy
s+lT4JR7D7LQb8F45tvMaRG59WOHXg/b/ZE4Ad1fJOh50VNg8UlknrI/3VcObxmkp3RHphFHtQfH
NtpTJc5eWA0RhIIOw1IVtyH7MxgdeRoW/PNPdtjD7OY53KZhPGuO4e4x8jeYBLbFht6O5/znjzRT
SlnVeIyEyJyCzGJXy+izIyar8EoyUbmzXcdp9Yrjw3F1xQ0euTno0cceYsPUxyRGxSFhBZicPFjf
lvMeldBmA888LyMxBzQetyqlQoliyur+ioVGx43eH2aGFqYBWyAR6mhTnZeofi81V2pLDY5Dq5jW
/3DH8+8PxC4LSAGUm4NrZzRNJnw5pOYS0oDhgd14rAy0RNkZJmmJHt5jxrRMt4S8SSE9gM4A8ofi
YJODpcxOE9i2ZGZdeT+9m5mXYEVIzvt+Jpu8IHBjsRRNDxSXcq0Md7ykWMbP8+u3xb3fsgOXNcqQ
pkNgpT8kpJhfcmUYXNK3waBtd8+4tjQxHEOEbIOxEs0yCWF8DBp49oW1dLhQezePeIYPbRsaqEfG
W7/+B6WCoLeXaEvu7pnbKQiieFuiJ3lvmEOdRKjM377bVmzxTOU2iHDuH94ZS25/TB19axntFjxj
BBf27JtDwFrYYt2uKmTWCmOX+NhsP1imJIOD8tZIc2+Al7xIn+UACiDbfKvytw+hPUfCXAPY9Eo+
hCGIiCKTqwRITXS34+2PdFPA+fLqAuXeoJtiGCdR1/Ssz2r8G+wZJ1er+zjYE5jNauSdp7SHZLs5
DWtNBvdgRExpHoi+RsHMAAtoNa7sbsktJL6jq2Cn3L/cYPB8jiRzMW6Hv8nF6zoERaHDWEqOOQrj
RM8KfSHSxzA1hJiNueKjAb/dQnhBlBJVGSKeCy9rEGj0v5IyprGS66CYLacSQlzginw0uT2R+HCe
8meIJwLfshxTV2Hj0+fTHY+5vV6bSEcPv9dTkKR1Pbvgg8Up80pIfp1Yu4v0PRmddfB46VhkDJKM
GBdVbszswnnTNvx/ldkXLuO5dUmOiCwKXp8LTbcP7372KsHwAFGwvARIbPradDH1VlEP+xVdLtGH
/UU8UjkeTq7o7uTSEbY0GPbU+vN/iD7UtQwGibwudmN0OEGoaAuqz5GZx5E5BBhQEh9jW0ssdE0w
3qkb+gV7czXA/byUrLsiDk4NBbeENTqCkY8ZQTfY3g7rVxc+Y7qR4nCd7lTO+hjbFcKRxsC4pZRe
7kFeaYi19aqid9QEq59SEcNOIzcvzo9kf8ha1Awur9Jf9b2Wx1VucB7CArYppT6DUbLxRy05T6o4
vzQ/I2FwSOs8GHiP7Rk2inl+KqfQVEsj0VUrPDF0vaOwg7tcZN2d+FHOdcr/08muytC4F3JNHUct
ZWUj/MygbGQyTeBDQLgYpl+0S0skJRssivJcMho8FY4EedwNE66oXJ1dVVO8h8GnCFnZhqa4HUBU
vU2htIjMeIaIgpTTbktF/e6bTU/dnDD1op+HdfaNhjE0q6lSLDTamMLQjWns10xq+z5tcXA4bBiN
OTsotkZ8cKG1XRBKrBiov+CN9kCcCbTlABYzIbqQbaEaGWksjcsOK7qaHDbv1KBoegBq/Xry4gHz
KK6Hm+gJs97OCuS5msfFcj5JKANxDtvbgY0ySY96QGmQSsM6xabM6FGgwvmAEa3OYmE57MYetrkP
kDXSgYKlnrqmoO/a0VgOLDDTonLTBz+3P2wkUiAjbGbsVQimsaoAAVld62Xu1a4SatGbBehH8YWP
CwZCqx8CJZwt8ni8UUwWkATFRYuLcBm4FsYU9MmUzPEKOwlBCfZ0p/AkKeVOQnZnHXRNuBdiKBjF
/osJTttLmkOe0OFgQkhuBMRfYUm5J9VZrR8m8iUWJT2yeb5GCs0C7InpKJA70Ylg8HtZDlq9Mgy9
67k6/do6E0j6Ofa3r5bGB6/miapp0gdTpIcKdw279gXvZv5IH80adOolexr9uRWX+HiPuxzChZgJ
7iBZlO6pnLGunQxIk7MOxdqkIXKl/Hs7I1wU00L28fzALGGRHkku1pBQlGI2HrPFkjMMlm9T043e
qZ7z3p1zybkLHbVXDhedlBBvP8iVYF4U2CdW0sfV5YIGL2tQOWWRsaiZbBw6Zmhlll4hMIWXxVCf
ypO9CwDNqEju7fv5Gljj3pTxaLGw5jEFPQfMyU4TBz7qzRUpC17SuVdrkVFhP+0PvWHCV1XOCOd0
qlP6lVij6FpfE3SmShmAd/F8TjY5SqclLepGDrKbuYqOBJcbIAJKn02JbYMyGpgfp7SQxZMxnL+a
GlDy/Yu2rIVZ+SkYUVmPiyHSawY9Okn1pRpyKasbzJIPlYFGYYfK+b460dd4WiQDGsQaSdhfEKW3
ZeN6AogBFPbddolVFLuahT/KyjLl4OOdW0wcN3RLus2ythYD42Bk/9HrwEcGVoiceIv+JaYEwBAw
Di3LgisvaAJQhsl+0z0CUYzQvIdNDNwV2G9Brk/j64nbC5PA9Jk51RJ9yG66NpQUpqVCTcXzjsPC
vNC+x4EjOD2Tms55tYNrFZsdZhGW5Sv1zZiG+jtSN1PV/i91ETr8RuNOB1AUsNPTeO+BBFuZrpdB
QvSllGIDYC3YnUn7vakRM9z/sx+uMSnTkn5fggyGTxpjPJL51nsXArbAJhtbIU8aP4WugJeG83H6
xYqua37ux/ytFg9lOcUGcZc5DLuhFpkNSMOrm8G8OxP44Xk3ZZEK2UK1cW2aSI44fo3xScdoSeS0
muj8xn7nPh3978UOwJIgCMFO9VgDZ/vmjCT8bmujSbvEDmlsQqQpvUo45sNxyQ8fEW+cqvV9wmEg
eMkh/vOnELw4JjOJFCnVoJnmkP8HwAtr+++bantBOtwXHPeiE9iUetQkkIdFZaAwZEZdGLEJ7x4U
8xt0fgpHGET4FYpqcymrYM1URrGsnWTfSxrPVR/h+MCTGgDQ/5o+Tt8UlLBz0wGBrhkJ8zN/q4VJ
5QHweYx+4tuNg/wORajKDYoaLi6ZqMTDFzI7tDjP6tgB3rVY8K3yS3WdZ1XHZfU9Lfd3suXAopHW
aRjrhiPUlYJWZSO6lsoXp6zM11sq/vEJeafovZYm/ATkUs4MzUw9V9M4vhiTepzPvpZ6ZN2kxQGx
x0+tMVP1OqPf7DWSECKaSJZiWdeGZyh0STG3iDWpTk8h6orFvGNgkPEzUC8FqQYAAacS379Y1+Yi
KHIeH1fmLS0ibERlnhThZObbkubpYVcK5pYsV1tb1lvy2LrfLbmqAPuBmyEIrEh/Y8svBfragEHb
TJ5WK4CooJy+IYTlP0pxWCoH26fV6AEWNaNuM51TzRSFOv6wHQy5U30NdoWILdaw5VWUDEE14HtJ
7NI2JgLBkMm7AgDD/u74VK3MDB+hKvVD/TtAVCntGpVhn9jccN13C9YicHseRN9aGzElzuqBHAc2
rO6FXzwr3crC7QA9bTDdNa5F5+Z7fwWwXpBRV8gC0M9jXUQ48kev2nBnLsE7rHJQCgcoVUkXVEQp
TEU0lU+wqa/9bUp9aqDVYJHlLxPZrq3/uVWeB9WfYsKH1jmYFxqB9BkRodGJRNyyDaBeAC3Fgdft
EyfOL52PTa68V1y2nbEwFvvGbV/Wr87GpSIP7nP7md20ocT5npTTTc6hmbVsmYctzZE322wkh6D4
7GUB/Z4S0zVO43q5tjG34QITe7qwzhbfQW8PBrxmBg12cN9BMYCC5ibR4GJ7TuL25kdGdjmktgGz
lFr4CaWWi37varKxJUx9OwqmXF/nUBxNd4/i2qr2xev32QaZEioytOo+x7qq+3sIMp/juTRuYTUx
wYEdyTBAgofXoKde/FLJDbtSDGCGanxgQDL2bgog7hxkxYumiEYLFWK1H45ZKOhI9VtHbtCcfbCT
+A5YVxm4kE+CM4SQBdxZfzue+rFZdcEMwREEIPQ+CPkZED4tHn8l9K9XyBxgXFqwJgu5SR0bn+9V
gpd4ZPVMz9r08kKLyuGWT5Md8C8lnXmCme1+unK0ytoZJdMVHzkC8qSbO7GczAL2Qu0sCQtom9JC
ZC98Ot/SrexGr7L3xq2PN1UGrmmb5jiuLJJW3hOeh7fmqfGd+IrXfSw3Wn0m2rXsNew9FMxiafVf
rmCC7KIOHn/ai1SgT9I28nPt385vwj3d2YLx72XAaXDLOhClsntkkbMdtdKBXxCVXXkB/1x4bkOO
Fr9QGSo9HBdfxJ7MzdYlj4WdXn2RchIorpuj56cYRJw56F2gyUmlO4f/hi4odU2OR2gDeDyzS0b6
8CBQPZLbqEudld7e0fjH6eeLftb6LZaSSMOxOkKHODiqBp88b8M0ursrYB2AMC1qcM0g8HGWRmJr
Q5qmcHB6m1rG/jH8gCdxACglN537689JiEtT4LNQ5F/ncTSGJFmZ/SR7z27rwEqwtd1V/Bbvr+iy
tQETO11JDnQedXhCRAfj8gTkMAb4zXqyie0XUZ6o2hSGL5HlUFLh3jNs2cUIwxlyR/wVYSCh7S9D
QmS2I7cjZ822EKfjNDlp3DuqZeGpAL2jvxZV3e2FtOStn/WnIQSDiWRnHk3vgx504D+N3Zln5nCA
gaEn53Bf4aq/5puM/l7SfVN2HeJ/VImuVReiJ6P9ulVLb4OHZwIXtQxCAQLdt2SYY5CIT+fIqBoi
rhqyZBaAk+YMyXF849o2iYeMglylM+ZrWwKOk5ZOLKd6oCu81HvAmFgIhh7FOtUekagMw93IDN98
1A9zNtPy9M2S1xjLDOyYZ27nwK2lSsFVM86xSzy5H9VVOkzz4pzqdQp8yyd4pLIP7Qi6S+SRIezg
Xa3VS70el7GDEs/xYBt6DOcqNHCgND+dpJeqz1NNet2m7TCqAIMF38ibNL55VTp8Pa14AU5o8K8T
W9dypv37DF021YEwBhBeYlMUCGIy63W93/RrSEFfK//AtC5zXuG7iizFotK+D+KQCkFosZOR69ti
beTLZeOjgGcrihyXk49r83SiobygfAlkK6T2NWiLx7E3qTJ5KwS2xBf+mondGGhosg2PIR4j6QJA
Z97Oxltg3OsFdjw6unDJ2juQ94MZ9lW5+wedKY5pxwRsiLQxD8e9O6EahvtDbZXgfvetR+ZI2K5i
upqnSrsGDRgpbbOKXDZFPxFmC9ISwmTcKWIWyNpFvdQo6IOZd1U3pF4vpwZrXxVXXM7eqj2GWPw5
wpQ6J+A3KQ2wT3+/bV6shxH0oCVJAuuobcL6YRwQGQ0ih2itanA+/cyBwM2weoik9d98hDCG7yD1
VV2FHAAmF66Hb5c49NpZNG25yunrjIeidVz/FPQ0Wwc+lUj7PjIhNthEUS0kJqq7su6X89Wt0Kn6
mXDJqm0TWqF6ZK54a3x7DgztVK6EXXKTXOyT5v3t2r+6uOBJ7f6oRKBttEI25tIcuV55gws/QJwS
wq1EBSJBF/XqTzS2k3wB7YTrg/aTsaVQbYC0bPcdoNJ+DnRyMaz6vblaPWG1cJr5AIQNSFOvnBJ3
hgp/Y6k3sGkqWa6eSDu7HAOKkyWA2oUfcrBugWspLGAwx6i2ncgkf1kBCJh4sIDf6klSQOEOI63r
/vPFrG02RWUwr1eSLjE023wK4YP+qEEVbDqSX5eLrPbJqc9brkzG4vKxcvIDduJVLjWUfcQrFl6t
hjqy2AZwdLnDWj+9ali0lF0wNZaQ7MmpZoZLOD2r8aMyZqLxvn81SNZTOHN7Pf2zRzB8I0p3l1vU
X8jLg9zDGxvwPAxKWH/Zz2//cLDg/eZefbA/DCiUDjJI+XiLSPRsoZfDC49uWbPYaGDtu1RYgZ+R
SqMZN00POt1DJARDYgorJsPEHcSlzQIUrKEqHEndx/MrlXOb0PLUy64gOuztJqfKjKJVEgWSzjlK
8itepSA216ibevDQbdQM9Me/o4atTVaewrSXL87Zf788e1fBW3iNBy10Fl4/W5XR4q+nKno0U51F
eOJTVoW79IP4APhz4bVHvelQEWjUxto0+LgvErSgAMdCpIs4i/FTrcOsWZfnupxF7xY9HcqzFUJW
QJSmTQcRRjJEHyjMl/gg/WanCNxUnYKEIveDR1b6TWDW1z3Q0jGxcH8QlDY+b3JOjFwe0/tZ0wDI
xkgd/ukY2283P9WvQldD0rFfkaY0/82Svq3r/EONkvW3m96mJpOu7mlsg47sU3y7dXnAFzxZ3icd
xWzIq2+TMk4QzOFj3S37KVCN2wiXI782Xo6NTARyzeLX01HbepTX9HVlFoFrKzbUU3PnyCxx80DV
H89sSMZBAPY7MuEq9+MXQkfw/Kc9aCNZC8Elod8ilZcsSuB9SNbG6Ji9ShyM1QpKtSsYG8TimFww
NTv+fna+/ezIMhGm7C2EpaRevi7vLoEZ5mqZu+HAx6agjR5DcBPo8G36IPRVrK6ENbpjoPaDEXwP
Fsn+/pSIJtnCfgWp3nCQ9Rs4lmxIKv5O/U3cYhqLEBx8ppnXqmCxwPm1qHG61qtSRyijjvOoGzq7
VuxzdEky09HgKipkvcfSUZczxhb/Zsv9uVgIUKxEwjOrNUzybfK8KIx6CRmvDb9bq9Zzbb0iaEd7
1W79TfBaVcPAqId3PegGA6w+YNkhxXPrWkxqUB/mM6ZLDlfYWT6JFXniFKL7vErycNs7zfEIE2q9
b22bDsB26KdH2cgOGPCi+ZqAVduHqZrEJB3yrqjldleBFnHzxHJ7hERsO5T6A3C7iAt2Yo5Unuyr
1ujfdharzENymwHXWOAkfGRQGLrdYJDge4DOSVwy6UXXsZSy2DAjbaeBmdR5Lkk/diOxiYOsg0SF
XjAixGwmaT3sIgTnlbE2kEw7VVC2J3f/HkQK/1HMOueMCFuD6ypkrp0D5yH25U/4sq4A+7v+Ahal
4ZAqj4R+349EmgYmPwkfoVp8IBcDWIrSlMFCY5M5O07GAXNeQGWdEZvlWji+nanfwJjQVeUfrpin
r0EQ8b4mnUjBb7pxLqiOp38XVCa0n604rw6Zh7MqCM/CRyx5wID9GnFWVo1eTeyy18MPh54wXySZ
kMs0WgjZEbDgIDw21unCAC+YO/0+GPnQ/t3Ssdf20gESoX5hsSpJi00lh6wkNAw8yuNAXUq4PEJ0
Fma8FELH0bsM+vVYJM8Pzf+ob26+aBkeugHiVUsJcOqEkZ9dzn0QOEg3i8H2LiSullzcm5D3XS39
DBG5EL73EfAa4acZ75xke3Vkiu2YkKDQGYDDVo7+Z+X+r9XuRPx0BqyNEqH8EGtThBx9Ied1+t6d
O8u8C0xUeMV1KGsP3fKSjtqeAn2hGfr1ySNQ3Pv9RH31rdfqi7GXNtqy9LYUtaOrQv/TJOFDX9Es
XxqTtp8LiTricPcLjrYCRdINIRRZYNVR4YkOkdy/1XZG1nYrj6JMrdZjQK5Gwb77JxMJuQ6gcvNH
2dNK8vvYm4clFhCR36cvva+lQeeSBXpulWG643WJe+8vKImav5jtMBnE1lfFz8dPhuQCiAdhCGHB
kA22YzAikmNH6O+1LWi0fMyxbJvoKP4E6Tguv5l3bctPizZqx52qssVY/nf7lLgqNiR4FwuHXlN8
X27daEa3oySzTNB8nz9ZOur0lcP3cjn1TaKEaRslMiyxrTYwCSGdQ+9ryxxOEaRExni/BaSvzZKa
gOX2ndgQbEbmU1oQ7lkQicDm4RsDQUV9aJPxFEWPTFhIdaiF1bTtxLOzzVjb9u8BZpy/LS7r0vT2
dvcYjrhJkYvUAgsBAn85O5wXFt24fQLejwNoMdciST7R2lVbqMy5a7vD7ghI28/Bufo0y3aW8e/E
GlKh0k/3s6xzuv7bKmioKcvWN/UfimSTDK60uQbt2uHCq0lJqTJjB8ww1rWf++h7VOSOdQVKZV0a
q2ilb2XzPAynMxeXh2mf65qUH/UrrtLtTOpObA/TYz0c1YvxFrccZa5CEhAsUWlhyDR6Dm7tsYMO
tw4MykPwDhKSlpxaQZZXbdWZA6SCHpvPhUvwfuSE182cEZRWIyN4aqmn3Ko4aQaUO6PSOVuPg0Cq
2PLC+4y6NBlxBKNo+ihV4AgXGt1LsBbIMccFCUnYyLn3iHH1QwFH1npB82+1bY+cnT9W819QXLff
Bt1sFqo6Iq8ubQmSbi4tAFDEb9i+7WhqYuRqCT8GL3n9vlZv65WuLzTNTk618W6226xAdzdw5Sxh
Z7TSN+zpQg105dmm6LqxgmeNisFijYaXg1AGVve51p+7Z8mgqTzW/ZjA2KP2DYwsFqIG1czL+NjK
H8unq9JM0WynhS7Pc3/SYW9LRsEQEBIypv2DlcLon7s6Th5NFIdejej+uZNv0pYQGSvZC1t0ID5r
C6K+R2AyBhdPl2DVlAlbTpPP4wHvhy2mMiMOeYez4s5nyg5dZAhXnDo8glvWMO6ugc4B693wGehm
94Dw+MIYsysnXPzI3SfDr5vgf8ozVkLuCMwTJXApHaT6eICambjDNnooac7qAe44PCYcxlbjDu6D
dkJL/2F9f2tlSDk9k36DrpXYlcS1BInal6GYDDy6bK1cfLhI790oXQVbSEv5U2oowJ5lsg2AVZcF
9agJUtvPtPN9QAb0vsZ3AIkKsLunLYFuLrEB9JIfqF+HDGL/5vxBfdQXp0G+jhCU+LQXvU2/uBPN
N9Ker0RGHsN7JXMmbw7ZWNqKySJVXtQwAgaURzM0Fqr+LMBNnCTUPIVGD/1DX9wdinRZsEsoUtCZ
w0J15fK2v2BjTCKuFUwAz9nU62M1Vb0ht6YaIBs6KEddCPaqnINvY8xgnexB3LrkzJ1BOsEaKzD8
pduZ/XwiepbgZYW2CTA+Y+PTRXJpuArKz2Q42BGgANs9p5tx5IWvVYEoNsiGjN/w/yvAzUWyEXNP
ZFuEBjofHRPOUkQB1CnFUfLWJkBd70g3+Dqx6zn/caogWP4jnjbA4iJ/FzSUWCPZZnGuuSlioicx
t6a9IjKFZp6TGvpWpvc0ToC25ZC+LmJvRv3EhrLxspsI9z+998tOd1stqVBZGIBQsGrbsCLcsO2a
PrtInTwJWq8yj0tMq4lbv6GUsRV8ifzC6h5xUl8JY1agXAZ9H4X/pR9kT0AGwQxBw1bmPtw8aDsU
ne54cFlgPUC84sN49boxEQC5BCoa2MONedolGbLCnhBZHyqph8Y5+sDrODLim/CSQy/QvDmyU4vG
GqJBzc35lYYtIdOQDM/Mg2vqChOJLCXE1ODJKFNnRayiuXfDrjon6FLy17YVgHdYhZpdSuqdja5n
Svg7qaWrWcyJqSXz0K00R82TRrLn+kE69yeCnYfU0sF0pJ0fIg4ec9x3EBKP4TtikAG/5cHjPMwN
w131SUwtOfkbX24xSvytcZ9qPxqszFURDuzCxIqm6sgDFze0hPEo/BbbYsnMetDfBtdySngAs/aa
zSoD4lBkAx7N/RLNWJrhky3Bid+BBEgqo19RhzA3bWzcV0g7eydHbcHwK1w/UUVs3Vp1hgsu00xH
02LoU+gngH4bRbAAsN1u2/UCQ1uT+VFwe+Kt1nV+aQm9BICd+pabypouh50tR0OiAflZlEE0+8ha
WGW5XvHuyghUyS4EgmlVkPeHyvEQf7kdu6SMovgTelFi71xResWwGSPL6yp4ur2zrKjID15TGvEE
Mbu339qXJ38NPkZGXfsOXx48zkcezUf+FO38DVjRqcdfX76N9XTnczKIvshSYhHZkVI+j9NZvsNn
6WCeWprRZ/rG5Nqpsw0EanLNXFDZEoK/6NFDVsAnU7c//KOzo92A6+hkotpv+YjrLXeXX2f8ibmn
FY4orNQ7dfETAglhx8V1BLSvh4IrOiDbwD6qIQ8gzi7MwYBs2vGVjY9CpVdyd5tW2esbJt2bBJpM
2R1bVkFNc/qWEl+OORPmMfALXdaeRE3zxBYUPLBk6sPZHIy/VX0mKJNcGh7f8QNoCXAsWLlX4IUK
xWfKfx9b1uNNW56JBkFi3y5XiIDHBd63XxlrRMmkVJwAmHvpuhpGorswJSTUbOm9iLRXewVouZvB
8lGyEx9ldH3edhzLAJTex80Xd1NkLo/aCzdI5ajW2Qdt5H6k9haizxFD84HEZdiKzLCeykuyACBn
RfZZ6rXDxO43iN/jBSoNvHJJpB5xVy/VX3Rahw4+2n6gcFV50pK4HmvWIkndNg50H/yoo+gv74D/
pc0EPDxaMsFORSnSaNcU2/WZC46YDALCXWXakRmhqrFktyj9hC3fIGji7GZplnMa9gVZdZoaPS/8
9/gDl/KgVwRqt5lCfIulhbize9XdVnvGFs8+ZzH/By2Gm/e5SmFC1fLJa6L+iA+rvE/QwNp6B5Wq
yH3mJFPSaYiOCisVw7Li/87cq+lMW8YWSBUh/kfxgU0aRV0dlA2HREJ58mEDvCMZ/RRw/wx+1OQn
z6iYYfie2vWscV7kNeFO6dpjRoAKLeFrvqZymGPdDQWTNuYh6xHS3mHWorR8uJ3+0RYw3uTnx2Fe
6S+jk9NVHG24hsUqzup7svL4hYmLxWeFYkpjSDrDAqWTQoo+XQ4+X99n2jlV4zkm793LWwECR+io
2JFP8JBaMW5i+0KgE9jaw81FHaspIYm7SLPrFPY9tA/F/lzOj6P0o0ik8/9o2sOS/naqtuP8eHdY
+BqX54EsOdO17SXGU2H1zDQvVa5kpHm+z1mFRC2nTSxGEz8ClfJIqYkkrAGoTwSLUSFjXiB6yFt1
uK17f8rtDzmDj2Qv7pnnRUbQbnuCYN10dS3oeyvaseYRJg8AFTBs5k7aykoRt3ds+55m7u4mpQzR
xsVm4pperFQUhvDh4UaChrz/gbSm2exZNGUh3FV3s+ZxH1nekwJ9YQCrQ3DVVMPN7VHGns+0+DIy
anI1apfLxT6WswU88xCdw1Kpha0naARzuwW8bQlrsUJT8z3R1Mswg8fIRrWmZNzj+i3x4XWeEzNo
ZKFzscmYlUb+Ksa7f7gQUG0sRyT5NwmynI+xf4yMVjeq4SzyEr1IqM2Ga+M6X/Z4rAwuLQx/BBmI
yyPoSlKZ3HEkqdMizRUmBN2xjuVxXWbtBrEVoBf2bP/RR6tBoH6mDH7HbW3ErzHmCFd5CvbkH+Hk
lyfzncnoHYFpRyaYgnuoKfbEZSqVJs4qHofWL3ZW3VhOF5wV6LoWqXXEvIM7KyrgmKG5guyLRLz5
zuEJcO4FG1085Y1wYTZ4i3WdSYk+lMdeaekGMTsGgdlf7L386Q5mjOELvvjJcXqETNzyP4dhvle0
tSK9DhFCue+FloZoLAequHvjFmxvYd02OYut5+Y6iSqQDXV4F0ec3xrB3Nm9GoaVW3xUe2enS54b
hzEzs9oPj8ylz4ylzhPf1GNBcIl/SrYSj3dz6jChqRw7g4JF6brTvFrOSx1Msqk4XTEogv7Ma3Le
skXt+/QfcixJ/kn6795uLXE4tkL+RqLp6ivLyyP0uS4APFerKqgfyTTmlPeM8Ul0NjfmfuCUSykc
Qc6zsywKTHeQlwwhuVplEQzVObVNN5cQhjLcnd3LCb0BIHrK3wlnZjanFspmw1BfiD0JjE4Z5dVz
2BhLUaNzSfO/qDL6NtvHBTGJ543rcbdAifba6hBPpoS3nUyb1G5T847f4GueOPKx0D65vYXyNxFj
UmUMzTFpF/DrJSsmVNV8YjbkiVKg5r7DvWdd0HXeiL5Dt/GBex5D16J+od73p3sx7D+1NicajpNp
zBQUj8Gxq6UNWdrqJoArCu8OzCJWs+FBJ/ci/pA2JuTJyvxYgoqhXfPabCc+3uirxvlBeXmkQYw4
dZqJ6/Vq2gizdGS6+/udY4AssaI8vax0KW8HzSLSBONb7GuKMISa+u5M+b7Tr9NMqqLkR69JrHWR
IUiYphGUBNSfbBzjUgQ1IPEdtA96X2RHaWsPmkjzn8Nh0zqWnNv1RT73EhaD9tzRA48wV/mZtkAn
GVq2A53A8u9LVbvCo3lAi+tlCJ89Zv8CCziBAv+EkbOFjwcKZcb4cXn9aqnCeYtsMEbuwFsnwB1k
z4Ofu2UK8A8L+eSdQAUezLtfqyyzxGnY/auFRZBtSCb9KI70R5LY4HhTKhjFO8SOHxG893PKoL7+
jgFIvejLUFBi0Uy9ucSh2+QmVMAfJO5K2VTWJYMRl5+mpAmx36U4FMCfvcLuMofKEk/1CeJ+PgBm
H4SoZVvNx+ugy/YAJtOb70hw3vOLVe1aRepMncbEDnMBaE1uK/mnhbdzo45ejiKJs69iTtVrZVC7
rtw6zt+cmvW6z/kpDi4NlW3NtTMxvEXVUvDJpg9No9t302YOvn/pEHerG4K3D0far8re3H8MRDsD
V5CD9jDj7iv31apsURnRObjMFGzY0sfufFr8snmMvDuawyFbpPtkNwJXeGIUJBQ+ifnN+VlfXRiS
sSJBagAoM/f8RrypZLqHEJkztDwcJD4cI7j7b+CpjN9w7L6+GPQmSoCOL6Qg/HNUu3Q60WkVwho4
YIev+Kz0wrm7DwcP39dJwckqNKOA7OTQe/bkAXmKy3qxHETE1UjTyJ1b5yuIe33U9t9Pm6L/6jPt
W4C5k/DQsvNKfJerQESF5C67Pilr516RlsclhnxQrZzJww2Vu0Bwkb3xZqtxMgEd4YweSEn4IonD
5V3vDWfDTdxljIouC2k9431iXI10URZJvOE8nColvBVNQUuDnpuRLQl8GIG1bM6k3xdXMudrMMmS
d8xzGtU/2M3mACLB1sL1fiLXTmUT7uXdRy1p30kelmw+Wuf0/6TA00nsg1bbTSjKh4XIL1mSWQN8
+0R4j1o0MOaXvNnrVI0QaIPjR5qE9I6mgUu6UYjeouxUgyC3+SY3SrSl51oyB0v3xybSVaOlvka3
V5r3wD/BeRA0N1/HVvBSTctvx9O+6ijz0KGjk59VRaqMi573Nf6/6qMMeFZK0XvqGf7l++V51Z++
Ofycv6YYeWYL1Op/wMTy9OKmsCXhDzDO5MqhHGEmBJmpLL31ArJMx3ZguoTgECqRL1al+G+CGE8u
3sTbu54GlTffPXerSO0/aTL+s79RNl7SJ7s2FG+e3ojmo+xdGpHSeu6NGRiplCIOPaENy/i7W2lF
07AxO0Rqhpqn9Xz1ckvUXgyCjqPsTgxecCcK81lgxa0rPIdbPc3LIXCJfAivut+dmcd5Qi3bbNvS
UB0+WS2r1KCkvTaClc+AKpnLtT90BkJLnIydW8BM6M+xeEdjkStfSBCaYI7/VA6F6Fsj+JiTcPaH
p3A6jIryaa0l6+rY3PYv80sF53h/cnNe159nU648YrETpZSuTTfIRAmedGONHO1zWMTGC28u/f+d
0xdnfLer+ZhqcsFzJHH/EqlkwBE+bLd0OolmVqHGcVDGhyhfcn7F24Fg2hlfSqCOBKXBwHKib5D7
xUOhBIEauXK4F5G2ZDsGvBKNVkQ6RH29VFDZhVVQNlt38xQuZk9fpd9k2jYlFVc6GLdyfNLsxl+p
9sGKd+86Gt0e1i5Gl9bneAOXlW9X4d/3cAVUm6sEreVkFfTUa++rsylnF1QsBvD+9/FVVZyILpMR
h5cD9wv37wC9QiR3vtgQmaYbr+aPC61kPEauM4yiLCYtiO9ZoZ3qQC/MRYGvPtxyFGxl5z3BCjat
IbMNV5/dvaHRydQ7cBDgMoghDk2vceZtygQoCOFQVJthJ+HtX3XgDnfS2wOgwp+ElngjPa3UAp8N
+3JVj4W9oOhE8ejnBZdLhV7xLWcXgnvBPZMoBZzxEXfSG12iMuT15AGQvnsWqonU3xApjF744l87
rlQm/IVWJA8TvV+pwDFsYFNbIgvTjBPtsZEAukMeVsuZY2OK4YTH+WZ7onW0lq+KP8MGzdbhRogy
qYnO/zpu+SuwobcJXUvb+i82PFRNh6LV1edHap476vBGAFJPqn1hQwWryXKQyCXfKlUwMmE2vPJU
kA8R5VKyCSx9jchXFJ2myTaRFaD+MWbIY1dzYdM7Uu3mSwS0U3FKNbxRwz6QfYqqlmUvcVpDC2bK
/jYIamgR1l6Pd2V6RgRlB3kAZXMDmhAF2IQBgiyKu5BqodD9f/EIYm9L9cnnWlI+jbsKch3DX0Sy
4ugtbCPUvqHxZejr4UP6f31kESUlt6SPufkLa30h4wx7rkL4hVqJP0nrUBDP4NT7e3vhUV9va317
HvREMX6mSu0s/HWBzDaMPaYMlZONjpwGj64eKCVryykJaZQPEPVmyN4zStgagu2PBPq/9YJABqvK
fPRNmWViseHDHYKH8xqpc/hX5UtAjjNxZVYA4p0c7riq1bwU2gyrpp0/IfOIetu9v9smTt0RZPsw
bsyzsifIbsC2ccBs2oBUFVR03wilNWeL+jJFA2zXgR0OFoZDpeL36V+icMxir+2MjxSpW9gG2wlN
R2jt2icnqBYc3PbPdev4XAtXju/LS020MTZ0MO+v+GfXwH+kWH5UdsGBQk8tMTCkAHyr1KHZRUxJ
40ZabLiBwG0GiPYNjmJoGLluNsTkpikF7Nq3wah9aEg/yKct0fbaE7zkSGRSmBA51n00WZ0rQu30
rYLlbxZegF67fvX8FscGMLpyELZENMfCAq1einOdWZdugvHBG9mtlBG/BnDqSOnTs85m0md9zHd0
kcPN9bXnK6WocWgRdlLZED+zE0FtBVc+dFUv5tkSszrR/1RPOZ33l8apgOX7eXrPBWsGxQYhfqEn
AYoCanPcJ38+Jv4HHuG/Not4W1EDdxa6QNvOPT93Snx3i46BUHq+xCXq+3GJ7jmQT/ptav3pOjD+
Nhj4sXKcnDwvwbYQKlaaOGGgn4r4HQSoTUtsmjRxuS6sl/C1GgGyCmAHt+BrC+yGNPYYQ7BibUPG
08yh4U2ym26A22TgeVqqYLi/NFaDzC7crkSZD+kG3pMB/qHPwGiqFkQmg85miOW9jI0mxQS0VsYi
x5uWHBq8HL20TpoQwDS/uyhJuDKv+hcL/g5vRNohGSg/YoyQzuWqYcZ6akPDc/QowD1F6w8GmI0n
9Y3H4UVQZTDXHWLkxWvrx/v4Z8dPv4Q/8g6OhCCekEJDHJ20OSMVx/2P4a3pfDn65EZPCxG48mhF
kG9cyoPAsKp6HnQHday2YKV2l/tPIo8MWfb8TkguyryH+J8krYUL0dQ77YnsPwvokPVFai0YXbfC
MmXb/dh/BUb3egwtcUSgpPV/bN167Gsx89kgp/9RqX7zOCvggQQrAzzpDCghtFz2j0nChPk2sVd6
C2NtAFwT9plLj8VmG6qxnojRvR7dWGBEoPuH74fgYaxQb2qb1eGCBkrhMVVytJwsGKWzdLjZ9TYb
stHdUZvtUyyKrcUmFSch0vIX++EwW0wQKFql4BMr2ZToIh53koiy+5SBci7wB97u9xpmzPsjElaC
t254UCEaml47c/uZiaVW944jBrIpmdQ17mjhmdk2SCG7XeAi8v5XpXGaGfZFgZzSq58ECGio7XxP
s/8o/vP7jF32WLpPh4ISmW4eGMyoDsQvvikByud+3jTie9QSM7ZzKENloi9v4y24MnHLB5tfEDsI
maB42kx5JjanL95d5i8KfTVJkY2NG/k4vt0kn0pygeKnmyThhXsvoSXEKAKPWOc27mhsMgVKYc8a
OzQS9ijH0g/efMY4KECwdZtw9mths3jHSnZIi7ygNui2d0tyOgo7VbLEBIgOEpVwt7A95ofiFywy
81geBi5mzhXXw6UOWxluQx3k3qEiSmzElJJF0pOsXDkTIcpU0/NW728QKT/FQthG++Su4J1Uivgy
IcewqGrq33GgGke9g/xT70ziFJAbhDN8pwl7wQRDuTp6ozOyRU5KUI/uHfsD7479pgKCHDJZsrid
MxEbfOWBSogBEiHjqwVD2V2c1/w1ZqXNIqqed+Iqfoxp77z99NuWyw9vMfwLBPCR6aQu3vC5o28f
+WKARbpqk6bJ91Vd4MzZ0bNuN1d+h7cnampmINWet8C6myiCz7offV1V1VcpuZXoSbdxtGtuhqU/
ebLCIqnsekjJ0X4ZvdB2VlH2h2KeoG2PmxeUiiSFmsQnmPMqxiq77p/Z0nYZY8qhOi1qF4GDxEMX
bPfKfnq4S9ssIyjD0AN5ZhzQs3BHNjZ0AnUVf4+fEhXRTeWO1MPFlKlq9IX5qdUPawQyBU24adku
T2rDj57Go7mNSf5cT9m3brj9GL5nu4RNhDTkSYw61mIQHtnfWbDAVLYdQTu932PeOSmEdubOC9B2
Xsl/guscj0fb0N3dzdui+j71NQcuOz7pqsalXPZYV7Riu8RTPCVjfwdfirbasiKwLFAPJc//AG8d
BILsmTOxdXOxya0kdDB02aejxyxDSWAyhR6n5pY7n2tTfHe0vVRyAgntRt8zSVY08YMR1dbIfXWT
guDzju7laohpsCznCi/2uiY1noKfeJ+vjJonR51tLAygtieB6yuqGEk8yGDkNXFwqzEVtS2L2Wra
iJIv1CrF92cFNzenTkjXbmAo78jlUjPLaFLv+EnEQ5axXZKR7jihDLU6d94EUzuvQsOtMp58vFzs
OALX2nk+oPQge6rs0bjdFNnna8l/gSmN2lNzURRNa6Kp/Gc7+M9pS5nFTk7zxGHSf+d8979zQUpi
RKJdNDD0z4gOMpw3e9ILTJ4C4kTHED5QPoK7UfCQmi6KJ+3dc/8WJUkmdEz6AqAcMrsG6lbDRnSB
ALFviFVDo+9mOVPJEOvD8by40yCJLKfa+vL3BpluC0qQjyVmvHLbmPl4FCmtv6zq2Fsks7ivY2LQ
+fX9RthplhS+7HOTdOksTlqqpjZuKVhG6U23WQL2KJgaA+GRqflYP2hfl41x2NQdV3SjbNzlMENw
YG11LA9ENA0ZUuPIEkKpeXoXUSVCzV9pT+vAeCAzRDjIGK/xb1apGqp1AoAtwxeoutRLIk3Mupex
FpevNJAgu0VfjzFz3mLXKN/YaUhJaHgIy5rsKzmZwH2ZMlCgI357c65wb3geQcq/R0hJVDzy1PKt
XpLCKqituD+4mgeYjyJ0Wr1nv5TdSdflJT7FrhkLLq7VdbHalLtzXvZkkVVBS7CWeOj+DPBM9MXH
EyEyuD3/4yNZIFS77BjtOcw9L7CPvLeqQHtMk4BZMtLXqLgLtb0vCMriBPHO6QGqsl2yCrJbl2Zx
JmKhEDUGLGzyodJpMae/h5+VuJCzwFZ7ynj0PM6PwMtZrSgMjFv98YWfs9qgd4RwYmJEF8fxdDhL
p3elTEhiLcEieWLxWDil2fqmJiPZSuMAhfDSCqH/nb3nBsQN3uaAhE9g0FosRjBIfXQy55w32HHP
1XNi7iq2y9N3TQS0V0bmVAYGq1Pdqle+b5XDGHXecRY5JxTG+0mxrjxk+EAN39pwpbfh56lCKvH1
WOi3v6xaIyVKQ51tJu5ZVEAFz7TsNZZBlfJ/ayDBGJTd08mEZw2aewRTWRxoiZYr9FLawIjk9MV1
F/xXC81MdlM1N4wiO5GRvk2yhmLntdKzMssCgpH+aTym089fh/81f2ECT9/X+bXOWEqPJ7cbSAor
FKCPgBEBkJzv0tCyi37Hr3+2YtUKcO/WrJYi+0rVfiZCRzxt5icM1zvzsYXojitmRbEgTvR1l73f
dmYmIiK88jhhpcHPHj4T/Lcae4kqbeXu3Cv6czBk7+EgrFkqV5aInPC31WtjRnDpeNfg89jAzA5c
IT3C4ATI9BxaSXYD/25tWPvTaWoXd+6w9nRC0R6OBNftPCueX9g0+s1u45WJ4ZhWrMviEhEA0k/K
1KHC4PIXSsp7u693+z8qwEDLJpMokOdI8ibQt4CbxAfW0VNJl0GBj+/NjZ+i30v4oYp377Gc16B2
19z3TP5QzUkn2lzfHWiqk2h69IBji3Bc6CygOGw6P/RKlBCSzSUNGaDx0VhjK7tavG7oNliPoo6n
qJ75Ovr4MVTFfa3eBFeLD3tSROkp5DKELlTHsgANkvtMlv5VIvro1u39hQz3flWm7ELf/fYxsUc8
3gE5Sjk8pLZSXzAFtYakCtzQ9EgLybHjxQnOj7wk4iLjpRr8PyqSUfI9r860x9K/nIQ0/qZmZQRK
+vyZ+9n9AEm/UDUA80vP5v1haM9BwQdDeT1MD6+Ryg566mHdmNK1Kku3GhfcUTRDqOeLNy4haanz
14A/HQGJ46rkdfi88TeUx/iRs5+Om3VVFVEOkyHHZyyqN/BT1v6RoziQdnA/gGftA5SHaPim/uym
rnOpIkyCcqaJ1pwmsjJRwvkWUzoaMHdECF0R22Dp7RbM1GyXLqbvDrBl88wO30NHqdmdhrTgsuUN
1OoHeQisN2rmm4BY71+RWlBZ4lWVuClkCZRd6i3Np8yzoBG0PvsPqOI38kgibB/hlMGsZ8tRTTtl
9xT5g04iror7Nk+Pl0eijrpRRRj7UXdlf5nsXHTFcBWAvmHG1pxrnPQ1K5fBHA09BY63oHDFYVcA
XFJsIKPZSMP5ct8s5NhT8m7gHciV8F3hErOX61IwbajuznKa/ha7LX7d6BNXWNN36DZI6aZGLkTB
+CcgCmSqNbINRRGua/gcr07jyfKvJYlq8NiJiexJL38ImBbiXIuhyo1xuZuZ7OYWu3oLb+qZfMUU
FoZbSLFvCWu/FwpI0xh8aqWxoZZFRubZLfhi5Whnt06nX5AS2Kysf/Iyg2YSwkFbp/kBztDnWqml
yTM0qugdgnq15xdxKjhcq6IZZrxkJLjZCmsJecRbnyXYh17rNUcPIX67SPni7QDr2PB9NwkTiPay
cfZa9CNeODpepVaCReiYKyKgD2QOQ/KsM4jm7AMsIGwKQNShX0jzgu6cSm87KYuxDpRKH8k6j2Rl
Y/8l8COU5C04pv352nHliP5A0fjuKOiDhOJhZwYeZee4WJ8Wm0Ail9ppRXwbDAxWng5agSy5YAOO
FKXVfwPVIru4xwTDGzmR/9MmyRhB4ZuqvbLJcg7iAmZ1J9SAuxFZiQDOEKdiWWMusdFiRux1gYK3
lj9x2hOiQYgXGv6vk3tUaKqznpcouNKEAQkfU2ukGUYO/CGXW7fCtKuPCk8+2PfX/hiB93d0qQyk
nmHuonLEKTBQH8DUhMV+7gpB6MJD2nPzifZawqhGtk3vJdEnnISAMsdL0sdBRkNucEVDaxYlaI6U
ZsYiFZiC1gwaIhnDFIhW9RvkwI7F2cXRg9yDUn3z+8dFCVTAo6UaxTRgAJpRL8riRbu/WcMS/foq
lI2WbDL+0ZBw8hI7G9NqYnqRQ//E6Hlf9FCmu46WEYXncKgWnjs9EzT6tfd41na6NCKjGSwJFrp6
6vT2LX10eSquq+1ICvTxhbbuXmasHxr5bN3ms4dtqPvkvWa3IzRyi5CVaylj31RMjj2N38ZeLu+P
sjnjto1owqCzLIX0p5Vrm/h54IfTNkMWNatrSMijEbKMPtXtogfBVNt1cUVniiqM6fKFqOOQWfUt
KHwGp9Yv5egNDIxGPl7XEZBq8hgKFxmWHjuEK3ulrdz1iclpyxLQIBfikh2SKNngj3ongSJrY/jX
557S3fEDwuKj1nkjk2lv6mBLXhqAlGrp2BYMGvjqBcax5MkqHTBiUzJKMh5av+Lwy4KvpKeViihs
QLMjQYTWVHKiPALy0+WJhaZFCACgV54gjjjDzoGXVPqqr2RwO3EFPFaZ0a/QVeZK9okVGKxUUy9a
Awyyt+Zdyrz5e17IS6ygZd2PQxTFBjQwvv74AXr3kMcgsMLfkUQGG38uo+Hh1oyUue5HUzippR+s
442yZA4uEWsIAh+DHPk1TewA0MqkMNZhqWPLzg46JuznQSlDaNsGc+ezP1dlGsQGN4ldedRPrPWD
ib40KTwmxlHJsiq8LJLsFW1/S/CXolPc8dy3vEFvPg9/PYyMTR0CNheDqnDLSBHJ35bR+tRgDcQY
6geMnmoFRDpjk5GQNxjpVL3lDfI8OrSTe/bubeRDZAUlzW3GTvOkgMiMt3d4cnGb+PS/BCsbzNqs
b0DISlUxhK0qwIZ6URDydzlY1lyu8x9i5W1BBB4UChKFRSBHy/tg/9Bor5cinFTEIReXTtyGtgkJ
gDc4I9mZg9i0Fktji1DwXz90dSP3JLTxRSr36VTR2680GkONgNatqSgHxBxnzpGb0dGH9wEVvG75
NuWJTJi5EsOOcfUfxH3mLh8sD6+NGqYUWL66Sz0mcIhNd7yJeJpCOADpPs8zG1lcUfarHWb3LH99
y71MlafNwjMTuSAtDo13D/NECleXonTDpReCPiuBPDO9UzJKciLlenz/oRmqB1486w3RE08YaMU7
83UHFfUOFH/kQZZ9YGWXAEP97p8TuWXbZEBzrazM+USV/y4z+37ffw2jiOE0229FmMsdv4r/fEJV
4kvUCrNA6VCntEgQ+PmEOKZ8+e0tm4jeGtNJMderti6sD+RYaowXxZzRocBeT7tlvpYKGXqsZ4iK
ETL6+AUMaPwLlClaSW1NWcsMoFwPM6wdCxsPpsQpRF+a+QA0poEGpHAszrwRc2ABX0pQ/Xg2ew8c
8cpM95/g2g02kEiPkLeFyh/meYV3a0A+CRtqvp3nYclj/B6i6p8BmaHELRCuLPs6cg0hzq3w3rto
zty7DuOmvVVKP6/2XQ13kCVJB05qKLBG1eP1Rye8+Ozi5H70/C5hYIQPa/BpUa0gTI1Jim1ol1O8
NE7HrKcKtp1nTSBDpP2u44lPqECWWdxEV8P3O7jTm6l1JlyF8G8VgEu1KbU8zeb3Q+K8Rv70WdUh
pWfeMOprMDB782yosbQM+UpgO8dENi123TcGI8wtCeuw3zKBA/p8OuILJVxNjEBt8Si+vIpD6KOP
5WRk5iJl9/tRyHXDaoc6zSzYoDQarNQ5xUJbqomUMMmUp2N8jpLwmhv7l7mfSFJ6RHacTuyHoUcd
ogfUxzLWfokuKi75F5nh+Fk+2OpvM5vzroE69AUt82tCpGA8RQVIJubD/XrvR9U1IRIu1hhjzSig
CnFWgAV3k6jM/NwYUKSRsJqatYbSqd7iSa4dPVMeWy/8GQ/W38IRkB+LFoP0PR7G3RnwsbQ2LPIG
dal/gaCanEHnx1f0I3iaAGb4O8AjvV2sg9Chqk0qUuxqvVoVlmQPglne8wLGOKbzZTQ4Ivqpq95q
k+WtNSS2RzKa9Y+eTUlxgZAC0kHnBYVJSyzP2IniYZXQddIAg/EGVHlMfxfVsp+qXShGyTc3OETS
thsrf5MyEMk+wdEC2mdjnM6pnLQ7cMpJ8y5hxC2khlGzK3i6AjO75fhzGLEpKMnilvFCxbVE5i5B
ObYiGMOQpZmocjil1r/VAPI+xG7RyLbkcfug6B/CUITgOMSpChNPMiOmPXubrmV34rfu/B69bfLA
DWS+g+BQmxnzAaknTZ+I8ddfmPhOKT7e8b2XzUeQ4bM7pYQxUiXeWjVKoPprzUfeqms1vG76p1hZ
flVWeqOzb7/KfbB58Ig7LJdFucm0VfyJ3hyrDkZry03i6kbk2nGTewjZwDhagHkzvVWKyKCuXm+y
RJVYswXZy0gK91OyONBKXlpPy7EbF93UfKRBYY5vZLtvi6AAIOrfdnf6Iuzs3nQSF0uAyJwAsxLo
XhWLNYVfRyhduSedyqGC5rCQLbfEwIBez0ONPN41iUGzb69WxaB6bLdMrFSVYGR9WeWX3ZgjRpfE
c8C1bh6pqClIvac2YKPCrmpSDmr85tsaZ3OoDFYPBUK+LZPB5vwb/r/ZJDSN8GgGmzrTAOR1BoN6
QXhC4PCf2F25WNvbnvO5mNdRBWYUfHnYNVuZJbF9MUrI5PqW9vsRatXyb+D4JugolJi+BGvmSCmA
PsB3n9u/M90hXzxIrgzeKIgBDk29SuTfEdlqQgiJdWHdcu1UkeFQzFiu8xakKzL6egQ6K51PJ7qz
U4gcCg/DXj29Jw1Th47O51WLdqO5rSwqCALhdqWnUWTP+cz0U1JhpCPPSracmy4r3jBUERWijfML
A62dMsqZkSydU32EJ5ddv/JItJ63hjOB15hd9eqYK23zMihWulwJv6WIqIxKSB4l//mduI2x73ga
qnTIgvdqIhEtHstfTheWzXbGM+WmEAwlzrAYCwsj4d1zkWME2WC2JqfAuQn/1mHhV/uJky1fXqFO
w5OwLckbPlY6CVOcxI9t1mDT9RxL6pelhDnO+wNpnd/IdYyHebCAbfVbzU/4pTPfnexhQXX7vIp/
fs/owz09Ujf5YNnyRHlfOm7SO/R3WT9fdh7WXZr3OjW/XyI0g8xP5Csyql+U5a3/f5wWV8uLKgF9
N0uLtiJj+Tb/U4eT1oQjvbDrpKKQRnvvR28UaCCm1GxKz6NOmA65UtSmVcpKsXNCgrOZPNpBZm/U
FtjHw5Hh/cNwl8H46EIgA3Hif/Q8gVvB1pIpkpBInLQuP4VLAM0N84/d+npZVL2VgiljvPDF5MDo
JydfWQeOt9xooVFTFaMOW8IVyOus01cPRoN4yrIy0chzokswuaokQPnvEYJNhoWyduDvLwBsm1A1
XINrCnwuPeVXX0GkWTCHdyfa2/D0bjId4ZruidSRlIJI73n7xgUb8qoFoUQxY75GDgD0Waivbhcu
FM1qCJ5CXt+psRtT+hKZRtDx9uvOtgTUrQVWt1QvGlQoSTZjXlyg7IQtObYuRTuJ15sC9Cuv5T7g
GHD0LcHNAtaHiOnULSOsLV/2p0BrQ3SC5CxAjDBbdmjqrVKf5vEizFpR3rLJR+000snguPF76BNX
YHwFnbeEo2aQXVsqwB3nTU2/D2xgj55vsXqO06TnZ/1a3TOoCXlMyJ+r66JVEDvG4cSfPnXQrOLJ
FV0bxLHiL4pCa4NN8A1wrIUPSgnfDmJNWlMeHZsSdzdGplx+mwMLyBG8GGKc9CVc5Y/k0cAH0hXV
vjA6EeMOeen7v3/l5Hq2dvoqkuRjJjqsoYutjnjjCeohu+FzWi8WyVzUp9AOBevp/T0HHUlj0TW2
+N8o92BFgWk67VNr2wvRb4PYrhRp/gnG0VkXhj2EUgg//ZmTP2AjgI1EUx+6ljhGIUnCuEanTbVZ
z5DczE9NIaluzpRaJkaNkx7ZSoIghOFDmEK/eyjlY9+Oqx45pzQvRLfw02edoLLb7Ev4YEsWZivx
Je2lT9HcFXDQ/9K2Nh4OWF12Qn4OdLB82L/EVga0V5jRAcQBrwRbSq9/filUTumXrN4dx4P0raMK
Eq9e4qk5jr79UCne8UuP5ZK0kGAjN28/HqJ9py6dxfbSZhC06gthANKISmuX3UAbh/Bou3SIBzg+
DhIoSfJ14aUC/D/JwxgRFs+LwZd9GVO0QH9xkDtEqXIXd+KlzZU38gONUoP/iEzfHs1hv1BvtiHE
plTOPSezrftkkOPIu3yCJzhEXejsS9XxFYOuyA68rHW9eYaxrcXJ4iJjKGbztCokmdV0SXIEpnMy
2DJaEq9uVrOD0RInX4tCKPQlixkAtG5p8YvYod0wYdSCeBYXx0Nqimeky7uHSEFACQc6TQ4s9CIU
tt+z/bupuMgt1FEU0z/wYrQI2NrGFgCOlhTw+HFFEbaTNG13qZiyrzdPgMxzfLdiyTbDee6Y5Gl5
VV0wi+gYF581327lD8IpnTud9t2rU46gaR5qZzhSHs/x4ekVsKyd3KWzZEWYOlijU4jqq/wwPAH2
UFvChKwFIssn/nDsLXDEGE0RPzaEv0/0robaqtPvUu4m1qQXEOp3zNoBaenNhTaLQLIVWDxKOZk4
UlJacWb8ZLLdYzVBggubDlFC4VWnSFTickr0y6iQmQzl8x55B2TJrnB1tflu/fMEfNQWXXVbISLX
Htez58a7cptxiEjpAHAVpJaK9pWA4n6zKypWdyDvwUR98hOntCGILAE+JWckBHvnrPwRQ8Xf7JUN
yjvUPZDbKw+BpBuQ270/uv2PDD9c4hq8H6Ecwq1NsZeVLwvjLtKIXnDdg8amEVYt1T6HjUr0jHhB
QFkqEbJ8kFvYcJ5CgY1+gn5WAYJe/+fKHjLITMRHwvQNQcP0IFzFU+x1kT0kHbZK8SCsTRF9Zdxz
D9rQmqhGM3MMeJeT+kqTUYzGx1A4HTfzIIwwA67K+3dGJly54ztPfXyXOnpFWdGOIuQSfO+lZZbW
L6PC9WkXDYvRjtfewwe77k26PlP2cPEtOR1jpkV6CRtHFg7PljPkfc+i9P/UhL11s2Of1GG+f/2W
WciSaP1u0TErRAHkHcJcFW17eSHeo+iAnAUphUY+EhzF2oGbjm060uWjZNAEgB5uGpE0/Y7S4vym
aZ9inkq/htyj8ff2JjxPW4Xw4SGbwInUkoIi+zgxagJvNhkbOU5+4TplnSkZBtwMRqIgM1O9G8If
RR52kqWlNeK8Kjz4ICnOXWrALQ80V8HDbQzo259BHJO3Byz68Whndhv1t7CTR6q5yHIfE3UDDQ26
udjRVkBZRh0DQjGPUMsfI3UK/EXYbn2+3qo5RrRvo/U1S9sPK22sLpVFm2rP0BQ91woBOawzyttl
+LTUKqzG9KQKA6VtBv9MIXDY+7uS7VBnjGAtffOQX38bWNYWGAr6rslpdCNRH7oKKLBWaKigXTTe
ifcbOgFiq9gERLID+bl4sA7ifrUQzZA9qURan7JuB+/NrckuljzW5fQghOoFXLgDgKUMBQbhk48c
IS9Qb9QJU0PyHd4hlOE6OGw5mRL2xsSYXgIe1ghbHZAR3zEjyifE4eAOuheqYzQTOBPn4vM54FAy
ZzqXmpATYwVlZTYDPS3IS/uxCdKgBsGmN99/weJPRdRec8UlZeZmPtM7Jo8N5oFy7GZgIrNIoFaT
jPmx9KD0VMLJ5VppqHxRr6Fe1hBfQdS1yvgbuRMLsyGaTPpnei/saKkqWXZQK7G8Lc0NKOAJqrdf
mCuWpc3Q0AReAmYpPHkhKXM2aJFv/KpdKX64ABD/7wNevpGoVw67oEL7+zsM9CB2iMTeUdhJFNy9
ODtgL0e7CEmY/S/OJ2b2RwfuoO1lBj8P9Xp+pIylEYFKYz9Nvh3DpkTxTZCaG/ewbP54Ta6rVt9N
m146ZOJJqeKealSDV2fAW3mib6HRYMQffgFAs5ImtJw1QXqdBXx5ZS9ieMgR6LbilR7ioTJHtd6w
GdlAxhGNwdZf399GMmnPTHUgpA4N61VLOUjwlnCKWvlBQ9CUSd90iGd3QHJ6ypRhRnpiP/1ps8JQ
yidzAPNHkIxsCszpIkcK91+GxolhmYKqOAoodAanVcwHFdNm5GPYwInN5UqghfJUvLNP1fnXA9Cw
c54mqR81LoZBsvBlx3ioC9tZV56rwMXyQAOuV9/bBgBFKxg/cWA9JmrCZjDoAXsRDtdhdHskOBwC
+jwOwxHrfGc1jlJW3xDN9TnzJpvTVdEWMu6JgVzeP7OYrC5HORIREhoUKmavyn6lzQIv/sS2Cxhj
Q4juaJhJjgyCDx4XUvZaIRn3Bd2znoFoC2Ja3pOnGRxYFCe1MyEMpNPf4ZrijgtHA4bdX9kWB1ir
9k+NkCNGEL3UUBLP9ZJ+9/YoWzS9yRXR9S2FODsvAVHnxHMn1yowpLOYnBl+zRMHdx81xOeN3ME+
5MbepBvjz9DF3X+B3XmTxJdB1n3d/wjamT2xJIVDoEKUP83/iHr3tuZZLnpYPYrjOLPkTbhHWi/M
QHrRrcxBbC1cSOUNWht8QtKuD+4TMIwJrr9OxlI9CSFLYZKnZvq0Tdn0aMHMIqKoSCyk4akrXQry
G8Qycb7+hTkuQzHcesO2MmB9mECxUu7JosUDS2YYpbWCdSIf3eIHYycal+rbRI3q5bBMYzyZVSe2
bRI82qq80QAp0ATFU/rse5Of2HV4wvCFIxGEjhDQV/sUASz2AGRh0h0B+5LTsdhGNXfImCRWRkde
ZYzqXyxJOHdaXxoIkLeh+vrG9RRdAqohG4STD72aUO0qQwxJNKhhOuIOddWfwSmBdH3Omdc/PAyW
M1WM+01mpbvj3wRkNVWotj1MvFhznLkZgG8Rb6JD2b6VIJq5NH+iWf2q8woVl/Ob9yV/NHK0CXBT
LjjalygqEZiyxCckRELxkEM32FFflpuY5wMVhgnTb4UOA8yNneX28rZvnKq2UMqisFIV//1M7LkY
XYbe4f6u2mk2tnW6jv1hq0Xm45lObBSOWW1DgYbjAZYKE6aAYRkpcHlMkI/7jxhnzJWhlkGmIvq3
85PtJ7pf6bGY6Sn5rDv13TUT58RsXZ8jOhm5FGKC4cOio9Cv4nyxfDCyVGK0njpRcbqtSk5W5Wcq
x0zvdhYTm97ML8Rm9CzFynLrfhpM6TPy0BUHzC+CBVWz47IPmgGFH+XnYC9io/7LQBLUnz8VO6d8
zq6TzAp0OecNyMS8h/B062qIqj/Li/F1Ou4Y+hDFQrJs3YTEb7sucy3MzwukfuY4CiNOzzrgjt81
9QeHVg+E6+fQVKhjJY5HqX3+tLMo5P3QEi7kahJRFg+lxWaLe7K5adtyuwQz0Is/XjGta4stoPr9
n8zFB3zI9MYUhmMbwKIPpRr1fDvbwflJeAcGmBS9yKZphzFPx859l9EmuRqQxLlhvSQhEBpG2mSU
64YCUvR3E+SmOFT6SVNIFWFePTO/vL2lgxqd/79Gmw3RcYJOK2ZYvgY5bmjIlHpaHwOkGjtobQvi
N6SY09xJFPvZaxA/DP6SwzIaw6/qYIKIpzmV+Abod2U33qDnINYckzNtpE8D+LCFAxR1LYKp6gH9
rcBnxEF6n1s+c0GR/MWEAi9mFHnQFkZqNQzs39VCbKIpahoRuH13vSYLIeEVekYyPuVM5sRTjNDP
AU+u4MghTNP38mLOe7tnCyznyNfZ4WbZEThGiqy/TOGcWnSwykhMIJtneOeD0i64SjgEluTYwtjv
QZPr+MhzRG/rcSQTfvSWOl1AhTfJ2U07RXs5V2lwqRmE/AId+qcQS/bcImL5S2+DF9lw546/E6u6
zcAJCAI+jfJ9neCK/PRFed9vL0Si7IBqZsH8XkwGcJWzN+tSyGdffXknwpgJLDQOfyK7nXZIiSJ+
ukJCM/xF/pUYojK/jDPubmQ3m+MF9MCnh82ABY5v1SWE9phxnQQr+Dj3WXZz23lEwoZk+/beMSXa
d00GwbF6Mak5FCdJPKalb1BXi4uCi/5ICjVzxw8oHzQMQCOn3NbCE97qRjQkPpNHXlrsXwM6vLXh
V3KUwHhSFT4Nz2VxVIfYaInA81IJgjP+yLHAzrBDftKLUD7N7fhPlS+fo+y4wZrrgwFtfKltQ/L4
eflfv+XlcZualAXhHAChF+S31hF+0uphc+GLkqs0k9MF+JJyqqAUluXgxjA/pMl7Yps4IBjwLG2u
z+n0YFmu/yDlUAhVLe1e/rhJum7zMZW9viLO1vh/qbDP6Z+HVwR+16nionIZgdZqDVNdqOh+P+Sx
QwwDiLJwe2F8kbRWdjaUKjTNdE8OD4rhgTbsJXnHkEeLaiDU0+sB59ykaBTWVQlXmXMU7XaK6p/H
P27BfCTN4z/ZVA+v62xEisNsdY3OrQp0Xg8ZxZMQqWdKcFljm98wxko/L2tqIh1YQVZiYTQH6ErN
RPV8fEMAYy1etXnGXG1VZiypOsJX4k+YHCNFXU700jGzNr5eJC48+1Px/OkGKzv/yYXNxo1Ge8oF
aeFROE1LXOzcSxqwzKQuMRYsEzT3aU88foXEfo9PpF9fpziOm/ugEDmS9kR8G++8XE9Num07XxiN
Aw53JnSbN5Gab8wnG1P23U00AmKKUsenwKvQ9CDuUO8Id+xXiuVbJxYsH3lS8dz10F/RvPcEuDS2
3lcIz5M7l7IPytx56l4y0QwEwzUYBa3Q3/ZylJPKE/gxTReaW1MMi1aQEccK/SU3+DJfMQ/jLM++
pPrJ1L4FRKzV4NF/wy9bPoicetvFxO4cDHmctPN9BywQieBq6wni3NwXEbRtA6w6h+k1jD02/Y3q
j6edbbI1c4gCcr/uKVFmr7EmTnbCyp6AoC0a5NPY7miLWtpmfA0JIiYMLuAX0SymZ1qMj203k4/I
B5fYs752DnNZ2Hs5/+i4Rp660pC9iPy8eks125kr/LMZe6V6I6FMGwqwFjHImnV9tS3SOtkR/76w
muOQZ8Kotp7iZ7Q1Ubr/SGCX1aNhUt5rkcBUjjTpVdG+Fgs/ujVXpS+BH+WTVa8fQz4a8J90msPY
8DKwACEj4XdMUhhosphyua15HYwlrk74GLXAgmQHjlk3eeTdr/OocSDonLI+3FywfHxkV6WvlpRL
UzSw7V064adf9SwivsD41tbLN0wA44AfranZcKc5jKfXL6QPQGAGNyGGphIJ49HhHQvkMrfWzJhw
jXEjWCnue0ZBtIhgdJhu9QX6Pg2fe4PUBA0S8MOeEkI851yeDUhPzD1AJP5+gH6asHYPeM36aokk
tVXynJWbiIRCmvFdSaJLNXNEiU0jxLQTjthr9SckyApDbI9YBvylQQ+RA6Dx37yFCM0WqeqbqvCZ
HEd/D1Dd5PCaOGM/KuVsAlP7DMqrQMu5J93EWNXZycbVvJKQt275Jcj/vZf2XVOCvSoYmtXJStlw
p6uJu+dNBh/ISu8d9ozILrRd9H65zdqMM9ex4INMIgSpsLjBP/JdHLQIsVpxIfn3w1YTxyaqjXCr
PYRRiIBgMZNeZ7f4Nha4TIuJpLjzvbTvyKa3YfKuRjACyiZ+SMQQNVlqT1ilEzqLgpgy9FgNmp7U
UCZBZsWpBGfYP3RQKlfb9e7qG8qqX4UMYTpz2DHdrbWp0TuikSwIAMBOGNRSNVEZb11+HspulRuk
PC2Ri2qjCrzZrhryLvlTOdMTCI3S18HVY5XwRgtQT68zQWja4kK0OOe8VfZL7llAp9/U+h5xn2wS
BbLFetwndk+Iebs9rqUVmOq1oYNyxCLXuuUyFw1CmR4Su+P30bDJcFBIH3ZBAu77CnCs9/VSWOcH
Xv2IClM7nNgls1ZGsF3EgPfkgbfansXYfymi+iXj3Zx42tdDkvm488EcBa+IJOwef5rhkgv8jI3V
hA+uiCQn9a7rMJRVPrFJiRoCMNnvLmVGxbLy1anejxXsz0EUYQ6OyZguzSzOXdsEnRNaGprbLJiI
4u+bkjmo76mYUzSXrhvdtPoT6ENMrMhJYAyHVGUwmeffQbMs91LLcrARijI4663Za3hb8JDxSrWg
6ml9Y2oletAwS7Sauzy7TBaVdF/qYKFPf3eVi5ly37hx3nNze/OMRg31Dxcs7j3xlL+XUH6Miw+w
eQOxP5cbhnAmZ/gKC+cHgWI8xoiHlhe+OcljrNxKw6G/kMn/IFze/AliM7xEfzKpi4mNarJDQHLG
eHbRLGOVBEtLiO3oPbyhyxv1Gz+dY/DiDnB0vK/POWWxs+WJLZIQP+/uYr3rmZzqxqAhshGMMmt4
qQ4Yp/RpzF89LwBdmQjdEXmWElht4E9MW66AX27990SCx33bANcGrQx7niLvelwZofNip7DYppGl
7148Yq1NSN8t8sNIBNHtwTOnDhioY77QU0+3/w1t5p+qCxhiAcPpfZvXTXRPoXzKKjyPpt4mV520
ojx4wswjP0kAnEKmy0JwN4hOoA4im5Q+XKYJ8AD0HngayeRwx1NEjUMv8EuyxO8aByhsav1qsrKs
RhLRg/QSLWhCUSZmFfwgvnFRqB92vlb/3v04+OxpaUrKJFRjowJwFtKCCK/7O6PS2O9O4xC6lGqR
ptFN7wqndETzTLrSYCl050ZkFgKl63F8ilyF6hvIukcNyqF2OMS+wXLVj+MfzhkTNVgFgt0nBPjo
n07RcRUzLrVVAYzEn4suVoQ7yJXcaGU4pRZoOO9mqnhvDdB8mHHME01u8a9FeMQCt1rIHZmb6BGr
V2vpUPMc0QYrwoohbQCsIs99kLypa714uxuE0pfHe0o+ZcycEdIIq9MfWcgEPKh15GKMg+btOcRd
A7Ji5LF8dfyNkhAVP3NmRL1J5z4cY0tyjQX/ipjvUWCld5Ytx7AT7r+maV1jqqrQKR3yduPn2cWx
LGmCXROxoys+tMyjq3T8qu6ORaMf8lXDwA4MjDNDa1c1N3ihc2NlSq98MuDRt59SnvPisifktfXQ
kjA+fHAai4tOMeVqHMSp22aJFOSvCRr6q5H+Iy4R304Mbqo8OERPxKhtNUUMOAiTp7uMqMt6Yl6F
+wGSvclDU2Av0hiFeE8LEEDYDY0Z99zWVDgQGmmsDYomGhGHDJY+iPgDrz6FXTb7kyvtjDJRyFVa
myl6kpDUsoCeuqiR86BXATqzh2V0qCaWZSeSwLo382p+MiksXyptX5ZdS1IhdpWb41dj9YuwoDe0
8hDqxF+AA4lvzN3v292EeCa1WlGbjR366fPaNtPy8uBY/APcwAP0PJdXpV7j7JJF+h86fgCDKehg
NpaAlpmwbnKtbPpnTc5nuqV8hVEzHa4/egWz/SIE/3a7Ee6tjUjJhvnoVmM2j78VLLM5+Tr0Ug+I
Cm8ann15/BJL8Z9yYIw7GjRNfk190J2LD9pYyAxQVsXa+dwEXHxEoOMBN9oocCYJ12NSsGBBob23
TRC875zmF5Euay8N3yespwff+AG/X03lM5BU6C7qoNhHj6ii16PkZgOhDRVfHPurYZmSzHcmzSPW
y6N4tAkWyV7EkVxA2XCdqEGd8t1OIVELpIRd8dIBKDqd5FzsrBJFx6TW/JRCH7n+CiXA3Gs/S76Q
5B1qk5uWKgl2tkc+9SbKy+90LkV+YpOXnDVZSJ9mjgJJC9/NAVGGZy423tMZ0RNEN6/mQ+l84ZTB
lQp0HiIcqfMubxzxeBZhtJIbITpswy6dbhyU00YecghwxzeGdrB7VTFj2wVItvIB96O4wSyTuk4Z
TlCbAjDH1roEeWijpVVBKnXyKrJQzIzzBVdNhfroNsyBzQiHlnR6voRhCPrCWFwePyqKanwMKb5h
A6hCspMLiuToIwYPuj2QqkeKL9dsvbBtjT8BFVOpHIZ2bkPAmPdpOD+5DSWiLKZU7MWfIB08vVZU
RTbXggLv5kBJ2e5gXsxI1amNX8AI/v7tP3lgduDZaMyGbRO984sWAWQoBK+iKtnv68t/iMNaYF2/
J65cCM5Z3qerc8YIfOZrcF6bUNnCfkFeFQWRODl682iE9Agt79GfeLFcSr1p032X3SJMgffvRmHe
Luuze1/YPqbfAjjeKvQ/r0o1L8MQeS1kxJKHa1qZgAimOLPF60KFVVtaH1719d9UYlWaQ1HHLhFd
6GZhx5hdEujzYxOhehO4GTRPbpjEY/Mg2oWcjO65Hkz2ae4UlQUElfhhZLp/xWF/9mVUx58Muzfb
KTlLyUtg9gDnR1aEuTO0njn9oEsC3Rbyd6Km465BkmUiAdDPBeuIShKI6liItJvxtAmCOy8HwLEC
mTQb/O7wRi+KDcxgyovJP9fJOT9PHpgcESjoGBlpsS/Dg1kSai4FPF9oW53qNzDPq9iLun1Vgty+
5IqrpxzP2+0dZdH2rIFYN2+OhDtWLqlyXhX1gpGTdlfp1G2fBf5T1Fry8bY1MenZgAYPRzkWXseC
2Rh6tR7O8W/SRm+UoY07SEreQ3LLn1jOxc+PsyBTUHv5Mr18BBaTTxxKnX+YbK9O6uFloXneKC7u
1nMVc5kwPpcs3IbCPchErNKyZWkTh9frsbmhRsdspgavJ3+sLEEvZB/Pncwz2c2Xi9L1z7rBzVTS
skZZfUZ4GWd3+Snuxxq6x+QJHEvOpd2LK1uZBuVSQG8Y/y6DpyHYw7GZI8ALGLhvO3NV7y2tpxWo
PkPIWf5aLAozaknsZBxk1MAJp6uiGaKInYstQzKEiBt36d3dBPaVk15y3uWITDlnOpCj8K3zLIMF
L0HPrWcSgqCIcE7dysqMPT/UIffEwI/e1geWszBkdJ7m8FI5VdNwjVN+9NsKNRsSbPFz7BmFtkT3
o/1pgtXA5BtO+TaXMDJ/z8P1dGZchDVS1Tecvak8hMb40QR0vnt8d/nHk3mvoCWVw6cK+bgG3Nkr
bivFTHpVc+KIiLj+L8f93dfcQ56T7SMJFNgYtt/9lI1wwHrBqYTNCyUI6J5AzYxdLkp7uyl0vXdt
bNfmOPrMFuJKilRdawwoHJOmCWIYqjxkAbWLSemKlifTwUsAgFzSKdP821kr2XKAO8X9Hlx8vlJK
D+GVYTDhNRw1RWH3HUqLOo3pwCgqnR/f37zht5BDv8YrGUgTnozoglXIXbG68rB17N7DZzs8OJEz
tACYr14G86/McIJhb7Lrn7eblttgo6AJbUSga+kp0ikZGWsh4XHFsnvn25P36lV5lxIkpNcqiDXD
iM1nlZ2BQ7/ruPkU5SfZgnhkhJbwZ8txts2FTY1WUS+oJxjNQi9CFyNKx0LL8xGF1PPA/JA0W35q
GIUS8v8Z2Z3wGEY/Sk9YzJ6inZoVMBm87VHUgX0t6oeqbR3ebzR4Fgll7m58pGM0nb4P9j8QTBoo
RBd7LWuLm4wOLGM20lz/32FAF9v7FJZ7DioU/VbbwTCLTLdwt52mgik3Z6b1kheQapGYHYgp2SsI
8u7zRbTn6wfUJaszbqMHYDj60glq6VOLCHNmV2+jOWdmb9Decsm9Ia5SVa2BaabyASxSndt8W5Em
+P0opx6ONAS4WE0W8U2KiUDMycE1aLBzdQulJYEsYETOddEFC+WkqdL4aeemnHWxYTGVVniq1aIC
RXnk8IJZl4NluHEnTPEmHuEes852d7S7IqRT8ADTgCTP5m0g6d/gY6tGZ0LesPfRDdXwxPhNOt29
4okdWeoh+nzfuk8G/Z7vKSzMFAaag8HI3mFKfHanUYtRNOr+lJXPnm8f7f+vHG+TNHKBy8jzBfHO
8XbwdJYaW96dJv9QgrUmMwUYDCWMCQ++RJJlig64zjPDLFnamRG3/JRGpA3NhwYBw710ZXh+jdeJ
fkKzFLtFTCLG7D2/kw77iT2DLKbuLFqfcUMpVAK+LzkDaYLJ2ifzCSuQjjFZ4veUVWePLflerNrx
azo8cSDJUNeWmyivacZip2Mw0SPUt9GcqgRCDSg3WIz+IeDCbNPh8hBSR2Z+aQdEzH7kkM0jxQjK
XlIrb/n/MSJyOmKKV2NlbAzjWoqW35biGF4sx4b3wwMuQyvgRAaA9knfaYYhWk7Fe6JgR4HtVZmb
vDSxm3d/pV5uH9Q4a3rpRZwdnQx+9VwL4Ym9WbRTrplTJAJSwwfoOzv4yB+ILYqV/4tUNqVr761J
YoVwVQOwOn1htofB8MW+mDDrHxXJ2Rwq8IfRg+f5tUGWGuHL5A1/HQnlKgntheThv3KFHC4bVz00
yNsOlF+VY2SAu0VKSuF0Acy9AyBA30bevnA6RgMgsm9ZRJH0fvtcd0BS7ksEBa4aJy8GStO5sVNR
jBtyhuDiiZ3bceTKo4tfS+7vq+tguteuzMlw25qt8Ie0Hx+cfYx2shdfuYY1zKrehSRNXNnGw1uT
lCTL0tH8R9e4K/SotHHuRVcN4OrGnKwANAjMm4E5pemiC0uTZRcQuC0vYWX5o/TiXp0VIt5v40ag
gUBiSyKyDICsw33QOsGl4olCvR+9eKPXIeNyj+KjSdacJniZtbFwBoLrZ6iZ8mzkXztPHEUVWQip
36hiTZ8a9petVvvPMc9KNGLgmYCvFLDVoz2GTnPkBCZg7VZyRJXfKQdmvhPfAk9FZr2OiaLORFko
Ozvj9px8dKPLRkhTfK7yOOhYs/59/63wQ+i+tt+yR5aw7c4Ck21PN83DO0QbQquzvfYaumRpjN/g
fKCVceA6CYb+tbN7PGz+m+/HtfzVv8DCRcRl8U6UG1gNgtg9svmdpYKl/vYD0TxUytUmdhwX8UJO
kc9fapVeMIG2McrZla2M1c3EWmrztuF3zCHTn3o09AvTHC3L2VWTI03xc5jTMzpANnZBcoadPe0k
xla2z+ihcyX7CTrBtaP+EdC+geZUaBx/5IOAN1e6qjdf/DuUGpB/TE33eLauB235hBSXYefchVSI
cTFpiMumtMZF4amHnVnEbFg14Iq9Crk4r2ZvDP6IeRIxr8Sftl976KU7f4lTiHEvBJLoAhEmAlik
u36E3tNyWr3QQg8NSqBTjRG8xQuGVvm+9q/JQ/balpkEMSqX5+yFlGdhEm6agbB7UTr1hYbfP8aa
UUd1XxNnSJiaMfPvnSPV7TKPtll+Vz8UZZYNMm2Nm1c/sDFJ+w3swVFW831h4Yyq1nsPXfYYRLWC
Ld0ndNfk+hYfnsdq0GQ4VB1bO0UVSNAyGACoNBQnxmIF0FgZASSzGiW6rF58kGBJk2DyPVM9gSnH
nI1QkoJDqCiaHsQqMSjZ/DSgKhdc7NnnaYraswSSLGLnAhWQ1frOzeJOLlocb4RxjEq2MF9fwKsr
1SOEzxuy/42G9ZAJ50im2WkR+zbST2aflZMGc9m4anCRLO0OztVxXBjBxY6jth8VLqMK9b7NLQS7
qSNufmYZMm4bvYlBV09c2jbbeRfUUey2qJWc+iEYCV2aoaeS+hWhBRpwQsJmHUq2ahNs2jh8oMtg
vpsC4EeCSjAMa33dPAb3QVjci7s7or5Y1W93j/UtYWe1MlYhEBs9D98wKovNp9zvW6opMcBRNWj2
UfldpNC6LVJ7BhMJQtFnkdd235xlC9QaokCHafrPY7w8oS6saUg1FpOeAN46k89Cocm5VeAm9D3j
3emuOmQk86QMcYqGTq0W/+08A2anMhXE8FI8++BV7t2NrX2sqi+UA3IhtzbLlrOGWaqtxZKTQusL
G0Xfug0ybmTbf1LjAb7WCY6GnCexAm/wfIm0s7Hf3wCHIeKfWt7xijcLoWKJo4hsKXBl4ptv2P4C
SWlOTFaLNbmgZIKesnIdCYoZSohGb46LNfqseHLpuykJYk6T6nsfqafzAd3kbQ9uMWi1iPJ9gQYu
ZxECu2eScRyRWbqDG4s9cUg+5tiSRwJhctXn9dFPe2VvQU0eHEUiEtWbW/355JK+BOVCvfS5h1tP
oEzU+bd38RaW92KFjY+S6/tnV9stXOwdEIfymagTPd0dBX3CFyAk9DrY6+VDOYb8T4j5CJoW/TmA
r/N9PcslMaOVGJVKy3iWjmbuSFmBqSDM6DFFVFsL8XgmCnjVrT8xMQL+b7ieUeVeQKmGc5ZSKL9P
KxBFIkB28G3zP1blEhhWgqpgUNu36xjJbjVeN/yqsGq8uv07CzSqEVfPfZUUPXeh3fobMX6q5MXg
MliAeaxl8MJ2L4eXtmv5pVjLFswEwObqr5s5KeFwOxhmEgpnlQBGGzSn6Jt7wknsLB8jXwWkPH/A
egxuNXh85U9MhtiZYF7H+EdDTAYgFXjHw/tgnRM4kf0HvmSTIJkyr6zaAW1ZbCi2FgA99ukgsGa3
LrtTrFRj652126yQO8KFXlH4cS3q+w05wJSr9Qel5prn53XQQoxJMGpSnyyD4HdrNoCwFDF0fG55
ElKNTZQ6Oo21+luuFe0DX+PltkcUivFimFf3hsb0j75tt7e7FM0U7Pau43nq5kdWrjwGOIJCId62
55hTor4s7YAzMkE913iNNDELly29DBZStRbCs0bAlxvetNW2Mc3nIaqAQRKtHNlKClA3sgm2fa3G
l+2qe1cbSzWGGsOV5n96+p4uKOYyJw3VoVbRqLbRzuOP70/i/G+bX6wCHWhbmEkh6ynABpWAR+vh
3vueJW9s0eUhhGf1E6hOGcMx6F/GCQ+jsTKO16/Kf9HHAw8cuP7Otbg9yCB3Hz50GnrU5Ix4PCd4
rBxnHippOTOrTRTYRZlTtkSNj8BVh7xHQQNgT+HGMfJ/3SRvkYU8naj3U46WBk8kz8G6D8T7mU6a
I6plJkJode5OuubHKQVQK7FuZIfj0DlupnEssaKm8Rwp1HHxDbgeIsBKU1mONdiko1QTD8j1lpFk
yVmVDfdx6tAaTmJVZ0CddreR6lQK1E8H7cfSSdXns3etYoq4IO4oSMrE458cSq7BX+U9ac6AOpkg
sZhwkSgPqYgN0kGxPmQfO4/cIOlAHUopPd40LCrbkr+UXaWN4ex1RHvfpsFOpXcWyR+a3xe5ESDu
+PCHjPEqSEQ3vQ+qUVHR/vc4+T4jyyr5EHv9CRMXtXDGI4++CvGL7PbF7YpW8mqb5H7T6rf2sgUT
gf2DNRsVb1LRLhaSPaUJYYzXgEMiKI0OFAedvFuapxFQl5hPPm+nbcZdesmskb/KMH1kppWg9R8J
Tqn2HSdeiN5UHwmv9DqJXJTHUZfa74IpKFJM5+FFUn0DMPtamD0VNjB5PmAM565vLIxqYwmU35ko
yXutDYdynBa/Eeyecchmi70pTbaej01+LUVXFO9/L6/7A057hKVGGqqCaiPWoVFlELfcaJ0pOUtk
FkcRqC+k98Twl7rFBbDuRd5k1IZlnp7I3u0ko7o6kRjxgTp2yZeF0jN77ctsujGam6gRTHsDvGY+
oA3W6mpQq8RJE2+3zDyqr8g0k+08JN00Vn20KU7eYN3WLv89i5tY8dx15ug7lXqfUct8tYBCxiDh
sjVYNQKG//7HDTocd50kS4LmSB98sYNHrlAm4wlqj2U2Yxmisr8t0fYKUuVcyHxIjKBa05JtwlbZ
UtwshBf8sP418VjpahCRXXLPVoJNPKPayrVKN4i31XyrBM66Qn1zAkhiirdPKPb1DhRGzRk6zvNY
wnsKVxckpSQsCucm9qNN2gLad3Xm7PoFmxQK41D0NxDIt6TbZxgQHSF+6GqUv+0XBMQHS4Uj6UqL
hjWErnLmHokV6ajDctAOSj9g80p0dQVyYoijSUczwFaVmjWTYKQ27qY2GtgdwKJAIcuPbQMROXsA
Yi5Db9iqnAN3x4nmyMOj2yVj4KmShYlU8p+22fQujaipev9vwRyZsSugcgRFPZ/MBUbNUAZ2dZju
7BGKT5oUNZh5GDT4n5ToI0visEYDuG+/aIb0rkES4zbZNL+MZgGlmWzQE7oOtrJuETgfheNqNv00
g+sZOJBsXxRg0+7trCXqJhPhlb3i3D027aGYAgNjN2Ka76np7Jf5tpQvdPtn/nJ+iH10npOsl8fS
x2mygwVz7yTkGjDq7dLqP+I889EHJHOjB+VSlazNiy7aceKTm9l1NRPIYsTjvfpXETJlhLEBWvlM
JvwTfIbVqVN0ZbIljHlPLOQoUoO3QCpYbzfgvABtRYuQudTStua6yVZJBtJtWKIPDhe7H2tWwIxk
ByIHv2S82xP2FnXUbJwHswJpToEiq6CzW9lrCa/keahDgA214AtnG6B5Mj4HTrg59MbV1Q9ciVJI
65dZ/DxVlAI23qXb8Odq164pbXnD+O4BA0582ap/M3fxuVs/T9IvUJ4rt2Ko2i2l8DODud17Z9Wk
IbSkDzPfZAJdTnlYCQotKBnX8eokXaCDfBFR6E4XmBznivfC7bPBSqQwQv3esjlAIJAMo9Iks/A8
HFS/LGHA4OmhHQLkN/wWe+iOmzTfU1doGV9b1bw0RwHO88oqA1LnTaJA2sCf3nkQp945WkoWA2nq
l9Z+XUqlqA5J1u2WJiuCqYmFIo53h8v6S7KnH+zteZgDSLXjJ58tIRDG0GOJJo86xI+F5HYaw734
gxlbnYZzl5rVo31ZyLhYe6l9U6767CyA7LJCKRs9MFQ7aRl8kraBQHZzgx3ygBUJuQFOAR53ZQkF
ZtBlUJYmXWAUIBFgZ37xn9ceVd0U3My8lD9vhQOcxWYBUO/UD+MTsxl+vPMZqVOQhHfhpQCTZQtU
yXGT9AVLoBqxLf7ySdVhgcNNilsINurDEVjqCgCh56/PbAu7jp9wrsZ0MAGFpJqanb6RnU+54GeI
gjMH7NO4w6MiLdBnQn68XVkurD/boii7kb6p6IEp2hh4EBwCohvzQ19NJejwjsp2Up7LQfSKG6sO
GJpMdQu1DY/+zbaH3AKCMQzMZ3H/ZfGFZz0lqYxmfXzDQUR2f8yUBKgQxt84zRZ7Jtom4eYPv54o
pnaBGChb8F+dAz5JbX2j4a2YQcq3tJu68HyMt53Zc3BIWTBCfYZ1l7aafxVqhiAqvI8AJh4vW9T1
oJcU7bko+95L7405yhiartSFart2jHs88ssS/JDeRoj6gnK7Iuhqwl+MpMqhWbsWH0rcDcI7CAEE
qAayzhEf0Ns+P3MGnAekRIv7hwK9/voC3gNnPJHyh4BaznXb1qd+94/HRkUdj06Tyg0DRnhptaz3
lxD+mhIl0Q3fM2WBE9fMBXRcHZdONuv/kamo6IH5/lJjWHdB6nUk1ZiV38M0szEmDz6TwWSWmeMU
0GXpqItPdn1u3Ir25xCPIaDpTeyxIKi3j7uIrhv+HSQ0FPv0oPQVpReOFYLe9mY5zertplAJqeGE
jdNbDrxir/pfzFQb9YqT6pblhD9OhpWmR7bv0YK88yYKStDZwS3UiYUgaUmEd54oP31gKO/PGhzE
sObi6/GCzMRxh2Mf7TSfaZMlMbobECuuSukUUBJIDkMtQNpYndjdvd1pGT940CR6ukXZas9x31rw
d5yQBsPSiHq04ORHTv/3dfY/jdccU9R1a9zYjyzviNjfLBycTmioCrPvZX3V4r6wCkAsSLdGLsj6
o7npiRn73MIRfmaAh2t0NyEvksh/VsXzBLdcZluz0UBmBLUgsPMuT1swyuTbkxdtqgfO6fODXv50
t/MSfrc9TAcy/WpaGDzkvwyUKGZ1MxEwctgj9pTF3aGfaxVBTAISgFBvFFpCcYJTWTwl9dHzb/M3
UM+ZaLcNzDJwXti+RLyKJL/42bFlLMZAXP/lb+56uy2+TwNatcOhkw3PHW2izYWeV9R0al8X6zBg
3lUY9zh8LYb6JizV1lATdXEfxLMsI8klH7oRqKxu9jEWs/gUUnt5hcP1RoHfQ35CRIOfmYrvqZm2
wYpW8pt41Opi5MK/n9OxUzX7mXUJlVHSovaWERFo30l1ba8oxclN4pXGoAAXeppbTLnwDRqf481I
gYI6BpH7vXA9A4Bqa4wlrzyK4fiMcAdis5abfF74oiGDqFg0bjTu67g6kia0q03twtkQzfxW7SAQ
sFXpA89dgth/lUNtvuHlTu3XQRFshPwlF6cnwmaoTDOGS9id+VMpgmWp3EpiO4vWkfnJg9gZuGfD
Anq/0wQ//BIXHSeWpXKj3lbSP/a8f4plodty86zmCnDsK8MP0Asn1K7v/STHLO8Ldms5a1ggo68N
El3HiHSLIEh2jSx59ELJGuupvkrnDbJD5GpB6K4jBQVxMMM3OmJUHZ59kzRlLrv6CPZ0MwDvvICC
wtm/05S97Mk698aUzGNGMsL0Z+WltmsSBIvAfK4SWn4kHDaWy7XyjcqjzqjZfozPoKKh5ug6+hpM
965Vl18H+RuN5T0IgrSEExUPNjgYwRhhitZXfWkpm70oVXHQ4RK6KR8ijzG6MX8maf3/4UeYl9sZ
VdEq/gvDw+zV+ji8SNRr1NVdSBHVNQp1YPfL8oa5RM11eJHF+/Em2dLF5jaUf96Sn7ZnuQQ2lwtF
8N56rHbuJTlYqEsnl0WZIxV5AwZTfwjQzFAQMnLfH+Uvz3lrq/9y6D2uSs9HckPDcQR1OnJB0u7w
uK4mv68WNoaO0Cynf7zqMZgYnWn28KoSKm+JwC5IODdEO/O9l+yQHqmi/RZOQg9ad7vecMfVHErM
LOTRVgWkjyN+xEg+HunhchoCoH2b63sF4X79vTRYSAdgYw5MUEVYktubvUhDqGcki8U+/ZZ3FFi/
e7Mp9rVN+q3zJ8BNiPMcuWq6KXvK4BLyzRlTH3aTFveM23thsb5ZhOnKrIkbJ9Vh8gLZ+1CsdF91
p/PIcc3oNR6nlQEUr6Li0ajXqHB0uoEb4fgyh9ZMiReu1zuEqfF/stnedJhYfROKn5TJLHBx3mH/
3vL8/mqYU6yTQR41zpV8+eGwfM9/fKdX42egAf2z8yObygjOr3wFttIm+WyAKdujfJE/b0dvUoqx
TAxlHj7zciBNwugceK5Wx1NQtii1KBJE9Vb3Ps2CmnHZTJ3bvS+hNUIp0k2luS6u8lfEn8BtDKuW
FD5eunFPYx02D520eZAJ6NDaapIZum6K8XBjzGgSaLhHD47sibm5Ysdx1c7okcGGvLAyznYYSGDm
A64GaZdacLLYZbfu/NflL4pBIqfM6KkIUunoA96iWJ43V8RL1E8Wxy/J4Xmmpm6ZsxlHSuMNesyv
o55OvstXNqpAJ08tjtOtwRex/5y5NhPGW4vLIRc2ji0LykSAeY8kfR4+MQ7Fsi/7Udo3KB5TqM+8
lnfh0nsTyGqydi3tKqjVjfRgS3pZLv2mXbjjbXli9SvoKlk+sMCGZZMx3Co78Vdqit5BCdg8idna
MTwSHmunpW4qc6zA0gMRM/8JE9IqYHp4ebkdaFxBCW4jAiBBOHzH0d8fTILcH3QmxloMIp5L6l5S
cbOPv1QXw+rNfdNGnPSMdzkPoC8b2T8kUi9m6ZZfITn+leFS24WJwd8s7JSN6mPDJm7f3Al3Ax/b
d5RxCNb9qcour5CKP6T6RL8OXzqv27H0w98moVkrEo46lcfDSFWmqNdnK49ssTazIKnQDPplIk+g
FJ23vfBNOfsvNy8pnKmVQ/4AXof1sgA6cPKd4kmW6HJPROKjFts1RNURPhnyoKL5DHz0KDVu0ZLy
MoPoFJOCADlWQgk5gWp6qXl3rDPHKFDLXj00BSu7tPO2g+xHWuCSU1xxPTjkPDhkUwREe64K3oLU
u870KSYjCQuxIwWWb2o6Xuw52GRybyTq0CIWSwVgXEY/eJfsC5gvxJ4S12sLrC8WEJVi7sL/NKMS
VWILEDCvhOFuX/0WMqrMZt04TPDK5+kTdDXHFOQQS+si3XmQRYVqf7gk+s39u6xxzHJgcRiLOQgE
GqX/UL5bU1r14JJ7anT9dGKyRUUSYSH0/mzt+ZYm1g1tOdpEY6VY45ACuAuOVI9nDUj49URiST2F
ByYbFYQwgy268g5NHv95tyDnIl7DeFIN0GpiNjdN5BpeF/XFFPT+sRHlceIyaqO/cEIf5GcNIOBk
chmuzm8fh7xmJKRxY4gTa9vMHY0df8AzuR2+yVcD2DewHWzegzXzm77eQ/r1QHTIsT5YTIFaWHzD
3erRZA/xaMNkG7DAWl48MOcNKZ+jhLf5aXmvmh4oy6dsPKx4VwdqZCiHPbH0RdaeESgz2GGeoYB1
cyF5LMyVPXOP26fbVGFyPjymTSmJFHFBR/L5mp1ttFzO/vF3mV2MKNnByQM6C/Rolu2S1jRfNKvi
TBywX/T54n8qwnlw8CHfcM+1+IigsBvNQVDxzkPPdK+XrE5fSYKTNZR5dws9DVs1/GAw4Hv4lt5E
SH2eP2RjaVvhOMTtCIV3s8Idf+B1Wcjk09BO8KPcupZBIvNYjG8rZXpyPJITutOQLHf+IvApbtgZ
QQcxw4523DsN/fdJS8AsTkVZO/7ANjtgkkN+JFakRxlzNvHFHVausKhouE0AECni03lxC5ViGugM
9Vo335QbPGBMEUPNI7HEA5FJ7Ai9VlmOgCcQqGG/r0wcDv9krP26L1DPDnXLMg+ZhlAUAHD/saDN
sUap1jZcw1EhiRQVYT2UfhVmxvCzjfnoNFTpLsyQbnIi8J8clrW/S3YgdwHFJdQbtoRgJqS1g5dt
n5HQZGkbIlau0dVLbcoWBMNqZl7EKOlqUXLqqzfSX8+IRYtgtINihB2CEOzRBPYT+fC659MWxC2w
mBESFK13a/MjyJ2RqToLluYwGW7XaTAx/HDO+HC1xVgZd5Dp3+6SMLuWT4x4iHJ0tY6e3n5qEtee
OVy3kqhN47tdw+x0YfxlTJKxTAlxHAXqv7O6aq+aMk/m7yQkxjK5v8cHOLJ7VF9u6HVB2CnLciGm
rzw8s2HEFwDa9SjcabFcBny8imCiZqHw6O42tKq3Y70NWleV8llFWFz1h+3LpuqpUVJvv+8OV11W
ky3t9W5BY0PWXsBnCc6auOr01dMlNYOtSRSJARMoJaNRmpDch3kvxGWtKMbhDNwJ0IbaqT5froAr
ZlxZWDcatp0XHiPsU91mQHZ9qYDC32SY3eBHA0B0ELwHPqay9yDtf5UXavrr64cBqzMj/NYF+84v
hlhatVI6OXuA5vqWCa2qkz1X7/1QBKdOmjsqtleZqwYZgv4AiPKDZLNijTJUqEVeecX3obAHa+W7
YuOZ2NVPwoRssyrxIJQSOLWYogW7LFED8zhwsvdoS6pNUQJwn0x+TfAz9Fadv7EymjOkZ4iCHiIo
YtyJxSVlQ856zFrUOl78KPqlM+jab5vftvJiU+13vTOe8zzue8aQX/nTPjoJl/u7e38HGTXhGALe
ZXD5fbOLXtqPdWB1EOeww2k1xCV44rfJFOZbvV8NwYPeS7ssq2clA2Sh0/b9i+/D3dRqbtCQKk9e
bu1ZEzw9RwaOFupyx54XsDuSjy52kI0f17qnntZNEc3oYFsSzWyOijtAnj7HyPIlH9OE0qBagu1Y
IlL9ojOJldtpvO1OTxDr60TCl1uSajpM/IpUCjzq0zM6O2zPR5/IEhlWIc+QtsRVuMe5ZxK5IynJ
hkZ3wN3w8jdDdmuyKXfcf0Y/pgwMsWmteuDd2rt6HZpOdAdu8qGRniWYcRs7PpFmT+b7FOXlO9MD
/e4xBHXBeawZlpfpItOQCrwOV+IxODFmz6jNmNz/av4iHodqqPn4zol6DjB/ev4yfy6v57LjIYtQ
yg3URSGmLBrt9fi1BvpvfvIaE1kePOF8Bcv0UkY5EZ+ZF27EykNKYtTP69/AS2sWSTLC0xT+tv/c
yzpvBrl7n8Tm4g6XKNrv1OsF5BBWlXljNvpnf6HDq3dKvB1FHpuB6zWjf84TzZ2BfYQuHRHDh/5z
fN0koWzpl4IltMTIrir+v970HQyvUgUn5VEmbhe/t9l2BpYcIdNlK2NfiD4md/R7oM8xaPJiqgaD
x7BF7gEv4nUb7RTSe8lyzUGXIgE4deP+R8kpwRSEV21jqhpWKRguVpWm/x4GgrPQKj/eU1PEmEe2
EkRbKT1bUM/QxuKabVZVZEZmgf4u1DHCO2cw0FMZtefqAtj8VOCYZbkdTtOmfrQXRXukUOsUlOWW
EZ+7TfmkCa5Z/SLrrzoMvJGcAKkZnB5DcTkfKsu7oWe8KKDYCpw1ONfbPsQLpVhW92fTI8aHZRK0
dgr6ao9CFaEfGIoCFVWZ5ZMZZEP3TTB8UKylxUv2WET7xzCAC/rOnAI0TXhSW5tLMmBgyTtfnSOv
MgWsqdnhjSFr6saI18sKkLebIm09alPiPjEQ++rXZ2yIh+l4wJz/UZ7Qonug0qe8PMHdtW2VcmXE
9lQDMMp/V5BzsL7bwF0MK9CzonqLw9cSba3P3hmWH5wzc6+ypJdjw76gm5MOyRlBSOiFrDr2ZECv
4PvvZTeW8ETFb8cCTGXWg+48ua08oaYARyvx1szJ5gXq67F8w1T1RZ+BrruDSdscfBLTPBGiglIr
KoAIecC89W4HxBpQY0Z5BL9knrK9FRM3FZGtPBJqfQkrUcaScLTDOs1o45sbyY83ZvrWuBODT77W
MZzRMXJyCcZSJBLE8oV8SuY95vfPApdRxDSwh2VkcC3g0okESmQX1LUvN/dTIfFj24t+nOkJIRP1
YGh95ecjOpLoKGnB2fUlt6Mf/POP5zmyJb/Wx20sWD8qokhmmv2aBW3GvJE87Z14wrDfeab4jQWM
9lVkL/LjBvtTMjDLKBgQr+5d2nwiuuTud55suwp8hJW3ujsJytA58or9nNZnKO6gSY5vVEfji2ST
/yOJGvtYlhQ7RwOyfCS4dUZOpth7kiHVcNtcILEvmz1kX4CKDuJvOIBTEbD+ULXjyUc6Xg4UUZ7m
PIXFqPcyl92vL+PHNXURAw52zlzGdfp0eAP9DXTvBg1JMKWDnSXynI9O7vgSQec+ibdd7ezDeFlg
ccOfmBFNiOxefX0Gu0LWHqlNtfjg3L2U8Z7RnRHODYdi+bUt3au63l7su58TXwCkRPAw0DwxEot8
pMT84aoYqwJztm5xDsSdl4AYPLMQ60THO2YnXxy2C/CH31aaMAOvVxD22kaCtysm9uIZJtqKZT2/
bVp0ncJ5rpxUeUlQWXSUFRZ3WRAS6MKHXPOypj1RlDcrSfs506k0/h62CP5oWsjLA7qX68ULCxo9
+YsgkZ2oDeYvWJYhKMlCpygx7eTR0bV3jbL+BhZdCEVkXE0Cd0UJ1zl3+5lGIb0cm5uXky+1nITk
XC89E2ZHPS8aRkGyNgSgE36/3G0jqjPHA93+y+6O1sEPk8fpBLmnq8M0NuaJePW/Yav8+r9KmwXt
/7/FMEaDY5e3o4tKLj1yzpmIimHiP+jIgRJoW8qPaJdqK73KVcJOuoJteyzthsv9zjZAa6yU3HZ+
pZ812uku4Jh3kKJbN32Y+XKy/cKL1fO9uSfrpgEAK+mruWxRlIOBA3aQDk8DaCBN+lWFp33PFrx4
MjFkWlQbktxaH3/L9BuMfmw0WhmU++TyFaEiPi4et9PX69kz+3nKPU3KbNdc1GBaXh8wYvdNcaot
F7a2lFORjN2a3N7amddoZNdNsO3pWwqJCPHsz7oAz4urcmsc+u5XLQiy6qrOMjCe5a09mbFiWx6k
rLEJdGorBGGwkjtWbS247EQ6adMQfjHiwsYtCXphGHZyLvf+tp4U1Y02gxnUKvYOavm35kYl8s4x
qMB1a0I8g0a3HA+Wk5DguKGJKIWR5Y7RXQQU4QkYKs+n3wy0so2bGXGUQadyOFQn3slvWMQpJDHc
lYVrYlUhvd9kmtnqqsBDB73vLVXcWOr8dr3tabTEQia1OspM9+/NLg13EqAP4PSJlnRtIrimHKVa
VbfgB/PP/DkUnBKbdlo8Y/cMM4D/vrLSrII43o7lFlzOzfpb4K3mi90UL4qfm+kkYKsC3lxmGbTr
xAwsIqODrtfV6MuYi7ywDYH1qiREM82dj/9Jg1PB3PjX/LP43E7MXmUp/iLOep2qb7xg6GwoEHVc
ji3qZrtl2OB8H6NYJMPfP+5kZyYg/mQKfxsG9dw5ZP9NDL6i7yO4eTu4Hc9JK36Ky5EqwUbWQsa6
Vcf2mAkmXx6+Ilxxm5CeFqEPEwKdxMGBqJCi39VSjpDOGSA1R8yDsmDOdH2ZisRKIQ7plY4Zv+aN
0JuYNS9Tz0oseWIhxgu7LtqcWIELDrmk5pNBJ6IlM/m63So/fdEo9VjIvQDy0kxyXo71WCpNkl7m
8+VKvZ9EjF849BdhiWVSzNArgXBSbUIOs57aUVLAkn0a5FANW7q/kLtml/q1U26/tuvlGYKEGrFL
GIiH8SEQlsR96arC3ysOeUHIO1lC8d8CmBKESSnjERB57jGN3JwwP6BjSxZa+YLs4EP0E7Wqs4aF
NdTtqDZV68yebdF8rQud4lUOoIWfi+ZfSCoSGc0BTPCjilUUZWIXBJ40Y/r6t1Q+6fqxpvIYqw0C
po3D2wddJ9hbk8UGeZ0zPyf/BcI0eOFTatT45JHg5YFkk1avHos/4fwaYjRi6pb/guje3NHJdQ5K
5TuQ7S7s0nPDPJ8OF//0onCvgIfFg9IGEka3ykICGBBf2kGgoM1DFPAlm14c1GuD5vqnt5jttUcw
TWJRtz+w4GlMIJN/qBH6bfl3lxOIqLDEfde6SkLNelwIo68LLeIt4XZGM5JCYII75oipUOyJLmL4
rP+3TCDyerUXuT4vrBgh3ewG5Bf2p7wlxZPMH6kQUMfpdsOUJpos4LDSJ4McGJmDFP5epl+uo/Xt
7i/WRbzGEgdrLS25smD/KMm7l+NSELvxvQENtUB/is0zFh2V++eXYpZVK5SvgaZHyDoFqrsf1KYX
eADCZ3JIN89yuvrCd7unq4IKAMi0TSSxFr4EJ6UurjtIi1NvqTJAJoDYvFo0l5tRwJtWremPEsf/
BTvEUhpqZaEaHmQOUIXbqBr4S2tvpltmfAhapZa+PsauovXT3vQWdn2FPuIORiSoBsxZdRX3dhA8
3Pm5YgLDVcYs/gneVKZY0wFFnpZe5sO8pAjCgHzZFcyFVaoYfObRyVa1jzonBNEuOKi+Dc4uphwl
5q44LKmoLh5UEPdbjOuQxWrXY7fXhOw6nkpUmp7wP+RNKfk6i9kW6LHGAcfWFdINnMQ0CFzg5050
e5085Jbz/CyXRQN9wL0mgSvX6p9KhbkI2myjF47oNbgMXqVXjYzNQqWKN3xIvmibH/v76VuaC9pP
fJJccNxYoXDO7w7NizhnBxQnIgTl4l6c4FnmYc+uJFCiLlieowt58LoRFeEzd9TN07yU3ibnw2Vl
RmghOy0PUcHOlyUopkmock/pcHMCawYB75vbkQaWKzMy8KjrPkFcVC0VTws7h7JWD7RBpDvAWk9B
WNHyO2YpynOOh6QifH0l8ibT7d7ZVyHwjptjWGmTMbnR6srgLSksQ35cSaWTr+1zbzfPXZilrihF
T4EglfXo45RF2XFFqK6auvPlnmFt9N4vFUY5DcGA5o+8owpGYvzU8AmIrCg4wStgeMIH1uNz+J/D
+kUPXJ3XDWPE/RwTjbtPfAxFIZWJ3rWS3nzsx/DA1PqFcdEUda8pQJpQFN2LUJdH5Tmyg14cSKLl
pbrNKAq4yGBsl3IyEDoUiQDncZIos7A3NtJObu1qQd0ceP8TVncwgD0c3on4XhIn8HKEnVw5Pu0y
mVBDKaIOsc0Zk2oQf2oAc/RG2UFtwxdik9uPgcjJd54Ku04siJaW8TrBvGQw7f/EDTce1+KtDI4Z
cNdDvW0NWn8H4IM0uER9vMdkMyWYdRGUUGp29cFCoY7TVDrGvVsSSqKG2mcEd2VucV/E6c330o81
JMlUgsJJsLRaJzdooWmLpO9XXPBeynxyoYiAGpvpFiLWF114f/kDwQjN13E7UMvEFExBn+Zq3zwa
yW67tNdDyECiAL8BUmV7lhuVucILvv3KvmNiinCwecrrZkVSeLMKcRQebZgP1YFuFuVzpFwSml6Z
Lbtkk0ccXL50rvJ5OE3H3zoaiV2QmHKCykk5n5h8WrXvCxvaR9++Ue1LdYY2VHEfXSoBM7BcuaLO
gNtlQw5efnT7zsitT5bYWgcE9Fra9yDLG3srWG2iRVrTz/6dUiI9yl22/dxTiRPNrgKmCJwYihQ+
lmGGGQnbFKFTUOf9UezesxcmjgU3mK2fx+rtGjeBSCXnaXs9GZ5wP43LIhxqejafZWjiZjgeMVlv
yyqDVwR22Bw2X8z4T/o/XFwEjc91vP8KIOfxuX20BIR060pJ0OjDCJ9StfYWfChuhTcmiZrbT4LZ
HfoD5cVrRbQR6KzLo6ioAjJeE04by6Cme9GRcxzeBsUCMalICAK0pl1fYBw4h0Qq4hHjYBxtUSfG
MhZaarl3FN6MTrUA8KWB3247VcQ5Uq7wMIzcuqu89Imkn/GDi+M5GWXsLU9s1vXbNWoPf/46nGfS
urOBHeRs/6hkHT50UloEka53VVen4zpDKUG5E31/g+BAHAlP+Q+1REVg2+ra5putUYjJ0xllwnxt
6n5DY/OzKXU0T5pwjySugi23UVOlWObCkuuLeXMMaiHrd/9+iFutzOVhCBcOhVmIYAYC8HACsoWN
ihvpY+ofUu4F4wOc1/a0doBVgtylX+kiKCdeUV4OiGCwO7Mo9mpHoyRgpAE8S3GZ/Uss1Y30CEFi
DttcndCCjP2maz262pc6mPu+JK3GLyrGKV2kLSA2Fe8/t6eNpAXAxB/MPhguV8/CEdS0U5tTt28v
Q9+0xKWAycRsv72UlR1M/kU+QS+EHJz4sg2vd/Pbvllq0IxJ7qs2OItml2JHTrj03afUPSnun2M5
UUGV8qPMfEIbYT2o+dguRWdEq+z9N9XdemJmLRxYgO9zZMTIin+EFOJ3Hem1ZuqNdvdRqyT/lpjl
GzGB8g3JFxYt4y51mNWHdYmyuJDSrTaxgHUOtZi4YMvx98U/2Po6jXSX0CGS1bQjsjpan9oZ7Gn3
Yiz1W4vR1QxxCcR1F/CJ4errnP4C99lim12X4nilTNoIkUdaVryCJUPyI3NkChDhiO0LFgssaiHF
ZPgaxZuXg5ydp2rZiWad3xjjAduQILJ9Safu9qOgObL84RG9eIspVUSiGDgHoGFTxArr1b/2+1Nf
wk0obXTwM404ySXRif8Dz31FWQAz254be083D9e2qWsEIQrFm1hp0v4JfUoSN/bX+2MjyqjTvkj7
Kb78IXnKoCt2RfqaYoTV3H2zrmkvJLCC5a/rhCd1ooqCPugZD3OfR4SBxJkDNwRk6dQbKvU14OcP
PHbcxCLkYedz/LfRK7mAwrvwBaZQEoHtPOMELSUU565mRr61PJJOJiN+tqjhR6l+VX0h49MqgK+Y
JmmvPvNj+HKOsFN9qY03CubnK3O//A+k2HfH5fHr0ERggWmjnqscEXzwn3t15/mrp71Ecaxw0o3P
lVXJ2r9r6VxnTP3IngzgMPLDItgten0nPjSd9dZ+/ACFQeUQ7VJdpAwz2r8Na9ulHLG7bsoJhyGi
h7jYcGkvVatgzjW5fzcxsKgt+L4cDAikeJkmBxPb28kKMm47srUQcZ1n/FGZsVJcb05jyEFhV/gk
i10XUPbI1Vg54Xd8G9F/P7hs1xkNigJo8qAaxsBruyUxJvjgYgDcUK0yorbr9wsu7LOcOMfOaihG
Jt9e3/mF2Q0U6tTLYEML1+nCNq3PeRLRT+6GcSBR/EAgiBHN+HbDWYrSD2nGPViPNeAzM8L5vYBL
cYzRRoANndXDMuVqPnRJXZucBOqbfXMT9DFhlqWyZrDKUAlXrBFC9nhXie4C26b8+US8X5+3aysT
uaLR2M8afe7r41yS8DFkL4HmPlCyWCsOgkDXKz7AXZLcUHTEAH4i8BApVvgSpLD6rgYRVNy6qtrx
iDL5/y6k0hyuEhlzqu7Y/QMdz0/tmay4Am+oHdhvTWOI2qnutDt57vjgmiSVFdLWnEpQOSmvpP/s
65mG7ffF4CuVRvf64exSxyOhgRpmnF5qShPy54B5xSTn/UDhB7NasTjV/kgwIADQ4sYW60lBMPwn
ezOmr+HAK4T/gVccIcC3IalGpzT3fl32MdoKStdEv9g/xODlTeDehaPGb/zByZY+MwSv4u3zX97n
lUYda+XaWd4ev91mF9H8R2KuLfNYAxJCDxakXQCQxwpS4/iduvtUcWK6JKse8q40Qxg1wTrce83m
YhMhiNXLMT8Tda7DAjgpr5uQ/TA2YqXvZkDYEJ50gnbNId/kknBkOjGUIBYVwNY7D8dkTjR/tQGJ
/3epSK0Ls5hVrOVXL336JUe4/daHPLWLFM+X2WChi62EMC1s44AehzAdDiERffXnQKnaxvM6mlag
xZbWkC99EXEJUYMGYnhwoGWUhU56FrP/sMnnMgFE/ixipBqZo1mLm3HwmQHrxjg2OJBE8rDq6Rqg
o71atlodNeH2BiLlj5kmYeUhfnuolnimg7pCSLz3bq9gP8I8rLMYPzDuv+5rnxKiDBrAqoUbQK2G
9gBvnJO3+G4dFme91TlXXg0xpHbbNGLjrisv79KV8LjM89tYaXPNELwvrxcUR3gbh88P7IGxSbAE
qrfmgxpT3m9TKGPbhqnBe2xg3GuoOeJtsLAJqQC5J77n7NqQZSD3WSsoGcJVLMST0NUu/9vRCoFV
ZLnzACrN73B2Uff2b9TvYXxv8i1+KsQfW7J+KHrRSaG268JPjpHyCJwVoWaMzLuoXJdVTc/Sbnw9
J74W1OL+gijexfvSm+Wgc09CUg9Fz+5VAuTwTCX1gMLiaiR9J7/mJu91685duQ2/gX7dROEM7vkY
LJ9Kpw0R0tMmAaX15CTP66x7hXW69R3Y8g2kpCIikCPVgXAccycQ9yiRw4X0tDeoGtP/fShci4JS
n5U5VcOO1bQF3c8SfuAhCMxBQnJCj2BIHleXfh3zAsyPxXzqgaNoAyr33A/GvkmYk689/Zsc7r4K
Pu2Je88N4SmNJ4zk8M6iyRpKhIedQor7rMIayAL8UC3BWS9NfDnrlJFIxXi8wqjZPN0ruHvZWg9u
3GGL/AG1D0xltSd5J2X8QoI+uJZnmhdjF9DA95nG7DN37eu9LSf9K3U9VEXC2SaFF+4cMcYiNvj5
XwEuip+uOYOW6C8qD8B7zx2uzZElrJJTIf5oRTCWAveOxIhga63vrTND/fSK/NlPd0TFClMSKI/z
7a0Yi0kPGFdwBhCodfgZaNeggIwz3tcEsBdesXdDWpc8G8bboYmQwlseb7XO3OSHYHfCmB+IeA0u
IfJebNLWmg/JvI9SIzl2aRLs96GzZjzC+on9k10MDxoDf3Jvy1F4s6FqApTFk/0WU+pLYPOh+XHk
rkBjh4Cf3xsvUGto7eGXD1Rr0DNclksgvViamhmlSP49mVfSvDzYUXC5PQSJejqp8AuuezdmO839
IpB5emNS24QMd1Ts4CHsCmhFcLZ1Owh3UTtVlfR9/QJA1DUJuD3IRn2GAT5zPWlQDQ0+es2wYFnL
QT1aeGQ/yLVCDkLG5bCkLMqEofXECPx07TdkuY4ufPrIj7lGc+8FN7qfMvi9V7ppkp2zU+fwcAvD
fDYUm4PZY3FoU+iGHLRmRlJR875+i8RsDhNM8Xo6SCIpGIYbFaUhUxEj5oESijFVTRNpakJBzPvI
idEXb9E8Jk1brIDIl60f738Q6tj2pidcDVa17iaNTfhBsneKCLsYdDN/adxR7ZM2aP2SEc5GQNSW
3RvTUSIO5CZtfq/35UxGFQ0sGyfAgmuDrR9sNucjrNEIYghWuN3MicV4sBPjLNNXe9Hve0YhNup2
VtZe3X+3fmNJZQQfCr8nIGTFGW0Bex9c5fZ1Et8g81LEVNIVsb6xx8kChwj0bUrqZh9sCSpsRYIi
Cyj6hze9/DA/BqTWVMdjzj3CYLRRVYhab/jN3kdihv+wAjFdRr6GUJuHyaaCmMFWWxanU+mIRCS8
C42WPXx49zKDqohO6zcFuzD2gEindEbGI/QoFbNAXhB0sTcICPF8NKRTArjof9dXhZJufXi5Iy+L
MGPH9mvdRb4j3sn8EzbCp6lkEd3IWOuDfcyyPl25iwyAW+JTIIGfwxZEOLB+SzuX1bSyfVTYrYUu
2fYJZNl3xkC3IAE/Ro5gGNRtPCJAfU6kJNuFa/7C3D/KymBUltquLEouFgxumY8u/1rz525QM79S
zIuAqzVne29GiaEESibzGYzd778okl9DNWrA660lVtEGboFA6B+47PJaUuGz2v43HHlt45LQii1a
pXbevKef0VxgLlMGNOfuw0it6u+6YXR6OHDQRCyEOIen85nl99Lx+Xvd5j6wcAFm32h4x444IxbB
oA3II+RXoCM7Ziu+Gs9KaCrAEMMyZlPL7HDGsj/+6vtR0fLzoietblx6NShvds2u/1v0SQZvOO8z
yXT/W0UAHEIEksgd0e88S/nRPSuNZ7XnAQPIL0eOZ7T5NZYct4mOI6PdvFaKbmt7s6EHD0IAmfrw
Teb/9QmFyV0uVVV0kWRijaSMdCDT4WGVTPou6UZgLRV3Hc8fRrUjWy6+hpY6zkhZvaxHGvZ8bFdv
RRpCeFCksOpmqS0bu11V3UKB4zf/pYZ0Qd154ubkb4aqzWaYM1lFu4JwuwJL9ek9B7aczgs4I1t1
1ptMLBB26wbp6bNShRBUEV2eWOmQzE/Sb+0F23/YZVQDPF+SOVoeelAOTLPwdHazEdoupuoFxk8V
2uD1OjeFsi+Nlu7eSuVOy/rASUcaVc0H/lvytduY7pQi4R4CC2+744fTawApHdfx/PbM9oY5j+Uy
Qr5XcW2WRoq5gvjjgCVROS+ngRKc7adSMuC9UMz2c9UQwem3VeUjLa1he094Db662fWvUs+iycY3
VxTrToBWYbdhnUFgfZ+pmRmMQA3W1m/ifWysktevc/dP9hh5bhKBoKTecsUB2mwyOYYjV35eZ1Ve
c7W6Mhd10T7pAdv5dY/G2H8TPiD0H7ms4U5ee+DX8m83PDpyQ2Ec6hBLzuv4O7nanz0Zv2AM0fAe
cUgyT/rZnq36U+5K5DaWa6TM7j+Art5ETEhWe0O65TOiwIIO0IcFVVZt1wvUZKuLE8jo1Zyw4dxL
VySx9+tmELfehDzeShg0hX3lPMmYNIxp2l9/aMnBth5UaNwNSV3jmxuziijyWCWQW+l/UK8bvdgq
0si56VnqbM/EMTFqYwQCCVo0aKsySZ5nCRwYDJDsm8w54w8EQSIQPQCij8rE3MsZEfRExfYHOLwF
ZxvfNA1bF7gIXC4YJw8dAeqRwqsWGZoJBNoxPVsJW9oRa3BLguOPzGwXly9R0eEBUoYz/aayu+Kp
HKAxchVEdwyXzFbRz38d99BSZsu+Di8+YGtp9wTihtl2uFwKsS5tPTowIRJxO2EZ96EWXPUtDi8p
tz7Hr2vOebHAhmbdlUDOl68EgbvymKP1q6vlHrgIqEJgPE1ytNNS3OaP4dbcbSwPvZRpg5e7j8Ry
QAQ75tMlQYspQdeHIkm0ZuQxcq2ZE9iFwuOK62rXjNNr/bzW2WVpc76mRPMqFILTn9qYkFdaHtpC
6Fnj3tbXnaXdj2D2FxgUzDR+GIvqeegF86Bt72GI0+uRhah8yjlVguC1nSobwIYd/EfTyo+lD+II
oXxz0o5H3CeFiql5URdLHzEqLb8faeh0H+F/z9QdXXT/iOgRqc0J7CDDX0ZxJ5T8TKpw13gt0zCd
4BOW2QthSNreCPZnUSHROVUuiBV+Fi/LhklYP5KGiMkngllvl1WtPKs67WY11g254HwEfiXVw4Ur
3F3SLuxsL2RMOC1yU4hfvPpaD0LndFcTCUjQpQcLJHb5fT48vITJF/iZahNPNQmGVWS8cxug6hnb
XsaakYwXeJgtff78PZZYT/zNskwNCNygkqSnU1LvldZB8d/T9Irfq/+5k5psvTZoeFX5X81e2+LT
hjCzy8l7/RPMIWwhf+NSb93P93n26Psy8H+Yl9g2v4UlO416DQ+2NBY6bMjkVieQuu4kpnzO/0YI
93yB6OQzpNSoDIeaQ8TEgB0sBdGKFwQu8Xq0wEHVUi7Y3nLBPf4QOXxRqm0DoAba6A8VKf5Qj8kg
1xHXtlTsfaZvBZjPSx107eh2eZ2WGZVpFdqYfOReenp4Y4Rs4cNamXryM3Yl8UKeqUTj9UFLZFYJ
PLczahpuSSB+yes3MF7JxgOY9zikZ0GOSuafcsQBRcGnvObjZsvtz95Sc7pW88uxUVGWq2fOMWWP
cpgdc2KnbbGUmUqiu3nVTIQr23Keg4SjbxoOym1eC0miDmRCcC+AwNh6bkCgurc1Gvk/9vrz0gpe
IHLzAcyTRbFZBuf6e3S5EKea6abAxBcNse5TspXJ0S0JIxK7+NoKd9L6i5e0sARntl3D13NXkVIL
DcaLkN6hmiL+Xb8+z5MldDc9F9/vbR3FFJEohT0BEYIpkrKNp9SrJfHjBrOD+KAzL3XGs0gbdU1e
4slBH2cWH50jQI21VwPEES2e0Hn1n8ilrgKkZK0l6MJNTYOQJkATIJdZA0k2oXRsXG63AnqD+TbV
geZYsISBjs9OKi+AH5RdFKIw4Ma22SV08uddFgIFbvXorW8JHQLsY401AhVXNBccKt3HTSKSzQ0C
Wiv3S9fkbzWQMfkFqh1mjuaiqJ7RTeWT3WBR1tHH2OKc37B24cvxOMwk9Bb23+k5ZSCFSK3Y8yPx
jorqM20ii8FQ2hbX/Vf4M9HFGNFmlGGT2l85I5WBMyM9eVdhahu864r8uieiLXbnqcrTJiwZAhcM
kTJmaz7b+94UdVjTrcxL0bpagsOUPK/mtOfhf0HS5UqbHjHcFKPnBHIosgJSP/ufqO797C8YbsGQ
kbbHiHWj8Dh+b6wPqA77cYZZHBU4UQTfnjsdeEEALzyWd2S9uSTlv5kawVIzXLaMaiZVLUpS+af6
CY0EP72cGPEoGgG/a/4NJ0ZNbE1S5163P2gmMLHuTs4ev0VA4DE5CnTr2KvQd7aJCv0Xy/p8dTWH
tNRd+vHYqkP85PAwWJT5z0Wm4yYNYCBrVEfzqwi7ZON8XYXuetXgY4n0sgvY4u08V6MDRGVy1VRw
T1wcy6IgarZLblhehWjWUYtCkxSuavx9J8LRXCsXonyFlpVFujs8LFlSoeeTkRP+trFmqC43csWB
BWjCNWVsq+gQwqlUXg00HCKnXNIrmpgZHoHZgA9lCCZZVytMx9RSY/0QeTpG7gK6YypNO8V8muX2
4Uo/yLTQ4bsD7gVyYAUh61GRlxZR36hcRaA6K8QWti4cg2PHCLFKnFCf6gPSv8N31YMkwJtOHYU8
9LO4dz1T7x75mAkG20T5mdfkiS/3SO2KWwXx4Ceo0yD0zWQTG8IX8o+63esEhXVrUcuhLNDJXafF
lc3hIJ4KDMEJ75Ud+nLV40/jC2cWGDgAM8nZMwHWA39zWBslT71rZSHn8+UW75MwrWKAABwqLBtG
xjXKDp+KCLSHj1jDVfkK6uXdBoWA94LUG/1RXt33ttAlvKyUIc9Kv14K21RYddx8u4N2eef4G5ND
Is3FVczc8g32V1OrgeGlG3FOUTAtN9sfO03BGOv1iCC7I1JmW1GPZFwdq7h0YeO3SglQq4D9HHJ6
/bCp90q/fe4WkQMdjcBy5qPcvovLkoGvBznXgmPHBcHIwCWMNn2weCbNsLPkvi79zsHLKTZiI5Nv
trc2WGLGOrnZltsXHlWNw+WX4pwQsV4c2rbT4NW9ny70xBDQ6kA8cwE9c/VA1UnSGMYU72mtW3Xr
Qg1Gd3/rB+ZELYsYhYfHESHVTg0GoNwILdgnyrJByg6wcFLHxBKRzNagSfa3Hk3qXOkIlWQDzTDL
UDtoloyb5Da3ASIe3gdPIbXGFPiBP35jmIzTPouiKJ6BtHo6C5MkBpE/lL+GKyvXolTdbMoK1EUu
M0ILHIZC6GN1vV5JmmsLXqjlWvEZ+X1+m8IZwg63I/IqXraJHCV5tVhHaMhxAGJtf4swbYtHgPGZ
4fI/FCZJAuj8pTzcqiqBI5TqmvP+SY3bsNukITn3aPyHCkUvg8hpiI3A4cN9yyEvECh3cI+rMN/t
c5BZ+e4ZE3G/0QnlKuBCWrqY47tqXXmRZAixcjAKuhzfwnHDHeb9RmJA+28wBBmk9+kjsn2afjOW
86LUxFd8GbDEY5T7U/+9BV1dz3CcTdy+bcOnQGJf7Ah6CqfMSJEHTpX6+omz6YSh2qd4dz2c84vl
058qQ9NFMllexI8gJoGfuexcDDCWCmu+HyANV5KJvreQPDq9hRxxv8tHOerPIzqZl1fOhAvUUeXK
LM4JX/XnVY+Mn3sacvLMHL1sZUcMQWOnKbstp5ZWmh5/sNxwLl6th4iXD8DwfNsiogdGvER2aCqv
CmgpOdTDM+oqaZmn4Nma/bWk/aSA7vNDxm7EDTUpMGu2RklsETHqVKtFcc/vBSerSXWK4C8Os+3z
5dVU43UpCChMRTcs9dgS3HUyMQLGk16YXitLkQrgLWGriNFxdKQgbXhsZaR5WRqwcwGcLcf8Dh4P
wJhRZx1cEyx2/nYV/8jpdKZZmmGtuXrIPMFg1SpZl4sQrLUWr/7dhLDxjdWYC+lLPpkx+nfEJgp5
WWbH/njXYNrpg6CGHYiEgiBYYytegsGRiXNDt8Ypemz1EfD8fiHWDDykMlKPXC3fDLFniMwyGNFu
dRZLGbbDKAxh9/cC0zW2grGTmacK7EB2qTJKXXG6j5iUwXmLZzH/61ND4EWDcDe9V2Tjg2/YQq6D
VLOTqlfNUSDjMDzaRDufQm0y3EWJqFwKvsjZHJX5Jp+dqHooK2Juxu/eIttkQzPl1dFY4tS0GvH9
2U1pyq8B5rAWUX4nlvDNONXGwWyvI/3CA5SccuqZLxGy5Fey3+q6U0xIK3erb4g+Uy3h1u9t6Yby
rmnA/bntojCJ5dRBinMJbcNhiQGa8BUg6SnSvncHwjGtBpd/tUO15/sBpWfd3V3WNN0LXIWq55SA
T3MB2rVl+yaJJKgKFTgcWuDpUlEcVJOd0R0kcnLwUWoWmPOb4XczwanOIJInmLL2HOec6bTlW6vm
ya1yWSfNvs29jOKIZmc6uBcquMqgUM1YiZlTP+jlu0PxXuVyZQ36yktTNoMbQGMiAFCpwRSGC0TB
sdxNCfLdTWFbx3mOO5XDrEblmz+tOzj6W2whLBvMNZSFZtgFbrp8gjpJsKs/31cUcalASwebBA2+
ckbjLQkb8E/C9Dp95t//kWW72kHwWhZHYmFSuPl0HCKsxWrS7q4DO2t15LHrhtlAcMvtezOib1Eo
Bf95TTUKzBGyOesBhd++livnifbZe4B5RRSB7s14nfgbIhwzdBwCyzFFVxjnHzOMJ02OqJHqvMiq
0vnJQ/U2i42LlL/Ctna9e5julaX80ghgLN3/rkseBkYb96rXldlFgz84gkb3mlUqZaQjEawz1N91
4nHFyMW0xd0KwV02bGUFPaJ+stw8kNhSfjBH9osGZOXB08LW45yixQ9LKpkbws1cBEKh3fdYp49A
l4EYNoKrjwo4iy9xaPZMk/hvxAqgKFNIQiQQXoJhssUz6oUxgFq1M9WDpRw66gtI256d4/EOxMBN
bPh/FUXj6M9fwI7ral1zk5lahbsOZmQ2MCVq0JegawcmBochLpgTXup3MkpGjDtrl0ViFPH/XdZ2
03/XbPPM6yKxH0n98grxQuh2oOWIqO4WY15k5qAIoNZ5nDCIpf9HHK6Tbj0dmuoS0Bs4DrgabHge
faSfu40GP5zGWZWeXpjRlretKEb/rj3MzF6rN16F/Ek3OMVc7jLggY0p5ySbU41NyoYhGP+2TmS0
3nLeJ8ChsTj92e4nC09JCdBWPRoWg7jyrhH0Q9HVo1eyI/ITQZ8lN7wQfw2BlcbGGXY40rBqTN67
6DttxZZeytd0//KZN6mFm2vh18cnPIjfRjf6mrKdLObA8wp+b6C+UwH1Do4OOjW8QtIogcuUEyS6
qAY3CZCWbeHKoWpL1vLYwz/nsdY2l0imtR0rXdphO80wMVgE/YKFG27LlEoX8la1cBhnQTr5xyRf
Ctev8WRwgK4CLuTfKfgzc+xk9/VLG+bDPn4qkYz9eGSjiZcMg4fqp3aplMDM2breLSJTnrMPDDkL
vaCyCPnENvZVp4s1Xxf57U6t+kLs459FToXrhYICOQ/vxS7ynjatsUjwZzZgo02kdUZ9C89zfOpz
Q9CWBjkD1T1cAKbvmW76Yh4m390oRqZN5jqWMnELtKqmgeVNtOfcNXqqZ8HFz1c+XcJEhpa+pDLV
YEa3Taa0W09vlmpfuZJEEkngTXfdhOQxUEjZt+KOb4yy+a6toOZYI8UPD6UaBnDEB6k6ICQ2ZVEo
UNtgNpzLIOpUdFdC7AfVPjP876TKo4eXEexPydpmrSPHj/qAp+EavaeR8Z+uuBdC+XSHGgQ6Xl51
Trpoj5apE58PGFD5b1n0KGSGPl4BNqf4gOS0tIC9fPqji72qu4zVqqLJLTJCCrWfG+CwhqCHCg3f
2QPy63pv1l8TUV+uqMbcRLeRV1+cNYrcKyPW8Vzme0Ic7c4LR/RKV6/8ZUG+RUDkV+IaGzWgmIya
Ov01ee+wY2QswcCXrqe8Bamez2S8fV5b+xud50DTtha27mNcqxI51+Wb//zYyckMtZa/NI0PmJP8
gjX72Dz5FBRU7C3mUcLv0SS/JSY/B8Bv7JnXiNnkFto8FQHmqk8CSeimZtyK1LjJd84he6fs8MII
a5yzSMRSGX3fTlBp44vESbN4mN3VrfztH6xuK1Oa6U0ksEa/4MHpjSYTlQWcY3p2yaKA/U+9iLz4
ZxPeUXxxwD3OZ7N32NQNFgr6WFjYosOjxFeb45ecsiF8ccb3owev4E+IDKGcDZCXNt/NzgqjdKbG
CkXdolSLp+YTGidoQVXYUICocYRyshhzH/Q7qpRxOD1HSaGuQ5o22mJl9PTGuP1lq2Fh0Yfs4J/K
Jy4MJV6XMSDU+G/LBhF0GIkL9m5qTv2tf42x7KCxo6hphcqjYaiW05iIG5wj/eoQc3bnz+cvGmR8
6OxnlLKnvsGsRUcV7E8j/IexOUV9ex1r3ESLraYtTtsSzJewG5CqjprUGrw46NPhmVsw8fzklFd5
DPqYJ7af8wiX36nMSS7IGeGk2eAcdi2xfgjr68Yf91m4yPvVaGo+3nfuBEgvQlg+It/7oGRkfzm1
4hEdJDhXvtg3/ZiAJ/ronmV4sZHbXR2yHhor7zsy99rnFDgvS9VZoRcTA7tYU95+lfu2kVxXt+v0
MSYquqT81KzbBMCl2/OaWwJQkbFSe0r/6clyZcQ843H8NjIaBxda/I7vCdf0I1vtkWjfbZh+n/FE
mu8nKjMHM8OB4QW2gHzGjsyg32IpFIKaIJkYt9EWqT7yoRxvPNQX84JHqcF5sof4Dl9CuShkWZ4e
hySAoyEu0UzgIx01HM4A38RYRDSzrbM8E+YPShjuLYYiDN+qHKnb/K/le9fAVOtF+gxsgCxV1sC6
oXHeJYeYsXU5qzR30D0cqZ0WEXXVNqMR5aZdPoPCcDDB81Au2rogdrEUEvlutWxIBDOXXN1HNEYB
5iaE0rJth7Kc31HxYWfgYK/+S1jDMA29g2EYz6rtJ675kImJ30NYWVyotdfWBtyJGhB6cciKE97b
J3EbkeDTrVNDNKB4SWri2mEVDy6z83TMjvi+K0hJeLKBn+KYnolYoQ6WWMljrOgcOU2Hlkw2GncV
RVkf/49zxfeoZFntFJH6VdLTOHZHOgbqYY9mIuZV4Cy72X6uKv30OOWlpWjp9BOoD45AtVRjo4AZ
VpiJuGtrScHwAdMrP5cpn+6hr3MlJ/28wHs4SNgPoQL2juES2YCzJCU0PAojpXKoaBGBnSfCtuJs
k+Un5S5nyGgE34WtKGDVeZv6UFBDFlQLanCI2AradqtnXFKfIBHxRcr7Iz0YBAn1xlbunx5c3BvB
zaDxSwLPccBJxteWn+2z6KgLZ5JJTrAOSC9nBmCAVf56vXymYvWzCBiHnuRGh0PKbO2qrsxAr7Xs
Y6ulLKfpphBmLA/NhXf6DQlJOc8AoB9PopoiGqX4LesjGjhrG3GNWYrMVKYzV/zqSeTljDT+bcWz
qVLubnTcvo6gbmyxOCVNk+by0IyuSzusrq7fkPN7YEoIJPkegA0/eCtU5pyQBoQZ8yiTAbPz3PWT
nzKylzAZJIAQWatxN88nuy4ryTuH8wVeL9muO6g/WXi/96HdL1tldq8E4iyDJBzl9SGUPE0q+Le3
2QlDOnsyCfxGAhTKUwPM6u6617sFyr2xxDMnNR25ElwAXC5fAj49nAbXKEEsG9m6FXX3zKi6unfY
jUWxTcCnJBELPcWH+JU7b3hmq8Wh7NWJZ5yaAXmjv410ZO1WnITurucRlddp0dyN7+n3IbQp7sVm
WyiOycJ91t930WFCnD/DUxkrWngLzeQWJk9ognI1UlBi+/OH3rzUXgcyGShIllynb0jAgtRy/+zG
vHC3O9Ctb0Xjm8IqJgcofbeXhRcWptCKlpIcgSDu71sIwsu910R8AWMtPglxzWwm03RlW4E7QCSs
+l6uEBKNHFJcrk0B+q3N7DKFRObS3qQC8qwk5T/oAjD0ldrvxunYgtrU/RZIGlMbPE8HvrQE63ht
YrR2ER8/yZ5PVgHg6+bNDJk5IPfngAA7hmgjzsKoYAliGnVPQWYy4aAQM3Uq+Tmm+YJI3V6l1Tcl
mqIYr2pyrUeZvoErSbsnj1cJ6/2/dNobDkXwvrx/ObA6F+QhRxR+nz1HZMtB5p1WjNS4daQFdxz2
ydsUikWkNZj22yNsc41G4d6msje2FJN9iw3keOhVAfCGgc8YO1rA5ovZ6x7RCx8bAvtRtu9/z55c
IVFbTbQpA5zinMsRulJVFbNKb5BmtQyBEHoe/7trxXuYJxsiLOnW1Om4EWX4oTs+EuR52gZ9uykT
7FK/sMAJ8s19/cX9MIKxGkp7K80bcmRc0+zI2vOcmskklEuqc/DOHZios4SrMSYuj8K3OSXj7v1L
G5EPxTmi3X2hSMDye6KphIXqaL4WQjY+b+Q11PxoH730EjjI168eobCzjNaC+Cz8tf/fumDprSjP
/GK1VsUcrvvKiQqWjhpTcy3dUSXX88yEboeIGHS5hIlXFX7QJyIJCSLtCLJa016Ww0/IP0Tey3H9
iZVGojQzfCFuOYF8f4NxV2QWzOwDOuRVBj2iG0h8+V2oQSv7XnNL55WhsBN3HXY4IgTebZ5xuEqP
5vgKOV6yFPTGVPezzZPM4KupJiJh+g6lWsoThT5/2NPuDC9RbI/grQMf3cXIUkaEiV7cWWkRd6C8
N/mTvIHmJcBzkoBJ93x5XK1K6fewpQkvNVduHExueDpM0Wk+jKBNLviRWiUeIEiFpJEgTtOcA1MZ
DxpsqYbExinJoHvJFhnykQELEgTo71i4p5E+2EfgJ5kIEQnOtASFbGNMQs1zmnoDeRTmQZduz7sT
Tke7/2WXjnnD2bCopvFoVXbvvmZM7SUS3KS1yAlVbp5OlqV75hsCXWmrxdMc1j/8eyzbD0Y3Hr+M
LNPmdOaYaMStz47qouseiLaafwNvuVqFTlZjJJgYLud+Ss5p8Isd7ojem0L72rOUnq51/1GToJpu
zRmB1MpDWjwJ7DwsdNBBUYmmg6nR80hnQCXE8DllwttRrLK4+auUJ396i+Ey86/sSRMwkHPX0AIy
Dc/tMTZ0ynFenM9dKsb7wOF2WaDGVrKbozqPwRHhI48qHZt8NQOn4yj0abFaHl1gMmoz8FaTlq5J
5f4aCmImpKjVfvgCbZd+pBzerPtS5/nwD2EK8ANHj2WjFWCCWWJ1vp2kAGJqPiMoSZwu2TazPixv
CTkNqrDNyVdgAK9o5U+5jIlOkCPZPuSOLDx4IFbc2a5q2VYTPsxq+2V15IuT9VQQi1a6xPS1eYFs
DNvKMCQmCUmutimHD4FqbCWqEGRHt/xAfQKQVMf9AbHrULBX2dkY3tPo2X1O0JcVjbBVGt83ffOa
kTQ8+v4xYeMcWzLnblmnfVPUcLspj8oPH0GVL6Ff3JR60MvIWzbUsQXX0skxpcFeAP68oxaq+2Il
X5EqAoETDsAY7VIG7R5FeIy5hNEFEe58u5CqWOZgdJv3J9BkFpHQGLoT8PhuvV7jBlDf7NESadGa
r8j3ryqcBblucH5/DmZ8A8HRe1J+6Nl287CSU9KVQTM9WNaB2+DnVAHnuOrICxKCM5l0w4baGQmw
fJH/SDolmFWRe1HLEPgzdSCv5KyRz1h1LXaOVDF7AS0ArG4W24ltBmWDRM/0dhzfzUN7D1hgHwa7
V7vqcNTxVA8Al5afL8nHPXeKRL3wB1UuG/Fq/FEe2oNx8muGVDQUDEO5MsJpiuk4eK6CWDYVt56o
NqWUXdrhd9x7yj+U8gvAbYW6t9NWXfSkovAmp/+Xxz0YCUYTC0s+LPMgHKnVu26wornylUgpvdyO
VEyhB7paO+mvTCmkGjcR9VBUxvJ8I0jJQ5yYdl/suKDMY0pEKEPB+gmSFmpafg8673V/yuACd6s9
pU4FRdbf1E97hniDBbQX7gy+f9HjEv6ZQ5bq35MKeqUgSA+XiVAxk4UqLNcmo1P39OLkJZCCDy+x
UZgLrhXKTKejjgvxryR5AUN/mmzN/k+kDJTBqZmgJisISYklea6Sqlkhc+1/BK/643J5AwIseDEC
rYYibaNQHFRM6DB1VffPlOSFp9tc+pPFHloHpDgCLTvu1paQCGTBP0Q3+BpvT+IphxBzWv9DcsOe
9BOY0uq7/BuSgZP4DbRxyR6kwVHdE0Lc2g3QxhBAkXUiQtBG/1cmuBN2ppethfamc1WOi8XzodkU
EQLfwiI6DWPUCpncVUCx16fhlpDgtkohLl1m0BYsV7+WOuaDaUq74l7Xd3MK42dMp9HGJEzMS65W
zhXKQhxlhO4H43Qp/8JopTHmSqayssCbyN/YwEbndlFQ1kh95CPNbj065ulwaI8Re12kumr+vrVr
HO0vhflf6MwifzQE9V1bOXd+AMFA2t3CRJswBOdHZnyiBB5w+LeTNuTsURaLbDiwXt+IKNd++TjH
q3mQoHmPpbE/nnzIXezNSrJ3g9DBswhDrThdE3EKSBklWdhigaC+bvIzhLlYwxRM/tSJfVdGDCRN
h1SEenjceOCOq+TkvNmXHuSZBXGiMUCN6HYN4I+3YXUgMuCOsqgGXjE9KkLlGJ03UkEOUe3YwdPz
xqX83CREY+Yl+IvjcoMNaCPIMXTUo3Bi9VAjRReHvLCwN0O20u/DFU0mjjhjtZttu/gRHDP6KbHF
rXgYJnrJVoPA+u2ivLlXHmHdcAs0tzGYV1iS6zIQQhWr20yc9oL65LYCdGzeQz7IM9YzUmH5fToY
vUQQzI64k6VdQr5rifxnh07hSLMu536c/SByKyLK6dJLw7966dKzNeR6WMTLh0kGEp5MXEz6cNw7
H6dCZRyQgMuu+0KjLzS079btWFcaHp4p/4I6yh5hVfsIJKRfKa3QnPwTeYgZWqrD+gjUZM5qoVi+
v+rwMf43dY0slBr3IqhgXzzzLIk2citbczoS7f117sQxWRx1CEEEmfKRaGMCD5sCN60c6OToGgtz
9MDteXZNAx5En/rMuHje53hVaiik72ZXuNHVJIWq4X4uZ1j0pk+iOuW15rhOfSP68Zgj7rHZl6n1
lzTF9ipC4MH5UdXdwhXUr9fNp/QJM25hHJrqSRGiVndnKF4UgAJnsWjppK43S0XVhTeNDJrkvqv7
K5FCToRGIRNkwuR0zeZTHmYGzC7h6Evn/NysI4uHT9w8KndYbXO++V16l310iU/l6NC9ndZbW31p
UROzhSB9UUY+dUgjYm0vqoUmQjvc0nG7kKEOWvpssBYs283h8YWeJ0sgzuy+8M4OLrEDRp4GElHB
ixQxwL+HGMBnsA2a6AY78SWqucAaS5St1rxEAFMSAI5qQ2jhopJuUP1MC8+rfuNA66mi9m1hAr3o
yPGDXEL8T6MRMZHd7PLSQLDP/s0v23jFWLyy0O9+Td9w9IsVSMOoMg07nkpnMT7B8ngclbrWMKDG
hMrQFHyiWCYF1yzZzTQVw9TNvhqnUIszvVe03xKoY2zohHFE7ON3rG4Fo+9WxYV9fQ2nUXe9U0xY
Nhn8m/zO4MEl+wvfpAXT42kHa254dFzasy/4+zUIZKIpw8vhKua1TeRaA+xRFhzCzEytn1H6oydA
bpjj+l2hdo2lPb43mHic/k7m2HMAAilLWT0hjeox4IHVK/W3udST4aVcG+0bP2o+ECAZfnVEppSy
q9KDtGdWu8GDOHWselwI8CPs8VdWPqdPtDH+7Uo9cPW5VLg4Bh8btHaQ8uZYfC8S+Tbp/gBjBFFq
b9qzc/kYfmc1LMslavSL0NPrJkRPhLgkqAvDuP+ShqQLmMArOCvbvpPPb2qpWNg+Cvuva0oOzQgd
gn2LzZK1QRe3OTjHKrzmAXGEdQtX8rCd4b53rhVYAqLwSVS5ckFrEZXjt9jnWUMvEjbaBB3oRAdc
rDmaSZk2CBLs8BNUV76LIdttJfAdhfjjpVsc3dctmsgbW6YVEjd26byvl9Ax6Uhd8PX5mkCMvB92
qCU6ZZ9H242SYI5KfEypg5u40gexpox47q4DP8x/LeGPW0yluuLciaH3pL9KLZe4O7p/rOhui/s0
lkjYzwhLwhU2A/AO4nCKGGgr4/B19mqXhDG2w6MrAnzhwjUOjColRGJvS5FIhNJ1wDKQ4HeSFDp9
V0CxFFndezKW9dZre1uH8ELS/1+1rf7GF9icrhF/9AMTW/rqbGvzfkx8YDa9d47aJtnZuLfBYFqB
a9T42UQPaFuQzo0XTebUAW5y3VCgHT6mxDv8aEQW9k8VKGv+nUKlsg4risFdehKzgvE8xtxKMMOs
KFnptaIeOFF5oZRh5psd0gprvtzRtEF4rYsiArYerqFmAM5DXyJu12cIhABu1rHAtDirZoGb0INk
pUBsFxwwry0fZ1g7x9umWY5mqsyaH1h+uYLWAuvXZT6bo1oEptzoZXbCHREix97zCkoZ4lbWF8OV
W4sIOfvZ5m8rXQ8myCglLwMSlbDasp44crGKMlNDd7u9ULj/OPoE2xOB8OFHzspaaTCNfHTfdeMY
T4uQsc4KYYtGdPjsaQoTzGvd04ey55kE1mHwo5BZnWaWsV9nNGIhiNDQpz2EN8HFce+treCSHP1i
JLxzlLCwjE5f/ltvaKBYelfh4Xe/LHlwCjKW/nazQ7Fk2bWmj5T0ne3ZqmRLaBnDQIJZLdF/IKuZ
C9ak/1eBezvqWaN+J21qJ3hENZjcEOTi5aQjr6I+ZAm0ubYUdMJLY6VNjAcJh70nKmxqX7m4cG7b
HMdhuywoBlwmgwEjns3mP6oWI3HaCFrAbWTjcRnWykOLSXGroP+8l5ZOxPWy9WI/Pdm6Bc85fqaH
f5XqMdxml+tI0UO4otZ4IvOq2W6ePcx0DayURzdJRQ0/ouxeP0o0ameScwMNikq6hQ2aE5Crq6u6
SCK/3mRw2WzatWkqQFkVPlD4+3sDON17A4NBW2v178eQ4l6kacVQZplR38kEKGRGvOS6eAazvgcl
SciFKt89gVQUMWIyq3XzlC2K+FPr7JtR4YvQb7dp307te+dJ+yBhzs24zrXRJZIuXgb1DQNhIoqp
X5RXTY+ruWEA/nGe71nFCi+smSQB4SSFBOW7Zvq1v2GLU0LKvUTDMXBYoEMnyYHDtedsWol+j4Xx
BaHxJqNz+064d6Qyt63yjELCtaVKuTxfNwIcrAp3Nm9f2XdTUA2Dwei8Wf0OLYryHJBHl1e5SCxe
qstaQ6No8mA/2TXmpTJYFnrT1izArJcBH1WduySC5/hyQ8+zxVfq/Piz+eVGpacNqKXUt1gT/50+
4ipulYes6s6LY13VxmoQq9962UZqqgBXQlQ8by6P+dEqTQtkuEvwEqdDvQuOZ5CGexJZF67aQ0Lc
gGXkIEWNj1LsZjWSO3ANH6HteKoGhfD4dRnWz0v5DdEEe83qDqmtLQVeb7itfHm4UXuZAh9t3kRO
m8yzmRbiXEFp2ZyMXKJ0fhaW9cMaavAb3pAQo7I4ihFpoXPV1NVINhsdV55wDxdWoswWBOgyvZlw
ONOaouK87SWSEn3mTI66QlyQwLDSWFAEcNqCLhgZaZkrezkGVddXVcD/k330ZA8d5AKXPo8VMEYN
uNNrfZMxwHNPKIr8rSFVfKeH+sCp+/qFueuK8FHDixp9IlD7geelrqVeFRzXcF/YdqrjUL5TswpK
BFwI6rErd3E2xdlclCjKKDLUq8ATevr2Vmp1CxeVeLx6k9+9WxIiih1O4vHdtSxgRy3ET0q29nu4
ttV7c+DkEd5mIeg2Nbulhmv9iP0wqi0bn2r++YfwRdg1kPAa8SLgtEG0XUl8e7vvpwBXvT/mbqlI
LaEs1V0U3x6HmdCU6hNpDvaOGNC2qgHSqQIJ6od2moDIZJeR4t5/yCArjfaoNDCZwPhwX8t+fgDh
5DscQjOt16/mhOuuc01BQf0Je3Q5XWIBA271CJXmT9o1DmLUGJzCIZu5YLpms3eB0HiIuKw6UVza
fTDvcSVv6tpOgDpRJu22qv5Y694ybQWad/Poa7/Tk6BaOFWccR6NqngfR6Qm5CmYzzSQA49lOqP9
XlOgIDZ5icm87K6u+skj7YImv70rZ5gFQ6dj1vM8g7DYbHfWLzgpkYFFrHauS6ijhLS+unXCXWRT
M6FB1/zXkMfze7+JoS3/GRAeltukOpYClAdgJ3ghraSdc7XxWE0hwRZhx4thN0JecHV3roKPKwug
bAi2rgQELmA3jwNIkAkChfvSfkUu0DuCS+Al/2QKPJidpYEVePaH5+uOGqFXvBhYDUEe6BcT/Rpt
VZNEiRhQecV5G3B9INR99HOn7ueXbaHfDnk1BnjqOWcfZT0SbMgQuL9D2SSOofG0isnI3JM2SFbK
7iOnpS/y47xfssAROZSiWZM3daCm/RwwhHkJrD0S5hAVsYs24e+9ZM8Yi1wnY/uWmcGXyC2xaxsP
cBPECsJR+z5iFJ9IViNNUGT4o62Bz+Pe7I9q0vUG1EbfszWdFE4cdyUDHnyyOktOUKLrJIdBPLdg
P2zOesqeB6UI7UYysd1lbZWH2SzrxOqTo+juPvE97TeockjSjhumsG32Yt17TG8AG3o8jDT+0PDF
+ql48fi1J+85cNMJMsrg+PJimk/UkkTiOcwxkBmfi51kNCpZHerruVx4yARqtKiZUWEfL92m4RHN
fpdLwq15cYR6y2ywTfw6OCa5Fkzxyb+5OZ/WJ3AGJK31uwnf3mTf8Eqs0LfLpe/jbFAHRcUHo3yU
qzDTJu6BehiMMLRLjJL1OtbYhTSpxINWAdepkKFDEhhxwG+uy6Ac6sKcAasvFCGAf14bXGNqzrhI
gkx04rBVFoiZU7F1+K0vxMaKxfDBn2/gxP/psjFaAO1ISM1J74BW6s0LkvfrUDUJ7YDpy/aB8zzS
QIfckVXnUKul7a3IfpkEaqewuY6uuIEo6wSO6u4+apzX/A6RMvLh/vSgRdACxS3zgl8QBDbJAxQ1
5z0WAt+ghfGTXy7WGbeUQVHXh464U/iEEKqa2I+45QCBQqCRe1fBgwNnXTFVuDh7qdSmt9uD/oSj
TirY/9DlqLGIO3esuLMOGAEzMRS60Bebqh130BjIVMzd3/snf2+0lgklnKgDHXioWLluEIaYY9z+
86WK2dJn8euFsr3eDr5sYFETE0IIBwy/Zw1WLsUL+MEdk+Bwzb5ZCHdWwrDv8F8OZz+zzR019Lj3
Ufy6B0f8IGPUDF/UBMUbPrTRsg9xOyy6OJ9VUBpxsYSUfK3kwQruuN1z1QgtGO5V5sb2FMQtNwd+
ZtQTzrSvk3/xgdF5DJHqaYjT3dZELuHIZYEjPkfQRsBdT4be9u8RQEmACEPR0jQOrMBflEv6lA8M
Bw4yrMaA9g47aqGF2r+VNdCS+DEwfuMsj0h59KXNK046U9IQMDeiKUxVM/YHNUrZwIXMycv0HxOu
IeXkEL6kikyZ9pTQfGYK2ep3Ub3tx1GhlfTF5uDiFK4GqbpLI3d1Zv41nsuioET55QFJ2STBHAm8
utDpzKj620YNnKs1gnKB9fnOdsNuiZQUCSzaj43BCVECvMJo+8qF/TYwfH5UrW+p1z7QY/oPyDyI
EXtBHbb6MVUS2HgvG357gx229A1MVNv/I5vM0j5K5MB1buLKmEwEiRohVJNFH0b0zVYvdPT0R4Li
UVApDaTWIXKyU5xkythCQ9MlJ+LNOyxKqO4xks6YMjWO/bbJbQqULE9eA+/YXw81RoauwZ6CwGNn
gOw9lAaGEqtgX1qJWZM3X8pd53u9mM0sU6HVRpyOKzjCCSpm42KirLLrgPHYQ4W+2yw2KjX5CVZp
9WLi0K8crSzUH8Co5E86wwIoMItNMwpPx0HsfJIE7h6XIw5QbOALfOUKX/gxLr4Mlkqf6pSvtQ4B
B1bzh2cX/YzSvNGaanY4kRZno6X+AtcaibZZwXLZEEB36ibqzjQ4dZ+df7xNFtOM/TQop/43biaL
W7feWMar+GyHXbzKcw7UPTDOQL+5EX37JpWsCDOKUuo3q8QRTZwaE6u6D0ZHUUrJLOfMCqGKTmtp
KWWgpq204VER8G6z66siZ9Ps4QnqI5wqw1D8guq/xq3HNJrryI6tk2dbxZ8TcAwkvSqXZcVP8APr
ukJlWfFT10Z31we2xJKdAjgi4Os6xzg3MbPxsXPDAWz/reqEPwJte/HIxqVddzVOCPZqsUbN6wis
YXxDoObH2osOvkTx9qNENuqBfleb8XiupHkVwbhhUzxw9t2mMnnRGKFoZftK+MUR3BOqF6/XJn5H
ELz2j72T9PSVOEct0AddiGsnYVDvw3/sruNzTiflqebrf6PKFLfPTe5VFbVSpUZcRckQeeCfyA8s
DsEh8RD6ZQTUng1Jm7nIVNInjtINZBtReTZjX90+mCyBUQpWx7P4mTlAprgXwO42FTfv/ffs7ghA
pTrJ7wO3zNhbfXSPZxogY/K/shW5uYRfyujlbTinOMGcg5uijpdC38wdLABIrrRCZq+k1LqsBrbY
86pXVXTB6H09oDDXr74mr63NxkgXVX+aMwFFoq6eTAcEaTC3qg0VF+63RycnjNrkxclGiUTzDNi8
oE4FZGmhClELdGLblorVFWE/w2AQrLv+bGTw32iNEhzHNwwVMak7g/3syAZBO6Vv74kDIx/V03T8
5snfBrFzS8uvVVOR41vdF+owGQrg6UE4W6soELy6MGFiUOkMEYdDDejbVTxK0CAiiCmr+ECa1xP/
NoDigTefDRk0gJ7AEepa2umls2GtvbW+s54ANobswDB8vsizSZQmTBe31Bn8qnT0o0UFldOVISbl
tK5wwS2uVx50C3L2jYpEk6c+PJom5b8xoS7gMoyjtsLrWcWwFPGr1GagBluYMYmhqkvRfAayUxz3
ag+BEsreGB+4Hl5lebL+VR+1HYQIvr/f0w7OTgLIN3fxllT5SpdLl9I3PJyMz/qsORoQ2yVzjcRg
ysf6dNO1r4U2lTBacOH5DiWTUdsOPFWIOqIy8C/z0ijkeOOEIYofql4nKRmCINMwuCVUnU9Gi7sL
E71qEOvDEORXxLnZG7UmcwHhw5DNMW69xproT6HfNFYixv7K3DYXZVWgQ8vAd4tnjtFs7whK1Yj7
cfpDOtagFQr84QK2T+uqhYOx5jjSraWMTfMNPHZXURTM9KkrFt7RpYMAZuG9F/ZbLAhlJ9JVcVzA
eZvcmUzEcwF/QopHf9W2qayD3US5Gu0FASr0HRWhQEyEta+P2nZDAKLK9YbTj7V36jviBtjn7fD3
/nCTuHNXjD9v4UPuYK3GutzFwA1FswIlBHOd9lPVcAcLOLjUiCuKsl5Q+IH/rQ1kg2qdnpkQFLMB
vXNFezL/EprGu8Qqd/XoOLsO85iCHOlzEXkQUKoPgg57E26kVZEetHps5jCY3i8KUheGLFqYaOEE
Go2U7vTJx3FZYjxFnIZlGPbO82RIpRZ/i9tRvZhAOjTAOqG37uiEsehDYJR4jMjiUvm2Fb/kLa39
WJRNBImPEWuShdtykhgfW4cBrP7bbuuaKEHrtMOlEHUBzkLyiUD9QoguQjR6O85honEiUoKhSUZm
xvHJ+2l5NCGR6vnNaD44b5K4NnTJcNbq7nBPkYjwNaZX9XQxEYar0MKLEXzJOwaycAcN8hjdzn9h
yl6LcpCHfZg+pBq3uoo05j0YXF9+3eUdEbjb2tPNIZTrmuradfcJ6j47ynt9h8LoR5fsi1NcfO+g
/La8+JWcqUQgfp4eQBzZX+zqvOKoRMsv3NWztad8Y0heVm2EXo6uzIEQEYgYDyEodSaVoKfp5c2u
xegEqYHu8GGcr7Q7r/diyaynYQ0nVJ+8agQPhARyarvaFCwUNVz46bQzcm06WOhXWagn/zAL59QU
+23kGSf+QluBnuk9TkR7s80b3Pi6wlRkMK/i0BhR4JPJvdE4+8muswjGkAiHoRW7L53kBFW3lk0Z
X5D27WQ+np20xxFw73DCBT7vzzfCkFVe7CG/pDQG+baENgS5IWTzTNKgNVh7osz4Fzlb/sQamz24
6qZdr2x+qPxKOWUG1+53Wc6BewtS15oOOgL33085WxkwEA4P//gn9DJzNpNxYjDptEpLIlj2iMHG
qYY193YxFR6xaVNS1Zfdy9K8zVusM3SV6lQktVK3H89YZngNocnRFN7JBey4VUib3peHYxuvEoTq
/QNqDNEAtCoxmEvpOoqO8N6vp60vIgrt61BrwCZQD0b+GnWLheEKc7obBUFklVTXx+IBTJYbHcPG
f2QERd5YWfjPxDjbL8Mg1KyxG96g/IxE6qsrc/49kascInApuz8jy2HMviVnR9j9OIsUvuP4Um6/
opdOy/FEjPvLpcJj28lfPmRQAo6GSzp4GYXARcLKnehA12AvkMtpF5tH3fx+MMJRWfpp10HcDNXj
z1otdEVwF7fCWJnokO7OzYuz0K81OmvBZ5mA+d2It8Zmb+O5J7uSyTiCdza1cSb2v0obu8JYRC5c
hUMS3wrd6U4R7q461AcxPW8uCgqSCdO4aiXOKy5MQcDqaBTwOe69fsl86ws/RbHFEYFrSi2bvwbY
pI7Ey6RbzN5E2Bh+C8S3PjvsO9Ce6A9X3xfcZ1rxzOVJ1E5PHBk7ejKnCh5sLoM/SaQ7k/dhMxRz
xnQjSsJc6sB72UGaC8Rhb7GY/HVmVAYtTmk1gJbvbvA1RIY4suGsVWhIxNJpWDCC+56yj5UK55aP
Fu5zQZoABKmzlgrX+raD/PVD1hohMRlrNNFdfUyDZABdf/wT+K36XUig9qDjHsGWNToOavXsyAyO
BmZX8EgMOa8TKW+oiaaYHfu+J4vH/31W5L4b6wdnpbK0hUZWTH3Ibrc3qU3qW5qrzpRw96DNNCpH
+b4H1lFvGWgY12y288OrB9X0qZeK4Izeu7/UP7rUa/t6PcMGYXMyxkGbUzQI8rEbHHZ9/RK10j2L
IiYMnnyITCzKmbcxE+4kMvsuCjQcyga36jTcpR54oHto02YC8/rhVTw1hLB3loncpjggiJuj6mGg
XrbNZZvCv1G4i7ntcyC5TekLUM6pgzffZS81twwnCAh51DVm7Jjx7L7tF33Rq249jTUWNaik+peh
EGwiVEYb1swBcPjtwKOHT00n9XHqDCjmEHI7wh8z9W5nYx98qkdbmBlTxVNs8zTZJL6cy3rrEugo
gTwvnXT5hwRkjHEjeib60mdfj04Db5TuD4nWoGlAc/17UtiWwfRieUnhdaEmISEjfmXYrbDi5LHv
azG4yX4uvgmI3P/2B1E8prgZkFbrXKhk1zd/2f9HW4IJvsUcFpGIKtWu5VDmkNgJ1lslG84hUHvu
4wByRSxOtgIHQaqhyKBkFpulIxNhypkrZX7IAvBqXvQevXEFsYjl8TahWb66A+dKaj55cSVV4yXk
hPjN3q8P9T2LZEK4yKzl3vUmXDrnRQmn76Qz6tf8NdYI4CTAJn9462n0uxF7tugJdN4f0xIiTnzf
FrwbIYHNIU69+MWo8FKoDNruPjD1eU2T6ohC2Zk85tF3UZykzRzIZHRI7EQMrws5fRSzvupwusbW
lO2fddYO6SeFGkSmGaEIKNFw8W30F7vRWWKTy4JVlmgrBMLbethRHh5PkE57r3VQDrtOT1B+FTqp
VQiWpABC89NeWBVwno66OLuTCgdq28jI/FVWyAREu9SKvwhtN73NtjNLqrekdXxcoIZCpl0YE7qR
UpRCMR5yHk7MYYzJDuEDqWFK3zkBLM87WJjfH1xrHlD8vRFEYmHdAn9RSajFjYH0VxhJ9l+EL+ou
ycGQXQ5fwhVwTqxufaiy2MtO48vSMeuhrjhBwK3OZOXVeOzl8pHo9rDYUc+PzQOSOXC5Ghxpc3uy
+I7hpeM/gOVMD3R9M/oWooA7tqmAKW//qnFJ/D17YhpGDkLffCOmfU1aAhsatSWq3Vcp/2Lm5VBA
2WMr8X081rwfcSvlejb0NSuNwW9otnUK9iIc4uq4EBxbgDDJqHXrKDBOsSeIb3/HLnlcKwOAEBcY
A9xxUn0qJFL+xdsQvCjAQUAoyKZE48XnCHLXvWaIUumNWk1pv6K2McsMjoKVJKAW3AnclHoMPvHG
H0/GHcdouZiQWXlIomuvjUq7Hq6Rw6RjOUhmmTspA344URNldr3MoNquz4LIRGD20pKa6DtvSQ4G
kYshBkySwaOFpOxun/AOLbC+WZ+4nYnLSEtArMDhbq6gWgoFucnBrtU+WnHa5eyem4ET3SG60jo0
GNmCjCcvPEL4rpat9l890RQVM80o2UkikBQH4ZC0E9cPpF2gz46HPdWoEOJoWKTMZ6i0TWvQmKJY
f48ZnpKoc35r7Qd2R8iXjV1jVPxU8sjqGuNoLydlatx5kk+opVMMqLKxfxdNKdOV5ZF58OSeZteQ
7tpL2IlYszp4IPlQdgFvicIlZ5KSLCPme/H8tBY5V4q8QnmHb8IFQpZ6g5RQgxxI216LTjqaRGdy
onNMJrPMLBSSY59hGtxdd+fnzFtvZmB3+ZeDZtSuMHK2b05Mif8U75PVM6OZqMl3fCCdUDc0h26X
EqFazO7bw9ZWlSQQCW7T/7/j07xX6jEl4vPt9OkRge95NN52lK0k4zh2C8K06UYdBV5J1zs0t1gP
KCktHqwCSNpuCLEdEgHQsrt7DeW87C7FSeBWyB5Y1O8FdJT86sEBKmoGigUwVfrKbrLuplj60lS6
gQ4LTEKpKwhZjTvyeJp2QhedMT/kkn8l/cHVIVxQnfyHAURYSCsyOvmybs/J5Fw9mBSJkIiM6C33
MJCiqtNxDS2ufpBusvwhk9lN36ZRxsoZ113MiljmGnZnGFlRdO3yFysJZ1HeVtgQJ8LBva8XD02P
ycuU07qTClnTH15fN7p19DTwJbZkY3r8IkhJl5OCbSuQojt7BS5ytFyX3J/N677KTwVRD3Neb7EP
LfJwiN3kZTtOZXIvNPQmgt0tUiDZKgj51e2ElB7nORXd0s72CtLbSPiarg81oJ7HO1MMsKkxuQI/
X8ZtWi2QBAxVWRilEo2VHwXkjxh8JTqEYbFUDUc4ZlpfgduoGQ5/QJnCX7QfbaDn0RXHEqXjSLK6
MXgv0xk9msPdDeKpCKYykO1QXXtOEgSL+iOKDweZ1HfNH4KN8j7vBY4Pmif0DeuQrlSVgGFfzZzT
veIco3+KmriADIepB3EUOebCFN4toUNsd9faCIwt8YJ0y6Ay/pYqyV9h7kJAFKVH8a1uVWxTzTpo
ivMHkdQPWC2XDnFCW3kFVFunD7DqhXc7NEuayp5gW5AjFWnLd6rwhQdTp0Sd11+3tRsIAON5RbAF
cWLGkMltlA9j0M3N3iYT7EaD+lX48vuub1dWjHZhu+vruU7p9YaLLM4CSPSYSv3pJ5TTndFNsoQW
/Y5zy8cA7UD7kyohi1VubVqyXllqeThiQdaC9/iitHvcLQef7Ii2GfeEXGLpqxlcLNMQUYMH44Oz
HLxBboREg6q44M6wgOx6UVdfKNL7Zxxq1/VG2Mpqdhkxw8hOlTMf0YfN/HmnVDEe8EeM95IU1Amk
QzZP0GiioQhKeY+vlpJxXb3XB6/e1o2cJR1Y9easIRSDVe5tCMWY2T8QcYCriVfwwzBjBllrUjWa
LRFBvQqXg+h96ootfxJiQ37OhEV4WUatQ9tlpnMqqB6b19/wAkLHmxtVi/JYaaEi8ITAlle9Nagq
P5ZEFG454eSnIYI7cLCcgY2x2BPVnxsKDkUPVkSgJFFMn8e0wOy2E5kGxrweHn4VhfbMbvFlBhPv
hqTi39p0b2ZRJGl8UeHY4mFvtvQFNfsdVIhGIHZG2gWIhiuuve5xMPX56pdeXsTlM62cUBT8KfbY
xKrJYPCmpl0IT8MUuWDI6NcWMXGIXXGvtu7/gZQ3IcKapZ/YKzZ4MB97bpcmYgaUkbGKH0d1124P
A8a7nkC7ZTza6FTUc4XIc6E9aqGv+c/t4Lg7BKFcWr1abgeqyn9JTK2b9/23noEOSNVnAmL+Ewxr
6a0I1RzvVmkekIeaECq08ow98aTSUsuNy8nHg4yMKeciuXl9c2a9rLCNhK4RPzqX72g5856URWq4
rVwUGw9Kcb0RJoK6zBHDedmsjVXliuepYO7nHAy0LB5blUdGu8FLT3A8nW/r8w5Tb/Yo5sHOqDnL
Fr9XKna4ZevTx/qaQwdIUJlB9bMmEZ5X9U6lvyuoNaz0bjuoD+9Vzp5y4RXawnz7Uhnt+PMVXYmW
+pazX/hE6NCL1JTqAUllHfegjupf4qoCE9L2buq5rymb7O1O/9zz68LZCsj4E8BFQvFXSv9sC0A6
JXE2zU8+tNdPvnjF90iH28tFqmD/ly0xJ2XPdaSbcBcx0Q/3DGl5SQMMq4T8cKE+t9A/Mm/g0uAZ
o/P3WWpjfGlGgN6qmvc3NOSVRMsK7k1DFiNfrdMSxbFfm6sUoaaMw00nkrB+yf/b6qkJyg2zkwIY
RMnW4FHOHec7iTItfBiI2Ta23ekYUBAGfLJuwMHBqGnBJiNA22P5cRbs10GoR1S/IGvYCuViCXGv
dWVbXI+RFis0ZdYooiPh2IZL4AptOSqGHEDWAN7irQrKn1zE9jlKQetFFIZU0GsWFmROPxJADzlx
wXt3kD0gchNhdbjvqzQoB4qVEI/PxWW7iFym9kn9qzPPZOJJZY4kZ857xFQ8OwqA9Q/N8yXFagTw
EYvnziJdIoslUg/W/me+g28pgIkDGOnox5MilAwR6igr9D6mzEiTLyssIriCnbU4ZlYehKjckOWB
oTGU/VCFZPvfJwKBzaMBxgngQPxQlE9BWEV7NlIdL4thVEY/drR+PnVZU4QkUgBv0pmuDGmmUZV+
vogHd0JFf9GO61O30hHNhy6mHjVHRnNmf01/TaGKh/+nvcrkiP2k+XD7UolO8E6GaXMA/yMxAa/j
4c8L3kAmJZgLATPqw6UDYKiluH8RpPurnw5UdOwSJ0TEMXnULtFv+iiP8OGJKu2VthC3WLNHJIcx
huaVeBfdDONqC/r5grlaSliqn0Rdj08AnoCQJAfbWg0y9FuneuW3BWnIt3hf/RlGDAod1CqBR64L
mxhC66c7Cq2ifs5Tert6V0T0JzK9iabf71lo6daNVHaVp0Sn5u1k318O3kc+cVAUh8f65L7vECnr
cdHwp6d8yau6bS4upfRUAaIfGXAzha/lvQMH5V4QWVwCMuga5KsqeSRMkCjqqcmnIJ2Y1TUa3OMt
7aXAJXdkyCxY7h8/ZXJimgCfswJ7SD9Mb5rpwDg0y2kDLL0xENMTrnk+M/JKt2RLR9dLRk7r3Od9
l+y+oPChu+guiMJlFR629hJ8iz53DPvHuSN1/MjMO0FiXE5XPPRehtfYIPf+rdUMk2EjtDcA0jgq
6V/cA8PKz6Fm3MKWFJz84WONJns74LBEUnVAvHD0zsbKHah/N7WhhzhlVVzpspzDvO2AddwO06tN
zTB6pL/5SspaXNQLVODh2ismKSJ6XJpkiPy0dDiY+o0ZP4bDsU6ukpY9ngQif9E8eWpsLyO8IHnw
QAygOgmgY8vqowDOPTE3NViBPT0OwQa7RBF55FSknAKl+MhdzzmSlYnGEqMNj88MnV8HR/fjIknd
Arl85wKBh4HQXS4ReOgu6dThOi8SR33bzKIMXEXsd3CcCb1qEZvnR5vhwRTyKXnK1PnFbtNd/ShS
ihL7vn3uI/H2QSIdPal/yRxyhjfOIMhTdOR8rYOjTOtvwOzY9IIo64Zbr1yUH3hEYyAaZoPxMmLP
ZqoexZNgeyrShZbC7YSmCVwMwo9us9v9/qFAGbs7QzaufLkFgk4iIyI3dFXBbHULO7UGu8BQvp6a
39zmTQTK8NCUguj5lI4rzqZEx9klOXjC5u4SGI+FO0Ll00k5geZGSG9LgEaHf1EKdLGUDnNldRnk
OTAvAM8CGVNm/60Vpr0ovexk7gFFy5AmKyt8byfxxrXh/iCyRGu/zVGCACM6ReYKjRgmz3VsOTZl
g56J9h5p/iYrFFSzWknTUkr7Kk6nv3rDe/oHtLoAVC17P2tzoc90z/JO0bMWSlSPheEw/PpoM9wf
LzzbbrXcMrzq+NujaKH1b4Ze5Qnoexiyg1AXZwfd4mDp6EHoPIrsSYOUSmNM26i6zGqcr7s3ZALg
ESBOGxwWzvunrTCa4il9AdOCMk8351bI+azjC3Qht9OTBkHFj18v4/M1vEb3tAQefOyAflz+rs0n
DLXizR+Ra/8bPM/SZNmbpiXNedNFSr03e5CrurhApsJyzEC9OkEFIemtvnqXiuG/wwBSdn+T4Fm8
nj4/hyk4vdusBgx1QOTdJ7GjoSK/+fLft/oMa+b0wgMzkJ4KaleTJi89zjCno5AXSrDkRuGsvCkT
uJq4C2uAcaZH5xisfDXALYbGURFqEwe9K+uLxsUbsIWkbRdmvovE7yZmFW8lG3pJZHjEaMHh9D3/
0zCFefZu5mp0ZOiQQywuRwcZGTfOtA5KFDUXjF8km8zUb5DVXnZgkzSjd/upzGBeAYAITnbzRARL
kpOr5YkZY87OzheEG1D8RaRHiXxVjhY+6RGgqAvJGkYVrZGB13io848952WoaexUypctfGVA4flM
rpwPiIUBPmqTxvlmO3qvncU382rAUFp6VEVWXrxGgu2a/R84oVWzzfTHpBf5Y3hYWDZa0IBEC5gp
RaKW9NNxofhVv5rK1VXSsO7/Hc30faDa8yh2G7M0Tjyd5SabCneo7F2dldoCBRxsjY/admplHpON
3VJObY2umyGI6wN28dY9515vuq094qdoCBa52G3r4Kk9d41kSf4aN+GasZFkY0hOSU8pON9UdgqG
e3pwDtBnfBQgiA0XEaFCwO17yjkajjoItk7JaPQNUfOt7vnojTSubEhujCd7XG2uMX5MtSR3dPk/
zNRihbWTM45749D1mAn3SFJNF76piBxh48suTTT5nuS5fCHyqUuBb0t16DVUHo4XNDBD4TK7PlF1
w8BPsyreg6gkvLb5Gu7O8M4YGQ/QY2zHoekujJtrOWMJxyiDVna7tl+rIj/9EV2J+pibGTnb1SH9
mesAbm3xwxckuE5kmEW8KP/koK2DXQum0IL5W8owsf5l+IlNmmaIkXe8RVKUHmnCEE58hZ2JTZT6
gRAmbwwJDOs4/4/ig/BrLUgVOrFuULBqWYeIobYSlXfuwxhXqyjh0Oi7Irhy2qw8Y5CAdVs2vcE2
JpRKGvd/p0JIsLjMukr3fNRh03y8svRD+TxVES641mEPdQicGpV6t3MqL7PVsvPrnrbWJ5aT8Ik1
DFCMk7U5OcjEnKmZjsx42qzZQ83ZU4W7vWhAY06xapDezmEVNoJ1Pr302X08HQQkA60Yt/ADp9dZ
UXPmLU19doGd4W6MwlX92zx43i3m/cyg4Nr/6TFHt+tXWxE0rEHUW9CNBYckZ/Uy5cj87tr15Qr3
xt7LrFCU277HT1680r3Eh5HqrtVZqTuGCCmeye4eQLr6fQA9b+/p4s4SV1AjE0y5IqLmzQBtpj9G
6325FuTpycxttKUU7CVV6qUID+j4/zUZ7QC0u+7uPpvTrMWhFFZQpqSQhkRqFSRvhB7wfWevINjY
iRlFtsmqj+2nk2m1E2bRHeK4QjIEo4e9YO3Zjg4FXS9qh2sISuNXt1UDVZvW7n1DtmdHfjfKlM1t
4ZxOFtxaBKHYTrhKAllbQnyvPhySqIleqetFHpSRcJL5QtES1d0K0lTkUtAnDvly7qv7ru6ILwRW
VnTy8DvAFONBSj+zYmLonlIsNTTRANNAXmjG0bVwMbKSkyWW2yM8ecUIxx2nU+2MAfcg8ZEg17a/
NGzPP8Uol12iwaLqAc2nBanuz/8AZ0e/2VAWiVPdpSUJ/I6sy81OIgiF/W5u9OD5R39sksICF6mL
1VY9/ugRY4b4JWGUxeMslDbWKaJ+kGdOPQVBwS0Dgv4p+MymwwEI6lZO4qnFEGrNsbK17FLHPrra
Reyf4grkEc0YPrsj9v+iWkwhOmx77Vlk1lYBk9+OJFYpPIIr/irGliQRfYS21/1XEjIAKHuxBgDa
8hD4WuGsUXYWSptLiiHEFQbxTP9TkJwroL/wYSmlopE2gUwrLNcaEkBVe8U+hFtJFGneUmtBtcS3
uNQxNZY9D6qC4SI6qNjjdeafC1KxgNU7dbWSYt27L3Uv9AFZnqmGf8Iy6Jo9FPPsb/8PZr4kLT+k
7BEuI1a92tVc5edVNBO4rPLTa0rDfn2W6m0yPZo476OHTDEckMcz2NV8ez5KuMfNqT3P65azWi27
cD0oQCt7SsYCatUGXQHNl5gCaaatx8azT27N8rLw7QLOUav4gLltEFIO2Dhq0EmskSo9ALAp/pJF
mIOcPirCkScnW0bAZtkN4C00WOaiiar9hhvpRAy+fUuNYdBE6AtSeGwULsc2jve0ZEw/OTLCaklM
0rkRP6OY5zT+vCVv8jxyJnzcCSdkBcmPIT/itzKv1RQWBDPSbdhaAdmXIXN7HO/MUq4iuOrq10SD
rq4rihrjbwcneTCe2izA5MgMRRS5MyxqX4qk/EacHnwYlOW2Jmn9jMQFPNjgK5mfALLajskfRNhb
+5RgiwXEO0muU5DzJ9vLjF1zSjOIT4HEf963YlIOCcBuF3rCPMMjKlEYFE5KE46eSr7NCHQ5BlY4
Kl7vG6Jxe5L5DO/F8hae095AwtbmTnnv6B95ii5VTbnj9m167chGtlcREW0+zJvTyMOoUcHJZPVD
GdaLIpyBt8lFhxcpTlQCxGIP9S0pJkODM0snyB7cRZeNOowB29MGD61j075o0YXZcQ3KzC1X7xEt
vqeDxL9sZkEe4hquwsHny2oeYc4apnB/uABO/WBU84j5YaRUSywtN4iPIBazkb1y8wb1Dpq+WJUY
FRzvvZVfOJbp/rhwX02+hVIrAMFrkASbAG+ZRpw3u+Xi7GnRIIPSCWkpkLQ/IFftX333PjAWctaW
BC3Wlq7srdYoJvWs6+mAHWQblRF+5sgc8TkDBZ+G0L3DGWN+/DU6NrkeYabZbxw8ITkkOfq16cyS
j2W9O5nBkYJnn3hGjTLfB/Snx798GkYOB8ZnDLqj9d/Alt6pzEUQlCIqKzEr1mGI/K57hGPPO0wy
sbeyhfJf/mp5EKpQCXsCiPyMYrnj3aGGPL4zAhO72cQbq8hb0e4RHQsYnSwLkwvQ071AOTtx2yE1
vOKTBfHNjToGdtgLYQNlQpn28D9NotE6rucRJpaRHycDijOJ+KYceF5DmYKjydr3RBM/ghCS/sKn
p28YP3RpjFWw4SDR8wdeKnRhSdaGzLbs11KUEUTXi4uAKfPqL3WBvBZ1Gg9aKNV2TxHzE/6kj8Yw
uBKtrE2sK4Wr24siZNSuG7ernL/V5fgr1WCNIjH7oAbIJxKQt/5LeVp492J3nTcO62lTpfxvPcgC
0e8R/kqIIBo0yWYmVzRYtguvIliKvePSUhTHlELY9HXz0w3VkQ9gsXb6+ZEOWoOpQj8swGpj76p0
cwlNsSxUjpGWMWBb9NRbsP8o/QDNgnNEAbqfRPJ9oyqZcdncE9hKInnuzh7bDVFZV15Wf13dMs/v
16EWKiRk9fGfuSKm/xVFAZOTm/OBrBJ1yydiSOcGQmQSi2dQ3/Tr7lBGKaFVn6wQgbibxic67Gd3
D/jf00/fQoGkZ36nXTYa/VhIWPVimfT/TIV7y+PMjf/yaJh71RyBXqXr7yUJlbw7mL9GOYY1gTA9
daoIwfwlPhHFwkt4CT2yHvr3v2B8HLqKKbjYy/k4GNBYCRoJfa9L/DiElnN2cTJbkAu5XMGPnPZn
2WzCxVM1ePhYPeoDy+TmY+UYgwaAis62QVVb0Lv84nkZLNV7mbTRg1+wvsQOFwn8G5Fih/pIoh8s
qo09n9pSBKkcpUe3mWAknGVZYP9UHwZN/Gp/8m/4AiajPbaqo3MIiY9UM149y5hds+HjVS32W7br
jl4LRNr5vPYJ6y5uCvx6OUHKt1KkkhBngup8C7MS4iGGzoptEeHpsiBC6H89aqnmaS/sP4XrlbuU
oG2fJLbD9F7FCVVcTktqVwH7avT7Ngh6dweiSrra2UsxSV+a5e091RGVF8aidwBB9sXK0qduT9Tz
Vf7lPItVCqnHVHFsRJRtVKuJEsKm/FyDnkEjbuaRAgAr4GXM3VBYmfIBlKLwn0+xLgpQsYKr0iKH
TE/f+58krJElrK5GOEjnG7Pg0w8Td7LQZnenzqcOC6x0bF7N4ZZYNzW7LZShZyyky/yj+je10/OL
po3+i7LY8zAJcd0hVzGN9GrVDca4gQM10XWnXBDkZ7eCQpd4AetXUMqTcs+9tqMWEHravPhdFJnk
c4vbGxNoZZh4hk+JMqsmaQPAxzK05nyCpQ4pLLCdGD9ANYU4UAvu20Ej3Tj2E+jnhZ8GcyvOuOZK
Sl/Lm6WtI8+d8hWMtuxmG6nC8vX9YPqGB5zgAtV7odvoQdihEIMbjaNdaqNh/z0dnti87LQkPoCp
q+moZpFDOydvyHCM10B6TmPTtDWlI6Ll++p6YjnFjDKyFrr+ot4PoBd6SO77U9WLQtQo31zz+THT
/PyjwgqnsNFEwWNvUrSrxOUnGJboQmhfUMMJ5B6Scgb0iVspXvEDVbwLEFUppv9Qe+AfeeSd8YvO
nmkwllEFJ/KLeKGndBkeWvf5QdLqq10/0MTyJXbUxMDgsdFfIEqd+BE4Mkjx35mxh6OiOaPVuliU
kWAxH/qEH+Dgl/x2CaKFz7+cuGNTADrBEdAyJRrkg28YjGq1w79lNu7jjfjKkXZjm7EouapQAq53
6uMtiAzsALFqBuRYmuK7ukh3rduhfI4ZCUEIbf2M26xYKBnV9qiCDkJQNDaK2GmTUyRS0++8cYsg
pP3amtiEZu90D4tJyAZQNKolzzNEKulDjnGjaieDbrISIBRZYiTJSC2iFp0DRd3Zffb/IYFPUp6I
E5XbsBc1bH7nylELySSGGoXo2yQus2VuJitRuC030QbwM8szO8Ww/KwCzIOMRamZWJFx1/AqYMR8
a/4Alb/H7uP9RS9S2kwlBfv9HTUP34dXCbLyeGhnXeGRHpAw/JnUVw6NbKf1EbTVWjO2V1lFb7RU
da6CAhaExyzyZmygXmbhN61pWzJSX3uaoxKQTT2jBybdtzlCbmhM5vpD0Q3JjEvaLYeVgHVvOVVj
NytKsZAGbZ1uUtZiEZi9vKLT24M8HTOQ0P+5J6/bNmhXT+ER41Ngx0zNV0v2skKDutieBB1h7r8p
tm9JHJSvjJoWa7Uqsumw0ynAAVZ2NRXKbwfNmZuMkPOxt9EJT+oWqLjxPgaojea68fKK18CVYwZs
Is2NdOo5DIywiwE+x/2chLnLGgi6ainuG2XNwFYQfMaI2KmPzvZkjtcJgjXb+SI+x1ltmgM90kEN
xDmAcLswKTpzLimB3H+sbxg55Z8lTyj39bEyZ6JJGKhmRuGKuKnvD7iF214W1o6fhlx3zspkSyKL
zN5+K3eVpv0a6X7iFu+cm+xmZ9E0t13K6wbW0TD4DnQum6oJT0PO9xSp6Gslx9WBpR1Mva+eCQNJ
/aFmrw==
`protect end_protected
