/*
 * Copyright 2013, Homer Hsing <homer.hsing@gmail.com>
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 * http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

/* "is_last" == 0 means byte number is 8, no matter what value "byte_num" is. */
/* if "in_ready" == 0, then "is_last" should be 0. */
/* the user switch to next "in" only if "ack" == 1. */

`define low_pos(w,b)    ((w)*64 + (b)*8)
`define low_pos2(w,b)   `low_pos(w,7-b)
`define high_pos(w,b)   (`low_pos(w,b) + 7)
`define high_pos2(w,b)  (`low_pos2(w,b) + 7)

module keccak #(
  parameter r       = 576,  // bitrate
  parameter c       = 1024, // capacity
  parameter d       = 512   // output length
) (clk, reset, in, in_ready, is_last, byte_num, buffer_full, out, out_ready);
  input                 clk, reset;
  input       [63:0]    in;
  input                 in_ready, is_last;
  input       [2:0]     byte_num;
  output                buffer_full;        /* to "user" module */
  output      [d-1:0]   out;
  output reg            out_ready;

  reg                   state;              /* state == 0: user will send more input data
                                             * state == 1: user will not send any data */
  wire        [r-1:0]   padder_out,
                        padder_out_1;       /* before reorder byte */
  wire                  padder_out_ready;
  wire                  f_ack;
  wire        [1599:0]  f_out;
  wire                  f_out_ready;
  wire        [d-1:0]   out1;               /* before reorder byte */
  reg         [10:0]    i;                  /* gen "out_ready" */
  
  genvar w, b;

  localparam OUTPUT_W = (d == 'd256) ? 4  : 8;  // padder output
  localparam PADDER_W = (d == 'd256) ? 17 : 9;  // padder output

  assign out1 = f_out[1599 -: d];

  always @ (posedge clk)
    if (reset)
      i <= 0;
    else
      i <= {i[9:0], state & f_ack};

  always @ (posedge clk)
    if (reset)
      state <= 0;
    else if (is_last)
      state <= 1;

  /* reorder byte ~ ~ */
  generate
    for(w=0; w<OUTPUT_W; w=w+1)
      begin : L0
        for(b=0; b<8; b=b+1)
          begin : L1
            assign out[`high_pos(w,b):`low_pos(w,b)] = out1[`high_pos2(w,b):`low_pos2(w,b)];
          end
      end
  endgenerate

  generate
    for(w=0; w<PADDER_W; w=w+1)
      begin : L2
        for(b=0; b<8; b=b+1)
          begin : L3
            assign padder_out[`high_pos(w,b):`low_pos(w,b)] = padder_out_1[`high_pos2(w,b):`low_pos2(w,b)];
          end
      end
  endgenerate

  always @ (posedge clk)
    if (reset)
      out_ready <= 0;
    else if (i[10])
      out_ready <= 1;

  padder #(.r(r), .c(c), .BUF_SZ(r/64)) /* BUF_SZ : words in message */
    padder_ (clk, reset, in, in_ready, is_last, byte_num, buffer_full, padder_out_1, padder_out_ready, f_ack);

  f_permutation #(.r(r), .c(c))
    f_permutation_ (clk, reset, padder_out, padder_out_ready, f_ack, f_out, f_out_ready);
endmodule

`undef low_pos
`undef low_pos2
`undef high_pos
`undef high_pos2
