`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
mDIOS8PXcK1kR53SwDDegCaYI252Xt/PIM9qOoHzBCBlvrVEgTfwXdYnFtcyEPAXpOFIMhuhuTg3
sjA9gZ9Vcw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kT/jNmiLcCvOm4mpYCI4eygVhjFrnC5AMm4j4uszeOK71Xgl/qVCrYxLPF4aDiq6Aw38Zd3EDkhF
WeY/0jcivGAjCONQZaHxaNOSv4VD4dsaZEspChn3rUxSKY8CAeCj57qCGOUg/jx/iZXNPzgXXAiw
EdFDmWu3pYcOmd5hOhA=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
rJH2B3YYUuS8PnW6+HTozZ7g9Msv4UCDaK7jjFTdMhbEVUe1n1O3cYT0d94U8bJ/e8qgYiXca3GL
5BzZ5xAcnGzGdiRH4RCfIrrnkEJ+vyo6aJftc0LlV130qCl2WsHqeh7pvyy8tMhy+P4KhhI35zY8
2GgrLu4ViZiS7U8ifybQfI0WVFp23O+tFqZXf0UcisnL6f3G+Q0/XadW3Wj7a+D5yf+J6OuU8E0Y
OInAHRgJFR4mFZ0tkQY0NveQsYlIUEubV+zKv/35VjXOhTmNX3afzW/Z8Tf40vOkCE5MLNezo+37
xsC6cWHbe5pE8L3QQQwddl5SR3NSw39JJXdcNg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XKLsO8R2L+p21gFpfS6RqZ/S+qwQZEYn7ET4lzv7ALj22WZjLj+T6sPGqeSo7jeqNmxGnae6P4CR
cLwbIbr1tyZRiz4SHfoXOoOR1aty4sliBFq0Gx+Xs8idPzzJrG79VClbilR4zmW0btnB2k8nMnjX
TxuoS6NKvxzNVz3oyQzntXhobenf0t+ximg9LIAfhbtgf1IR/EUVHUcl0i0TtXRVTdAQAMJO0N6h
NSu8KAMg0q0yIPD61otHRMUsDIQIoBmQkoOxWa4pKUy41SO2RAKYDHEC7t3OAoSvi8kGJtEyxxRq
41HPKlN1NcTyh3+ghtXW+46UZSbOauWYV9/FUw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YBSdxLYu8i7Kfsn7jaZ0PXbcgVeMZ11qZ/BxILsQQ2rKc9jSxY2S4+7MC9GY/Bn20R9RXBpqQ5zS
NQQHA8UaJJbD8e5Se1k8ajJSHJORcrESnmeVvX+vRd0R02OV4TLOlQkqgg+wbQnFucszdCeYXGrw
MRZ/9fFI4bW8r19V/32eFIsxHm9J7+asY9fb3gk3V5y7zbKR7OiczF5ObPdO67evw8RRO8bxy1PK
SfRhfq2Lzchy3J8BTMeJ41PGhA/CqGO8aJ5PPQjACln6YEAcEvaKGfisSc1hSwHmMLuz7SUCQo8H
DqXqF1Orp2OqPummRTbSja6a84gVBxFIrjLbhg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Iv6aKH1p+Zl+lBu2Jm9rauXPIgtYGRzAItQkUm4ImgGxvI96zhFJ1u+Fs2Qd5a7bWLqXL7gpjEmh
ecEPwGXx8SCe/5HvJ1JuD7W4LNSw6SKxzYVFIjaMajuVZkfi/QXZEHwyL1Vu2I6eReWlK4tzpWWw
9Vom1a2LQuS3niLiEMM=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
KUKtpJlLjwg/TkSq/EVPQ3IHPY7bbmJUxOefnagc1ktTJZybwntUvupr9vmVg7KIwX41BupXsbLo
xT7CeSLx14bXAptml5AoDeAW3bXY1Vf7YMUyTtck9Pq769VUDFRLs+VsewBxZQm+a2LHlB0UPrVn
puZbhOqa3/KisEAv4IaljomjCrOr0N793QaLWKnL6b+pvYemk9SW4fYAFNDmEH4ZctSsVu3CgYyt
OArlPhNFvvaIi0mSCV2s73hHff9eONeqUxR1OKvFZPtbsj5TaKbHKqaDSVwnHffj5qUrmNVBT9MK
PA7eNEddw1lMA9StJu2sDqVdD07cietzt90Jqw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 133280)
`protect data_block
BOiq+9cM2w2lAKzhhrczNsl7bNcWJi842xHAalNrK3bm8vW66MR0911aRKdJZCU4FfGJf78H8hhT
fGRPETDZfSiSyDnSCe21ebwr+0MFHWvPKir+HPc1j4kpiiuytbk3FIKodu7+G02dLTMoLow5cbYP
qen9ud2iJ8YB/AIbHLrxczYUd+xoyeAGN1qg/1V7q3mfAfQRRw7b43e8glFvn0L3a/pmfb1120ki
+k0e89ONfZAiPZlNZrU4agMctXHY2/aftQfOlH7vslwzYYC9+AIq7fZFElqJIf+QDOnhIT9mxSfU
C9uPLbjpAju3j8zLVI6J4u+bTg955PVTLYhNHn6iplXKPtQyLgf/GDJQyC/EvRsxh0qSq4X5BQQX
kzqhR4NKrYDbe90D2GzYEM/zECgTNfY+SBSsE8uKQt/YZPOx3FRcOExWtti1l0SYEVln00I1fO0O
7+bTCpR7d1blsvnSbbkWqXTzC/418pnmXSQukycsUygqJqQy5Bj0PVau0qMs0hHFU4GwNo2+C/Xw
Cly3+VHzBnWE+a5b/j+2CahTHWJdPpWUl0V8SfQocCe2d3kaYYp/dmk/AgZRzxmYS6nCOb0jlZjf
LAMSm4MK832E2ONnhDFgL1lgg5FVUcj/JAUGX+ms5CRn3OGQl4AtmwZTMa2h5A/oyMZcrOot3lqf
tyRk5bWmLyDicwzDBtOp0VKjMJ7felFH/UE82dJKoKJwMlIO/ES0/DQkRzC6zVeHhQAPS+sf4AFf
wU6/pVLwZxgY8hE8ps2wagERvSy9yHppsU3tWqMsYdGUiJsBzpbLu1vlXaDKL1wANqW3RwMrXyNH
nyJyBqpt9/fM6o/6iLjh70KjgeBShpdSKrbJkmw+zj0F+azVYxG1QHAJP6zUhBHEnqdkThgaNkVG
S1jMkJA3YNJTWmTZZW3jK7m5SRRrgEBBgfeXdFzAO97Tt8OU+S69cnjCqKTHoElvySq9O2PEXVsO
13fS32Hvc5mlyRyEJTPtrrqElTiJ6Oyeg/yy9NDdYUMrclN4DtVHYlba2nffZn9JOqXUekDLyxCl
Pufl0Hhj6yS4FP7Sp3+KM1xolbT9q36gx5Dmvy+w+8hHr+k/ytc1WpqrB4mPvHO23xSeGmJTX0As
XxNNhi9k7SWQQH+T2wn4sPNGusGS2RUwcOG+rYui6k0pDJJ9XZ+OFIS/crkjM0nDltpUMZM0gOs9
L44cxObchvH4vb+85Nw2Mulz25jtxPZDJHkuy2DM4CCIJZ6bbKrgFqhxN68viV2SLWcWP1hBdk13
CgoZmC0Tiu8wvpGeutxqJnucwtjdG+S9IMIkVhd+j4gC5vYUewZTphWZCi6Mh52kQgcYppmH37Gj
iibP4y9dycaVQK0C7EemarBSVR3wwE+OPJQSE1mcwnIJfFONNKespUWF4UbvQ9Aw58uafTPeWdgi
yfF85/Cer3vAmx9Q98wrRtAFlS660rLLRmkysSrrvN2riHyiQzcWU9moTaGOVVjGhydSDKT1+c2y
D0tvfH5RVHNsBjGUOVQ1REWHvgkS0J8kxp3dYCGz8V9JdYyLKt8Q3NbrEv6IrF9T6ncoDqTtMHJy
3qMiRvbJb1VHgplOBDiXkeTPZlThL5Zdp5z+aryP5CYyg5SPpRYdFBAtWL7vtX6Yziwya/MB3ouP
YSyI3h6/zV/VQtu4XDL0SmifDaL1SYIMAPdEjl3z1GDlHTatMWNlHjt35RZkgXVZI8OGaE8c4OAT
FoHD17uirYK41cM/+b4GQ75eVL0AI2hY606ZIaUcjZGn/FSJqTkSPKZGamI/OurMW1dV2N6h/dUs
tGRav8XQ7ye6gMya/wQrUYwyZc79AGu5UPZH//Vj0lvoIK508B4To6ebLPAkVXl8+XvfG8lhyT6B
y9cd+p1lqW/IAcBCc1UvR78wT5VkVMiDfHzCyKphONWQdm6miodjTZmYkx6Digwr3dKmQ03MuIGc
YYDJZ5lDpXX/FYu0qvV9cp6oz2sBzNQb3s+GPqX5AbRdQGFtaNhBEYc3OeGJlMSAHsteNLia0GPI
O8hT8gdBHhNrmvSMP8xHfRReZy/Z1VukcuaGE/G/jVwQia4obwWvVarjpde/6vvEtjTxfVMC5kj/
88JUMi0R69AYrD8cO5AN5WuNtzQdjgcdeCcnFjUN+bDGloqHFRSR0toYdDy0Tni9YTxrcHkHbIV4
R2z1fq+adnjqIKy2x6mP1Tv+MFyhlwyqvctvCLWZg01xz4/hKaU+XxZjDRdCggA6Giq2W3c6Rf0R
G+i9HLqdOS5UzdqiFfZdUXE0DAkQl/gpNSAIb1FrOpN8LYJUe4oHV588EiF0HmTcVrkrzozt+yBq
/Hh3nu6FjiX+Prf1/DDItI9ytNt5RS4zfFGkx63oLCuGe8jsH/W4keVpEH+f7iMd1AB15Jgcv1iI
zod3M2Zl4IbWkWSJhXqS0qwYB86pqRN4uMCdTIrARfgyMICGO72KlGATRSDYOA23KBxwQWX5Zd6l
M5wO+JMvXNfXMxS4ddzP9ZUky5eb0tWhSTCLLHZ/9gr5aTWb7G8rk2jIUMWGjrLgO3h1nhVqfHB7
MQo8cDuFtkFXvGThMqVvFw6EaRof91+7uL2l65lNXG8/8BQQmR34gpElvFNaX7jJS8P/tzsxJoOx
+qnLiphfVkWUBjjlPI3S4fK+cDg4iktAmgA+TnokwJSr0M5IF6W2iYrhGz+nWcWlz6Ob0SHGJKXK
iWrIGLUxVZSe6QVSfMWfmuakOTJ3HDXT7RKeofrN46wNNbQu4mhlqArIYXtXGwTtA7F/PncB5Jpw
+IAALBkZX4zZFjt+byeCQbYYLH0fjK1aWeY1xJvQMZNHCOrnjJQMJNV7LyaVSdq0I4pSAGwt2ivp
uPZgpWF0Ntm+QYG2blQWuwqaQKT8bJTnSYfqJgAGtZGfR39zE1jwiNu+jipuyxm/6EeT8DAXCOHQ
KrexHfP4t5XObSj6A0p09IZ0e7ZhAE2kpyD5xk4zjRvfCJywlUvUHQDY1Gm5WN8QtVXBazrc/ZQc
7ElUrICAKjldZZtwNDNT0SusbAfEYuWkk3UkJb2406Qmzhh0B6BJi5nRuI5bhV1eG/z71H/OMGCx
hc7UGcDHJBHogycA25P7IEoA/vu9lidFhVhZPe10aXSZwk9ohA+fmPoM33LE209GmDBMVIyOTWOL
J5pd223kvMYQ+1c0NXawkWqU28HsWc7RwTaVBqsBDlvhH1CZUXp4AOk3c+hxt5/oEiD3h4xtQiF5
UiBOqZHsWT8EyX9IGm+ZOqm7b/JY7tsNc5YwmCmbTpAhHZICZN2jFzIjWuTOfpnQduwWVX1y6lGT
I45gyBe4sPjYVlvqY0vQ/y766041efy9adSKJBVJTWB01gUX6t1zLg4YXu+fMAAeC9Utxbn/qt+r
yqobGT0FprQudvxvF4S3Vrvb+NTOkDYCo/IjEM1GyeFGsU2Wf0YlFDey9ESTVhw7PxO2A/63/qT3
kPW/W1bCU5LNcRASQrGhrOpDHW651PSrtCGD3A0w1mzKM0Zk4qoEb1pAlBE9gPid2hkA1GJu0kDx
Zou29ieYGwYoa73He8XYu6HO3kW20znBBTrjsMUvUfvC+S22UMlT5WT67oGfQqJA5gcI9Ms7Qd8m
XVP7nHcboU7AmLYHudnevAy49iF0Kv+/W7L448bDB4AvR7xjTQrJ8GHkRBbNUDn3Moih253OTIUd
HqJlHA/JVyLufb01Ne6MchnqpBnCI0Ag2S6+XMdOr4ggS0UOA4N9cDd1+KFbL0lDTeCUiJpfIUQc
wJft1TgLunhCMO7WS85bgMQClJVque/XxpW0MZUPOoT1oT9ESIGGJZ8tAZZ7f0h7pBxLK1wpar1P
ycn6+xqcQysrhFxfJYqrwo+AeOH505ib9VpT7/adToWBPDIPNa8cL8t2yTnisu76EVqzaWgNQRFV
X9JpU6oRRA9AJZ2usqPgLIXe4zfQjN4m/7cH1Q9i4CUCjyUnKKhOo7OmWJlROsMpxjn/9xNGdWWh
pqdr59DAR4OzzSQ4aqoTeMtmhu+Z+QmlsFL4qo+Qid0IE1rOTks80SFL18eSQRUg4azzR5wqw3TN
JVHbjzF+HERgrYci8FAtzsvj5yueIPNuSQBDFAs6woaL89yD6l9uxfQ/7paKiO0+cBSwIWTrsVc6
VmSYqrij6XaQQzmLCHvkyJ2s10atNdEisFdKrzpoe+h9eWeORIC1Tm4gbCjDroIo43lWEVUQmRs3
xhmEvQQO8N01A3g5TuAT6OERzjWgPQ9YqaRfCc58yAahRSMwJp5VOrI28knHz4OnzKuVlfjnDr2b
K3XOIEMvE72kaRO3M43PQWjGA/fYK9gW3vBtohHcFPu4N/sGfGGuHBdibceNZweQvacTo5H+4whg
bT7L/p0lUd6v8xODmmQSrF6DBm5QBPLznFkB6F+IkyZ3kGzZziZHm/1hol7ttBPAA2NoM7eVIzwl
77aGCBkGa0iNTybHkF5WE2xq2gEQtc+YaiWhQhUh8bx8DKThiJZuD6/d+mXIJhw7XcpfHRO9RGww
36VporvwoGZb8xrgihsOXI9aUWRFWrioKLgE3ZOMGNunc8W/qBFU7W/Lkrl99vYX9rypCibQlKbS
+C1QYQBL2GKazwlLj67rIBW/igpG+j4YsJ26RZ1pjyZWunPdkSBt+KWCcXKSqlxAX/Bn+UmBg4fV
jH07KcnFwwEczd+IpTQqSoxRO0jdnInMUmDDxt58CuEm9ll2lBNyvoDb/qxjCsYwwkh5Laad18Bb
HV+B6EEG9T4oEeHxm86JhY4K1fEXzblMVwSj1xnuasemb9WbxPhubJssxa1oGor4sUH87mopM9vN
/JPHDp9Jdt+JgrRZy3yMvYpScbej5COdpCuPoJulVa+NndY2ERd6FGoX8ajHLwmowRB+/vgUK5en
3mcMofr5tfgIHVj7CDP9jG3dzKUHSd9mg9kzV/Pf/unG9DsYBBOyidaCJoJTj+PomEWZ9CC70FpQ
xNH6LUM4fQ4l+wIphGE/0fN9AY1aLINrUTy1qD1hSaWz3it3XGTiEiPbOASdAbVoeexUdUzZwmbF
vTFJNNtgOhlCTaw0qsAePuwbqK7VlPrs8LmU/CcoAQTf+Y5MXOo3o5C8LscmOK1/wbzjxu0fdeRP
0AiCDOGsWkB1DlaQIC4OrpJz7FmCQjqQhloqH1dKz5X06TH9be4/ag9NEvBu6pU3G7Lhven3Fizc
fqAO6kM54gHvvbrW3yLRKwy626PLYlbI9i8m9seVhwlcoRyuZ+cX7JcKrIzQPAmE7S/khgZ7nAJ5
xhAdAu1oL3ivSh+jAAyaaMjcIcDSpI5vi6kEzOhliT97yG9BeqK7W/B0vrHKD7BdVncGH2ntf3j1
YAB2p5Dl0zV9/eeQwx4OLqxkYxa/gZtkFlyBtLoTXSOMUdfoHppzJV70IEKcJ/R+FZ0BE1HHhZfy
x++Bvsri6EFBWPrFgQlHgYqOF7FUWCcA3n+dSlOmakQJKYnuvAls16IvYpfYgsI8qIMbaAVZBavR
ROdTcJdUD5wA72x/jp3a9qtQxFNsBrAooOTpKKTak5xTn142wWbJ8EBZgeu1W/9aQIoT86XGTYul
26p+RZ/A6Ly4kIoLCG4r3oOXFK4qUKj7On4pP5Tdc6mEoA2AT1IztTOgLHRhNnZZSUKSJ3ocf+8A
1VxZSqjnVuDtHBGFj0FQnjKrva/L10JOre8pfm295pl9Myh1MnGPIDZ6e48rnHMfjxiQj6K3WKV5
OgdEoQ9ZX27DN07tg0tri57aMuLDxYnrjmBVWm7zh9xmlPube7IclC35Pbd9CGX3Y9EF+0PDjh+i
dkStQnNUILbisycL3+cn4ieUraDLJqPMTHjTSP8cr2F38jSUnxQZRxFmbHA5KQZcfWMngOmkA0MJ
RBL4p5ErVQb9s9mMj7r/0dzwerrwHBi1vrjIjEZnt7sFbMUgsBSO2XO5JYMGXvmOuieuvzPwWWEG
mWxiJ5AqrOHLSsZYgjy6cdix245sD9E9he9r7NPXHvw07gWsQnUfbCx+ZDItsa4vlxLhUyDlrQcb
r9kzYWAGlIpgNqAwNGvyWfMJt5fZT7pnUWvQa5/jZTiEdxOW9DmSCYvo4a6PWmzHrYmJS//uR3VV
wUBH+rXSk4Y2h8bb8/XZ/X8s5iTX2yJZRtButzuf9g9UL2rte/IT0s6dFsnLcygfL7NDGVIrQ6QQ
qXtS1S7i/9ill7ar71zsgQuROTqnSQKdmY+oe4TvpBC/7BRUyZxJOUvDTavt8FmmZ1YaMhYTjPwB
OHl2/06B/AfutiZ3KBJ+VqDs9U7BEMkbV1LPZgR9cJDARDDyibmSujWUpZS9vyQUbR5vGdP9lwbH
4QFhoNpNkzq8F8hpWK+2JHXjWx5Vq/KwGuq0WS9iCLrs4KSboATpRoCZ/W1ZGVKC5zmafan85Tui
NBVaEpOP5DhEuHQVX9vYE7FFVvoEinoLIxVAr6tzA0NpNCfG9z4kSqyZiMiHnSM1Ubpkln52McVe
mY/lkLjgRz+LPpXopYEdf5mhQ98jVFLHr09ctC/k+nzV0RKsfsifZsXhp36K6YrCO39vH3Vg6Qj7
De4l9iyfzvgHLEyjLkXiidw6rFjVJItuSyvBGxnpNam1usyWTN0r7N4y3Hh5Ka8C/+F1+s+2HHsT
rtsUJjNk24MOCa95cvfXevA6yKyOxBTXyzWK+jmAICdIOPGyOKpi6d3HN6AvwetD0XMImvAQuym8
yhGN8cN9ZZugXyJpkXFesD7GVYdAFxww3lVeKTIvJNAzREjWj0Fr6OT/yUBTqZ8gVhGc4O8+d9nf
bttf41lyrvHLC8gmX+HGJN92ZeRO1Rbl01iAYp9IqnBXh/R3FPYR7QGqmgkIRbBRzlfRQ0y1Pl75
GAJkSdbIVESKdeQcml5kfGUi0ZmygtFKnSl2bvWnf9WLDOXPmm/VGphMBX4QlQF8gu3ozjR+rtze
90gxpGVSx/yEDnRU/eDflGQUzdI0aQV5Og1e3gN83xDntVjo6akvcg908zUco4prLX4GUv81yQ4A
19CpMXYDfnG/OAPRoBsDMWG/BvHCAtSfaV2yiRkZIur3FpxmDN9TueVwwhwKbclgoXdPKQddtaZL
ne1bZdecGs2bJ0cKDU2Gu315lpNm8yZAch6VJ+vNKiyPhVcYo+tZK6gmMuCyv+jbUSuSbvqSMVy2
rDesW+ZQf7OKA7SqQ1W+Gjw97oc8ew+cNEEJ0NTMGWUvK1dPFwjNTHAR6aohxNNYd8eRZ2AHyiP7
e3PAkzkhJWEAsVOPL+Y9IZF2Ke/6YIfp1gAw0rt21ZNJ/j6+IC8hVrkw9IqBSpnegBe4YDn793AW
C33tOP3/NlAjRKQO9Z8xkXxV7MzBRmMk7Y8nGhhYf447vAtiPZ5GZeOBaY9f6bIvx3VfeeN6slSB
H6lw+MoIQIFHUJ1NYRWXay7GPp/pTvL8hhe5WebxUYvEydj2sibDTnx16Xu7d6LTFAnIZle40UZs
2TxcU28tfvvsH7NLILdoXhFKNi76b7XgIddY5CHevp+MLBkr3jBFQWB3XXc/fHn6ZhpuwKGWoCHn
jGZCsD5uJhFbK4wCV3Iuy8/SSrYlMTQVKIUgHn6CWeZFCqdqkNqDMbGvm+o14qEpgTLq859Ha7vD
FhZygqSsVI7EItVZAvAxSEP9D/ZCH4IaMLzvQoLyB3Dt+LuwuIlMke55Cx3N4zBfYIY8omO77Pi4
sqvn6xqTbkrxbRuHL13wKaDU3mLOL5fkUhq6RIoSo3UOc3paaYG23QXvE27foxY/7rDVqdgY0eGE
EOcq6FbaoW62ePnDaDd0e9KG1+uRY+cBzzYwi2vEWhGkhVhM+DCVXu6JmmmLdUolPIaDg++2nO7a
kkAHolI2/48O78QgFcNEn04ZXESIaXExAlAI+bSl4bEFtfNtyzjMtBOPt5b5GYEL3EQhuaXd32iP
OqanzT3q0xUVrRSbRRKZUqHkBril5EjWeMhMFlINXU7teioARltOTGiVqZZ28X7VOzNq0df0ntWs
pUjEJktec0ejFj8Fo+0mJZO+I6CndSGkHSjOgjq+KuCzm+XatLDnzBBte4EQ+zPbEY5fouS0H+a5
pj6Vh4RQP6wjYXFqCmSe0dwNRbjnF4H9sFFKN601tIWLTXWTOalptIcF8GDzVybYcVnfRyPDdjbW
gONt89t6WehfjXYhlm74ZCuwEJR64exCkXHEimJihUTaO4R6IWV2sFlQ66gcPRgK+QhoAezJ6KX/
JhWwXAoE/aflmObO9E0/BwhFPnwkLYw3lU7oF4dWaqsKS0WQjGX9icd+UZZgR1E/jy/1eh57JR36
WDYD2GY+6H8iaIkE0b4fagXwNTJKf6wlg2Wko1VloGw28+vjeXuKRcEJ2cS3kth2KORIH3qa+x+E
mWYtm3KyJrx+RicSG+xgDvKdGUL2IoAFGjcsA4JQNzy9CCKKm3zKwMsgPAJkvUpx00ZhyNy/WF1D
WyRK7L9I7dZrFwNvw57Crgek8B1PQcnTVQ3SGUnaWH20a+PfwGaZtxaAu8Y+FF4euRLYOic4G8NK
yBzyxVbt55biW2+5b0ITglgn7OlJJMzz2xepJ/lkSOsq4x4ckn5vlrNQvurLfIMPrTsSekDqdHwm
U/0rswYcdk1TVJzGFeUf6TXnKNFCb3E5NbtJBZVWWhCR2IKZKSLEqQjW25v2bqpcfY46rD+VQZ4x
H6I3oWIOj92j/m4CYZxFn5+ikvKzQWiNIJj2KuaIIWzy2iUv2nBswQiIAQerAYSXGiqOauK04MZ0
wagjrf8ij85oBY9iQ0iIJKjqSpNeuMWHd4KatcEMCVgn+9yEzN+kByfagodJFJKkyXCJHRhRmbMS
wnsDZCvFvZYUikieS0OW2lobZxkP8g/zF7yDEtRQONt2aSlYWiHE3o43EhathPL2ku0wKabFfUJl
avirrUYodS8K5cjM2GEA9G7Y/ESNCqLJ3TNZB+UkPBTSeI8+GPFP/CwwuVbe4O1EnL7B4gheyxcl
aeAXAFXeuW9KCMWZbzCd0l4bcnXyNAKygaPmam3b2ugm5cAOzrkXaXEdnY/J5txoiLgb1TeLVnfu
LiZmptefCxj9JZoV/r/IQb3VyiDP03RTYry2lJQ8qKhvmEMD3m5yzqxeSVS/HbfajfrXwLohIirI
6rHIj82/eKXxhHYd9/OXaL7C8L/JkkFt0ADTHshIvYjdGxP6aUbkU+SFrUj2TA+H9kQL33QFLYoG
rkrG/PmeQ/JS9L6CnjkjZsK92hciyTcHoA4UC79hNyMQeSVdItvbqoxALazrveuWzwa83zlR/p8z
IIfb8mqqxH6ourSzHvXQo1jJYyDGrg73WBWFoHqd2J7yTnvu2pL71cneKwozliVHddhhccMjk27D
xRue6rRtOXSdL6tWy9m1sXJpBFeFrdbkmmIwFJYLAjyg08W0XIut7RlIhtvZNecPOZnbmh1Mc9ut
/E4KqLqC6oUojlE/uULJm2bHHJ3Bkr1061LWVHhLbcI0UpAFSrJVBT79Q4ZSDmutkUqjp6fkS8yQ
9V/JIM7riFnxI+yvmoidVnLr78CfjfL1+nfvC0mLjkcQaa+p51VFzSEs9dtZ2hLGFYM/Eh2fNBJf
vQq5Dltxuv23aLZE8q++ygrCJ1F+9ZgN4yf+QWcRp1fnQMPnOY6KD8hzAoUZWGKgBHWxPZRMhhYF
QGc4QefUcceW+gk0TxJNzbAiMujKiK3KvFV7rjWTM2PRXr62+bW+RlgiXAK/uuORNCEuhAwOrFaz
cxwv3Ce589Zt+TcH3leLgZVpl+2EG1f1XaSDpyqaySmXcGaKiPF/AO9fTgkMYb1N45Hi2EvfiYcw
hyQod/eq1nQiSmkzP5msQzqd/FFnVte4jxYF5hsQuhM5gzJZP2C+41xqC/0TpGKKM6AXm71o3NBX
NeJOz4gT2FzYOa2Yp8G4kJxiGVWkR8NFdKItnD3EHEakVKNOzeEK+SI6s5Ny/jV0g7U+JxyAePmC
5UCJPo7Vo00zJYKF1JzbQVKEwPkODOK0kJw/u1GB63M+1Q8oAwg0DCNAu/TM9E/DCBZQ33j/HTgZ
e3qa6HVZ/BA8FVtIT5ZBVUvTgQpxXfe2GmRaGOiwnp2FIXnAFwx7awVPvAxfcAtTZM28O1lJV1rK
tL0ERnI964EpaMgSsDXNDHvMDhEKiiFrchTBxdRGybHh9FeX47Up0X3YvJIC7bU1rMJFjba6O3Hb
ZyBLY2xCW+lMf3fuZB/sEx0GfwpHuUf2FomIxlYpKVqBcQ1KoYM/ZIZQMK0Epv0ZoNIVP28oNt0M
jPj15L/YvuJkcFZHR6DjMcHYFpkXEdK3xPTJvPcfoOdafHVfzFh8nEmQ/uTa3iA+nrHsjfKMA7pp
T7bN8W/CH3DtHD2TVm3nl9Bp7jhvdDAS75RVumALi+aVzj0uYhY5SBVM7MpRYPHrID9qlV6lDTa0
8URkDd1JMaaEWNOXYVfWr8+2ke7pnPkqJbatRoqCWq3DjDFb6XjEsz3qfV/CPagTNANhKmSzigeo
rY0kIK05zx5VobW3lwhyfw++7ToCwwZKWJPhM+b8ugMwqKcSGUK3J/MkkiTgRLsNB3cWBwqvHea4
fl0V/5BijALnh4F/XWMra1WnLMM/PwdFi0xGOFG5JWIpMv+RgU4OmWVqAq3NrJvx8dH55u3ekr12
9/bckY0cdMcNop7yLBAOZ/3WjPC3rZJqAGQR3g9jd+6WJFYQiHj5N0e8rMW0urAh+NDo//78/1QL
broWfikdto2QHwtyb9VcpD0DxsG3Ge+cJahbZ+V/5AMcy+6s8c8FVvlfGlw+cTllUCnLRYWAWPUV
3tA7MjwHnHOYQpODj4YJB1gCzIEosMTfFHXkcfyam5PZ6egyTeTVPHlO1hBCA3Jq92qF+npm3rCo
eezaa95a7sKPy88S15K2q37emO0MJeXNUmb+2K/i+i9Ee2mKUoZLPBH5Y7KjFWmBLGv8/VgVsP/V
+PQDM22/7ZvgcbCh/LysL/EdPiUGvS9RixNHWETEe77Uvf+H2ppF832M4ecBnkyF43/6ZPoAIzH/
hcdlztB1kRehfPUg6S4sMz4Dol+c2qCRi6Cj5wmcHNSABaLYSUkN2BhvrV8t6/HaTXMI6DgdKRz4
e9qwx3JOZvZdZRwAPk/sjdjA5kofbzC0afWNF/RDZf2/mmOgJJXyb9kl6KCV3GFl4KTxGl/o5cy1
/HSkhIGh2KHzS65m/ApneAgqzV/rXHt5HzXpRd9KFXZId7VCZu0tnxSKthFB9lCi7+kt+ugBUKLY
/VZIOnVKiV0yOSqPab3SsrACRoGJ257XPTAHKWy0K/6d6cgYPm0q76N6MGBTPKuhVaeaC1pjqatM
f6Eh3WUOTTeCf2FN57tu5+RchgFbRkLSP0vztKlue5CIQxBqcuNjH8NqO+hgfaGwLGCImOIHxsYk
saP+qfLZjomnCcuCOBa8F0Qe8QLLsGvBGLydeX9GJmFZf/c3WAxgRxyYKMZGFBEu28Pw+Zq7IVHo
Zl2BhKHqniNGFZSD5rXP+/QzFviU1A4a4CdpMupOwVDNJPKGjNf4G2jI9aj4FNywHoN9LUZWRWN2
gIO6MhzxYZpaLHOMU/uVTni6RVr9lrVP5B+48nvazxychyYkXIr72oLB5Zj5b5k38xLvH5sNuSiz
SNoMgRDJNeUHJTkTy6gGqcN1KctjfqXzxUtz6d+89nBtAy3MRco65jM1YzyOnBHlgbS5SljMaFWF
XCM2DMtFayxVD36AWfR00cK2tJLah7o7CHXxbNbmVxFJ0avBnVebEpqJhwHTXeapacF6DA+lFPze
38AGI8SjIwdnFBDLv4lClPumFd56xfNOOY1cuNYVvGf9663nW3Q4NQzAYxyw9oduD0la4Zg/jkEp
14ssF0YF7Zn+XFAjK5Uv7lgjYH1rd7wGN8XORkm63S5zPr8ACHwstnnZD0pq8TlLVLYkpHaym4/o
e2b8I7xomv0UGVTR4YcTh4bCDOgLrep4T0QER0MvGUcmkzLMR3te1TJxb3+Lrj/JSQCSYJjCk/Ji
DFxu8+crW5ynogzvmSK25caAhTA+TsCFbbGLpOQUIyYepjCf1Ovgmi4sCXNOfzA+5jzXBS11jVI3
ao7Cvnz5msBsQZqSHNjYfTyqLdUasL4z1Ucp+0Ragkr5LT9WV0GOqxo8N1H21Sge7J3hXYoOqtxY
3oyTS8K+P08RN7RBU8i9bGSGEd2U+nIj7FwtRC2PSXDcjD7wEtvGxBrDyrgPugLoidH+5Ywf53lk
pYDEpbXkHX/U4Iex+BanS+xvrLkzzHfkNxVAqSqT4nedBveM8cd6TClXZUMofsNpW4wyiru0w95d
yXjPSRzL83/nZuexb+sNkCnQKX+Q0D50KHw6Qaf7HYOE2tcnaYc8knQT9QY4hmAFB+QgCSGDWxmq
ipPbY/bfDCDEEjC6be0mWtbduSPl/jbTRnDBSBqlWWGkhblsoejyQ4JLZF+hInJp1N7wPPcNAaZY
B2LDFgjbqI3LV8yTUXiFE+GGpJyLGzp2bqDsphW3XaBmkJAf0KgfW3wGl1IIr+k84ergGM5HKO0+
rd6vuGYTsnZ3l2ZJY0Eg+8SQ2CO74UfrQVz+dwsIQkrPPe+ihNPIwzjVGqswWsw24AG1ldwUz0+8
5lQ/7QnTRrQr8+EqRZfGIDwkQG8L57NNuZCFO8F9T5Nwo4r9oAii8d0lwwr7lh8wzU+kV7/ozf5A
FcXvih/oCmlZcFu2PeZ0FWO96OmXUeTsMmX0AgzxsnGF4J8j2TlgiwlK5RjB0ILMOKmRcv+P37Bf
Wmiq/OK+rC8tUS2fPD4xx1DfX3gjyQxWJk2cqYkA0EE4s/BfU3dg6+7Mk+k3AZ6wIHLBmFMVsQUt
hjeRnBbYTSy0QNhDd6RVGzKT2Ln36lZqVfh8Q639ouVZp6k5w6hU6xqgDu0hX91rF85V6jijM0aD
KjvujVRB6z9xI0Q3rV99XEeASYdrdguq6bN83tQDxbaUxQSmWM06b2lTmNg/vo9vyVwAzhQA6mPi
tFh/c0JJKmzQdGXrl3erhoGwg/lNYymLikrRCNersVXksuCCT9imtg5Au/Oqo30WcWFF0I8F3Shc
cfHhjl63C1R0AMAd8r1ffXzMPI5bvIG8XGolVTVGwRp7jxl1ZhwGXoSR0aYIUikHk/RwUYMrKTRS
fxSgOIG4qc1e3KSutMf9NfK9xbK4pCDHe7aAR7vgv2EgVYqvuHwvv4sl0+y+fFJSxqquM8tbyX3e
kl4bmWXMuz9KvfUVxuf38mgrOcfEpdsF3wqnvgNdsMyLjY/+U51opbo5YbOv0CIrfU1D2UPMzHJy
mxq7Fc5Hkz4A9wE4p83/6hAfR1lt6vTgwCgpFH6Pi9DssUiQ0bErHT7VVAGuvI5b36iaL6Eo/tl7
JPwk48bPeB/s3675dnk8S+X2kJGlgIwGtJmu49Iih+UQGhG/75iMwvYgjr87h9GlsrpwvA6H2KZm
6Ev1c0VQB5WsvkxnxalqOaCUdm4wsB5gDk1ocWbDL6FIwy+WVwqpz9FjDh7d99MngxqVoS5ZRc8y
c2M08Rlml+AXowXgIMECLLcfnjd6K9Dq6sKC/oSk/0kRykhCKpWztlvIQHmZV73pcJYXk2XeTqVf
FE3hchrC1w7wSRnW92SCqsTCEcOwIl44F6WuX+QXWB2KUKPR/UHh9PaTtJcRRdciyMX//Uja1wgW
CPlGRKfKFBCXQVgzlWrGe+15v6pPn6RxO513SD3i9ok7BihHfpjhPhsP4xupQBP7WCrBVzKsepsS
HNvB2XSUs34hB5IiQWdOlAaydyqrFt+F2qWVvJh+7yWDeB7KfzCX0glpB3b/4AvFFLGVhtNz1HFH
JkuhDoJ4aHQM2L+WukazC5RDarGHgk8X5RtmHcVqCICGAnnJa4O1E6i/XGcxmYxLtnKVqXBnPgMk
GGfG6huJ17LrWtq7ad+SY2EU+Z2Q5QAOK4M/UEEjp/h8L42f6xHqCvzhEUawt7Yn6m6wmKbJsCiD
C27cD7DM+4KFYtiF7LocUgQ/vDxTuOjSUIkscPUuRYreDIxAMyZba6D785h1uKOnwZ9uMC04byVo
V5uDTYfELsAO8+VNukVNmhBF/TS0vLtz1nl9V9+xAZ6SEhCyzXO1IRCxheCPdpg2I2KdssJvpCqv
UNfN3DiMJlggDbHrKrXrHBgYrOlLzL99DIWAlhB78D4QsJmXfs7K8cW+HH3geQla9K6WraT6bXn2
CSejWbwcx6Q+pL6mNnpxP5enEu+6+Z3vp8qES+JjA9hJwZDCZTLvv8FNStKDloa/K48mVHvufC0z
dXNAafKKFin348zabJjTeNelNGdtPLzD0UscUsJsBSoypxgEmjNHzrIoVA1VRpBs+xeRpYvf6Fqb
Hh1VJo1xW6UY7adOoLcuRWTe0QwerG3q4l0cwDBvxii9AZlXOb5kokwt7MVqhIiWwRINZDN5kIGU
mPXNOIYjR8zeYyam2XoMkXybfNgmA9KYNt/AnrGnC7Xyf9ysOWEDwFblDQ2IgQU+48woGCFcqBvt
dsSiiA22IcwuNEGLXiC8sj1yciKeylbYhAK318cG1CyQzOOn31EUiLytQrDLXgTe1BQkCijgDWBU
PWSDoIZfoCjs9IjzKmmwOD2brfUbn05R/5MVZcjY78OHPQmgif2fv2KVRLLhHDvU/uMZ0sh76BXZ
Lk1YzHmv4v+CHbVFoKh+4GCX0Dsl90eP7AnTs1CVlUkt7Du6A8UUaS8W9Pac0gC18xCGTtQOrLiL
gb/6aUpLr0AdaKO1oMvJiCAoPUFI1cARuGmR6MyijaFVWNbHJrUM4IY5i9maYXGoWUQHX0Vzln+F
yquKiKfDEjQSWudXqzID74JQeQ+KEx9R5yUoqUq3uv6B4wRVzk1jIYqPzArwQhlp0ecPXkKp8y8y
PtKpDw99HRio7DHP5ltKwIv9AT6J9HROJQ6iEd7muy79cTjby+ERMGJBuk0UFO4ufazm364aENaN
MSDSkmbMdUEwI/+sfrG5EmG37TvY4Q0MKXj19heKz5Tcl+2X6IFiWXMdY7gzxOWF5kSMqCF6x8a3
vvb8Hgj/cdNh+pzBMa869lMm9ZSiSEU5gZXwvjpnSGxavZUlnDice5GBS//0QNsEw8xcZqXndKTN
NifQgf6eBKLVVC4+r1cMMrUprqlOpPgthRVEsnJ/DUr1r3+zJsZnrJDOBnENpuZBhmbMwr34YAwR
GgXHxnyp9NEybuQcurDZd4q84kIF83Khjp3qF67rdUEnS4jdQiUrRbyAMpv1j09gwF9RcUSSBuK3
qXRpaI4Seb2GKCHCAVYkM48IRMO+D/pVJu1lRR/tisILovxr8Pg9xS6HetbwbhH7I5THkYRXUeyf
bTsuVH0ZB0Y+BcziMQ+h3Jif2qgpusVOqrnAs+J8o46tS9pNKzCwwQbUNnvqwPCXlZDtcisobHCE
czdUc2yjj0WA3iowrSa4Bu1UAXCBOKK+tVVe/6ETjC1FaUmD4BYhaCwZq6Q23auUwU3fFuFJ/U9A
8hmsoDqKbl7HukurkgbI81B619Lh1PEnj7aE9POwJd/EB02VanhTveYMpLEnZnNHe2pb9UiLTzVN
USqGaHHpSEhy0AqzmIEdU6P9I+84JOjhew36j+255mIiFPBcQ/7ADoLTGDkK5qdYoeJNn/guR7/K
orCjQSV5pp9OSgBEhsy6CSMMfPUMWExjFmjI1D/KPGR+w6vtXOd/kxSovdQ4WwkqkZa4KGBtToYP
C8/79isK6TFRWcnPac9wMrqXKFVa5QtALryz7WDODZFiyENMTZK71Fs3ikenxzJznLkJGy5uVquF
TgjijDUED4qidj13AvkYMoOaFawcHyRi7CVmqmP2pNzacWKqk0y3nXmsenYFfoYac7Dw562QWbqf
L8psG0WX2O1QqC7d6S36px9i76cPms0/DA2ELK8HmL21NF6lvxZO3w69zMuYOtmluVRiQFlJLoxP
FuPk/iDxWwt6beuuraxyoK2lSYKL+SbCOqJw2T618nTuKZbMUXkrZe78P97lTJhgGovRFyJ4Cb0x
ItD9TSm1KJCGGmGGZYv4Lk1oe9NetRffnvSwA+NWvBGG1X2NMd9dAWIFDiHg/Aq+KmVhHIo3dwMN
XTJ64AOKDVk6/BZ7t2uR/4lzq05eJLaplK65n8eJVCUjTnkaFofcinG5lRbXySySEgaQZM1NQG+J
IR/mnArCC9d2BY5PByqUghkktyDWx/v3HHs/mlsxxaqkobko8D84FJMaIs9JxvxmYaqQDrUpZkV0
nU41IZPtcRqk5qq5T1fNFwFikf0vUbncxH0w+8u81G0qaiBecu7tuh3hemR7PY+XwD1xfWmwaifx
T/auxcyDAJt008gq7U/Dc5ov7yGLQM66w//hqzL7Nc/dSeETdEvtwA4glGcfD5LmqEz4gBK1PlNS
56hxBmIRHhZ6Jxxjk9r+NZcDMDR3w2Erog1RCVIp/am5MOz/Eh2rWfVZJcN3KWj7yybBw9ODTJ8r
VbZ4zApHNKBJiXF/BlFakS7ANnW/02f5ULTw+8FmrPf0kSnI7ak+WIlsPcKHJvdUa85MoHMv33Q+
SL8r8jfDkxqhS2uh4uymtnN/AJuZyQagHbR5areQi20BV10LVYlwYByIN9fvUQBkYQRQCeQm62g1
aov9DtrbdmxLIgTXNNsy0snOTt/zRpdStcD2j6BW3AfX8Iy2K9+wSGwLIKT7KThWyNZONs+9SdQl
7aJFQn/G0Z9kMWq9I4nIg9IxUuqW6hVZk1DnNrU4ioFlvFIO9n03tT+r7/FfqKgM9SvOkpMTD0qs
Mi277rpT9lR8QTlztzIRsvEhfXjVSH5ExW1FBWpST/GGVMF36CfxUzLYsWEZ3x0z8a32Jr4lFUJg
wxRZaR4PqASi/+wg5YQ5spo+nm7yG0gUa9m8f9qHO7c8yeCYseXBECqvlR8OGmkatQkOQ5b02sUE
olAViF2iL9+VzLRa+n3ZuFWCf09C/HnxuCe18ByXAP/j1c8gOrEN9JL8aVcvmDHo/ALthx4RKzci
hgmxMd1OtG6OlmRCId5tCunyTi/aIDVT/hqLEboqNPQarVvjDZnOqP0g23T4IFiD2GuxQiLfChNi
zQQo6b2QTWd1od6UojjAI0DzqW+YvZBzdpqKtccHGOq4SSxzUQjkSdm8RyFuSBXszyVUoaKUaQqE
mvkulRMxHna/1BXbwEyi4Wmd7PpsO4LP8F7Fp0Chf/+SbMCyhN4heG0nK2Bn+dKstf/393LUQZfc
X5p3GXj66hlTdTuLdeo9YVn0ROQoOiiLWBw7EK3BjUAl7ZFSxlZhCt3OMmIF+tS4VAGD2jPsbvNo
w1WRF7qd7mwV8RXhaBLaZ7IVvl+9h4aeGwIrKBl79MhTGcMqtCHYXV02oI3uNtvL5w9yPgaTXVrn
MW6eKBPydnZcKvLcoen44EyEGl1lnQFRIr1aW1kHPFoaGfk/tDvb+C7wDUMQsNW9OIb3UxlyeXG9
ZYYzzrad7aQj08MbE5nuf/67V0oui6qhASht/37zECjKkp1/PCIsISFuMinXhz7bwz+dsB/Y0ZOK
k6tT0bji83PMQCd8hX4HM5tnFuT3m2AwtESxzUIHOmOxd3F54/INLd+UP1RMKvKSvd7gkyYiY3OD
k9YPu0x7yp2xQd355kkIm6u+CKR4+f5zs9losh/2O3NHhCGzri+oZkB4BMSDQvg+/7EZcOVI0wtz
OZUSobRb/lQvC53FglShnCNqhBgZDMBvq0IrtFIZph2COeCMGLqPbV3I9cHFH7hBlO6Jg1E5wul/
7IWkaFVB+XXSkzz8Aprmc8FcEvmM56XxX3u8nlkXUG0mS9sgGDBRHwuKBdZKdIK/5S61wmoL/6GR
0ouE/EdkFB5quxy+TuPD+qwUQF3QQWQ4GCQcz2qt+7nhMm3ij52ovMzbBIAF1g2/twwB0Lxdilba
3h48sd+heBl3umscfb2GgBg3J5UGt1LvDtlV8yCdEfaMaz4Tq8ok3oZpKiyKDj7rdBZZvVFTy3ZB
BTG/LN3S9PecsOKuvngV7jAs28kEQ6NYxw2AElg+2PkWZqsgvA3O9dHZkKUFmY38YwevhCUqIWS2
K5MXo+qo7wUVK5CANvc5bg+TIKHPVG66oTb6wdNrP7QIdQUDvxc9G/MBm+tDbG66GyEi0c1WCpN2
ogsXPItUUhTVD8XJqVaJgGtGuO3d4FICVSEnqG6Jj2Io4JME2iJCB1I/Bvo/Ka6rq4vi7smnNi6S
zOal2lSnbZkGpcwXKYj2xGDqERFrsart5z6oS/Jv6YYG7S4VfHV/ti1Je+jp6bytgSKkFVYNTpGS
DgfkeOlH9a2Gt42S2YVf70BymLnc2aL9RgK9PGM1Zg++xl3+D5FwwMIYyS4ZTX6rbsEDWOH1IocD
OYEhMjbQ1DXHnoJHAmlEK7AFsKNRsTn8oX2oRXBhHq2nKRdYRSQ67BbwtCnVsLiLJoh/XxQBIzPX
USXft4nJUfBwM1ePeiGAWC4RkabhglpJn9TbTi4cwLwYubl4xwGWU8Tuu4ZBpjQO3sndMLTHcShs
PLikXpIuRafCdDlEEDc0DOsYIOIC4HxZedRVL+of0fiMhxCcotsqSqxAsniuPBUElrRtWY0lTZuq
NiAoi+Yqzaw6DOcUDbfVvkP21j6cOFn4u1YNWwncwFr4wCohXtPFW7T4vliyt+94tjnFBlyfYQhY
xEj6GcGoDpT7xVcwOfaRKdzv/+lfCgXOLBzv12gbMzwaFaYLLHsW0ZXja2U2PXl7BZEuGnvnI7BH
WTLZGLQheaJ7F4b4h1ByyM75cDz/PQ5Tbc5GRgcwl7X2BBULklvV3zEHiJXOFKHayF5IUYS2Nz0B
HZFBNKFONccuf6+AbIzEI85zQ3ZuyLrEWpVlxIBreJqFhKXlPisUCdzY7mE2SnZZXCPRwFnX7+FW
ESy2ApYdMG2fgkBHl/EfdBseKMUmCte7j1pYmDWyUBc40AznXU52pVivDof3wbIOGdHHuVB1ED58
yuSAso4iyG3zdzs70RkcO41mtQl8adRZsXbW+T7J7WDBi7fDTcCoccDq/5dMUAmIgNV3E/zhkffG
peb7Cf1xMEaL+BGsNnPm3rMs/5mJDbXvXAYZcf5zrWcagbt6goxVhj2gFFK2MPBJIsCFjDDZpHxx
zSO+enlHbZYj2r5uiV8nOR5adlbdAeaY36cAfTfvkLkwX3302Beq7ZwqdcFcNs/INz8U3kV3bAnv
g9TK4hef6QCIx7QYYHt0yJ3FX3/7NLE9Vwn5+PZasSmeBEfykcgJojjuSMZsOE8NgL6YBosY14mr
wmNWnlBNBbfLOd0ZAVQsmJLTETkQZPq7lj3z+WR3YD2t1ScO+LnpYNSQQJqUMsEWKZ2fSkGDxa5j
nns5PWyOIL2BuJe8v97hu7R+0SDTPnZr63aYWO1o8V5OuLg/0V1YkV+32qQ5Zg5DvoG3yCPT3x9s
k3JL5hZFiLkR3guHtn0hEjq0f36k4zzI0UetHhZLCuPrA/5yGncv1qmj/s+QdkUv6XnpQiDUCar6
4mlVQvsanKw4KzIevy3WIIlio9z/iRLmVXBdfIEeMeHezXYMrdaHWGAX4fEPHgrgytRO44fn3xMa
cUt/sdl159ARQ5GyAEIwJFwS/9TBhhpA91b7kHKby9sZY4DUhZ1u4FP+kJlwJl+e5UEnoISHDBXF
8gTHZpABbDpnF47YPBHQY+wz5PlsN4lCcYrjyROI3OlR4lvqx7V49/bNkq0W1BH3GrTHuErXZ85d
ix7vG/37Ot32NIBgHUrA7RO7bPVhUWyFciGCk5G2+Iy+QpLiC/WNU3uGzRU6un/EqOTWj/I5HC9d
8Wq3TtzYieTQfeSocPVATMlsOXxm7coGZ5MkpvRwR9+LD770HdfHPR2isXqNdE/4F7HoBbNWZG1O
jBUyRE/f5ZOYAYu8OORj4ejCzsWGqFcaSiAldW8UPjNRClkX9hNBthlPSXtWYnt6S/F7OtKJrrX9
t8AlO0M5Jg/rpth5Hj/RjOUONBBZTYyhHDwCom1SMQq8YbuPIdOaeNAd0cfSYncim5JRdz8yOCQz
naQyTeZCyF4SSKx7gBl3w9+OgO9nYh4lqZwmubEcQ8wEjFgV9v1neOWN6q2hBkXiBWRIZPBPjzDz
g4/Nz0CYhFF7X/V0cPI7L5OKBF+QWfkqiT8atNfEsR7L9ioFyTfICpMuplMoxQ/f877MDg22DVaI
bwWdvFQYIhoiNSoJYNigwvcS8wqVm2oBFyYiRL9gJZW6euxRHqGfJ+beq++Gj4RFZ2KQsLAY4Wgr
m7YHUjZV0qHjeFimq93fQDWaSAg93upKshExWN+Y3FpC0F5VUtqWt5Un5NO/P2mghRpOJR61gGSb
74wr+cfwcKiLOI9Tlzxo37xlG0/8ccPn2qvYPnohnUTGyF7HvmdBVAo9C+JBgipNfYuz+lAMnqL1
ygq3LZKHGzirS6ipfhs9R1mVs+RGO4+lXfgL6+pRkLxb2Yoe7abr0Yv9OphuD3rPEz4N8LhTFac/
Do27OLhbCe1wUpIiEbPvPIOueKSSNYkdCe3Cf7uvI3ItGChj/z5qWzu1DnPdB59r76BzpE4Z7PEh
gXXJVhhhq5a4/kK0p+2JK0U7w4qvnLi/vO1vr2c94UXrYfhy/6PeYqZuGwFG6MFfJ5X8eRtC60AX
4PPEeK2hnLiALITXYiJNG2LLmmfoX1IAc+F2PwLIO0oXREkvqMegaH9koO4jFv2RInniPd/mAb0u
WmUBpKACOPcvNlvVJYNPaQkJz9aWH6Vsnd5TCnQE6zhB6ItWCNnnYlTKOOvJnuyn1KDl80/f2ouK
XVUIUmHD2AbvIXj2W6de4JHNcugbyJ9lio9iuzuXP3Jmgg27/5m+thzFUICSCNM/xU0kSOJQ/2m8
efdmpEWednr53OyWk+1PrtmCAJ6BJgBze8C3FEb3PwZ5l+pBQa/3T086OqpA2mapdmU/JCKYG1jv
Zf13VAon0Xp1Fo8WacJJ1byrwZQn+pHylMS19tlJXP7bwUHBqMc1J8M/Q1oUMcyriHqXbEeZMXyT
pLEDwpmoW5BP9L8tE5CVxi4l83bY+ynkKYNycvWGPSaY2iV46vqkVC1oPmp5D3r7hSnvbmF9S/MV
mNt94lyyxUXpHTKOk6EGikl3+8MouI+H7ic8bBHbvKxs7UHYamXU5ePsj36K/UBvnJ0FulmjFqrc
8IonlVBrhpr8GMMU/Zdxi0GUfzpPfhPdB+1nZw6d51klgEB5tAfE0ffBDY3zDYj1lvOMff12wPy5
FZY+DEGZDcsvWvldv6fxweySnoZTZnl51ejrRH7k8VYZLBz7V5Q1VPfbRHuc5qmLu62t+R5kqrAB
CT6ZYhh6Rp9wVVey6fCtC+KsiemAyJQWS8gox/eo1FxZQvWS1TdRZv9+ZnLn5H3N2pRD5dctIvat
QR1HCorh5GyUb7YYJKEdfvspNx4PXNStC6uvpAJ9oEN9xpjlE9NyID59K+Rg5d701qOnWqUqc46+
oDufPpO6a4O219g5rEvFZGqGfjdyeugWiU3sc6szk6qzMTFAJuCrVi1bDZTIuMzBlYyiCnfEkl1n
5/ZI3Qb7hgyrwE3C9qPadtI9MOXchANb4Tz2p5VbPCuAJyZjbHyuC9O/9DDlBxof3B/0+C30tz1g
o8BR8tCC/9VQSbsRI3/aTU37iX0wX7vI3Iqzu587lhHxTbWOIaIupTE/j7B47OVoXmyd9KUHqaK1
01qNfzw57sjESR51QB+ur28rE99J4IMxPsFaglOE28WmsLHmogEmGOxZf6FXFxRORFR5bqOhjNae
w64JFUID1wFfBs3C+q9Xq5wwmk6elB7F/a0X84oe8f/WvZxQdFlwItcnMtR3UpUUi9d7TdFq5xTT
YBm1unPSiTC2aeV4TeZ4KLqF2B3tfA+88dZHxBCFNx1ybymWvRtklZnq7b7Os3JT9Fs4c5qreTEh
vVkYWzhBmSY+pWheueXpzYrf6RBHt4oObuD12ppxVyGCToijCKHTfPwfkA5PF8/p2u/N7ZPnJ8zQ
QKC3OvWxsrP55BO8t/VlnmhXB6BoaXTFVw6/pIFB/dMDBJ94vzCcD5iTv/6GEYI9jMRHzoHy4O71
HNyejXyJVSN8jIyeqcNes2r8gwXDJHfNFZPkt+JKYk/Wwe2WChElhAEOvqoLwGPMBtXjv7eeZ6mo
D9F2sobWtbhE9+9aDktEk8zkYJktsdeCXP7NeUM0c8lL3geihmpuqD6ClImxI4sOy8Gdz7OLhg1s
WWg7T3T5VsTgJdEM2RNf9HF5IOCtlgfyQuQ/gNId7SbldOHsfabCWbCWaXA9hgYlUOHX9js0EkCR
zkzix+paWedJYIS+hyKg8Wu1CW3hpI8udy1XWIWI/SvctA32YIk+gpzoiaKacSwaZ5si5NTIzFUt
DSyRAF981GwkO86OEpo/pJQLPdF9WFf1hzvyvtGYDGE6oQvH0pDcjyE3KyG/ecfaNBzVfa1K4TSs
mvRwpq8FY0yZHhJhkZ8o0PZvGPfx4403dCUWOimw7tM6sMyucoBOBaSN7s+UpprHveOO18ZPasVV
Ur7y1UQpqvmQJMXn3mXZ8nIYav5PzOLzZPsHwjM9jjVihMlEkeKCMmB/qTk6TcBOgErR7HnlZmth
9bPFLASVK42qznks3Y5WNnK7wYJlRNuhpFRmfwEv5xHnHSvBYAPBkFgqCUTDLSzyd2sOpqXh4E30
yOkeJ+QK7ETEXPc9zQ4z+NIf8ij3RydDv75dpDkHpapSwHN4LmfKgQVvN2g58pbDgrwnvkIfYHjq
hBnqxAr29Jw8vRkfQz0SgArVGUBnbMTeP81AlVMFcRV6yOjeXMBK3u+8NIeFswfa9Ot0d+MZng6+
taYeGVD5uQEryE0dXpyrMZS4oxN3Wge21mP49Q2G3m77TcedzNrD0vg+2cCiWqCFe7maZs+AGVmY
8+jbPPFbdKwAzMDltiVr59gp7mrAy65tpRLxFCi05tpyUH/IApzYUopIzvDbt2YcNpdZcnctassL
suSrvSr0oy1c9JB9WFOp1U+79OAyOnMzkW8TsugYtH5T6ZlppwJWxOGRGYj28vVKiDnjMGiVQeON
hDqGktFqNRPrUrzyeFyBONtPEEoFHvlk1AH7eV4Xq5gp2HvNvSApVCtk8ADKxGXG1H8nJkSqAr5A
RkreTQBpkLBReES3bie688Pu2LxwSeKeeg2huMiqCDuqz7DKS01mYkI+ilc6Nf4tdHukGSkry5Xd
h7pNI3vwLec+Sp16/X9QOVWpRF8OpEPvIWFQEiqMATSxmB0EyiohULsajexj38SkZR68iMpvDb/R
9KnpQO7I7vKy2g55ftWkmgZcimS9eME4zUUqMjag+0Wb5kcpJkYZ9TlyCEZ0C9Wq6byl/etbbu0p
Xgz3iqcSVPWMcfcNDpdOV55aZVLLG0sYzUjRA03Bci14uHe6/fyBBXOTdIB0xFRRM8Djs/EEA7cX
W159xRkXhqSTnGDInxcpPoNG5+fXr+2kVGetCtQj5WkRTSS5KoKbSXcShfCnHTXbX4ST1vj7c88H
XGpOUpFrRL+txme37xcLcxJdIaNcxrD+SgW++0ANwwpfvcLif6tE00oKXM00M2MuXvxAjk7RAf5d
Sw28HL+8OF9DWm8dyBfjDbaecehD9/029h1xpYcFfVe3LcsY5fmzt4fu7Bf0sF/GRuEJJ9un0Ru1
oqGRUFk3xlCkdthB8wKlFvpG82SbRfWWg1KKTMqtoUzJoguEl3DwBiDNudaB3XgN5tp1VEe4UREI
XCE1a887XxyvFsYUF9xTEiqEOeVSnidMVRtxME3aDe99CvGdW0e0bt9p01C0tdNuuU7laKC6Pgme
0GHNt/JQGqtG1tZKoJiwwoILj6od+AqrlOoLXSvA0n9i/bzQoszU7oZHBf58LJfJkHQFD3qPrXVO
ECw7ErDufWoTXak4JfH7LZWLohDaKAUbvTfuzXhJCm3P2baxBJ/2HCY4NE4obxAY77QxlwN6fT+Q
yvX925WumhmgIEm56qVbbEgP8ct/5ZkHWgfSt4RRyIs3QFDm9h4w6yuyN0ez/HK9yVpN9RIPxWhV
Kn5he9pAKu5yxuo0rn23SWJDjd1NCvgDqmzcD3c+IQKH280p79kWjnvnC8ygtepA18nen+Wjmbj9
ihT0T9zXBilgsuhx6JzlCYj/C8EKh7W11xT9fY31HdjJ2njZyV2dWMzghjLriLDUWWa/ZmB8Xq4z
oX8peVK6OvDi9m5/DgJQ/Xw5KP9VjHDvXDZmG2zvVIwuUowxZy8Jxv18cfVvb3d9R6EEq8/pfCFV
vWh3ooGWc2jCi1U8gN2m37NmXDNJra3luWAeIak15Ad+u2LuIbw8OXqI/d0yorqgbXG8P+8TPZN0
se2MiCynuBLT/v7HQfZjI2Vdm5VZp2Yxq8+Izilswu5MzL9MaiRKD2NcT2LUwysiwR1ShYEJuF51
4CH5GLLhMakg0GgRdvYOcAo0xpW1OQNguMHDqFJfYi2pidZB9K2xzR3VT4a09T9trumqVBdpx7Ct
9uhdjh4uYreGXQydYnfl4XDRyDMjX7wvZQsxOcbdYZWxsqUVDWhWq7yjH5fzEzb/1MyYNRPE4oop
kx4ommNhfwYQawrB+5hAScVYNBAmZpjFVyXcfAitrbu5bOR90EFpDpuZR6LWYej0fXrDqASpUbni
q3BceeVPGmUnvThNrZfhdxShv5dLYT5a1pUtX4aD5IkZhIzHQKwTj6kJa03GyXK1l74uAMNTaXMM
PX4o4xxkDRS6ccYp+zi+ZKQt5QE8undm9g1bRmZfIT8n7hTTo/Q7ajbHCME24L+2ce4/ZxDOo86o
cdWdT+YPCtxSxx7xc6Zt4sJmhx/D3ockopcWuavjk145hhXMiqIGweE0vbsOHcodWfKI4aX5fmu7
i1qCVsbMyWgChHbD1gWYRXn06fqETjGig+sb3yhOv0FSWOTy4SMVZA00sundOxRxoupDYfxU1Nvy
ZJPAHFkrEE16sIvAiS16csVfY9HqphPwV3JSBZ1J06snqnS1jJvISSFNuUTIjCQftuJweIDBYyUb
aAhtLPZ8Q6fGjrrXpXQN4QlZbBuyzLlBIx1JNMkyWkj9rJKl7EK+lP0deKSddfA3eT0jMi1mmIdE
3grgUr/+Id6+UKH6IF+ix4zM9CrLvj0jaFf48e3iNKGbkatfMx481F+WxulAx/6Ics4NW/4JPsm8
1eg0EpOAiOISxJF85P2/lXbH/3sGT72QTbObOnnMBa+w7QKuH3Y98gOg057BaN41KvvnoH2XsFpV
UGCFrqZm8TvgrR8XQPb6dF27VRuWvxrPzOxo0Tr744RrjK5ROs9rEGWh1zBULL4qQrXwKf7ZjS4b
FFGIYETS4Goj35YropTjd/+b6aTCYZUzsbFrvMo1A2NaWPNAWgZwAN6VmzjK4n056/7TkitirlzX
RquKG8TJ+5fCj2bmtj9Qsa1GSfiMG/OKAgO1i1lnbc2xpZdkHBlfhFcRg5VWuuOTLM0fyRxL/X+C
05QsgpnHDbTtEcAEYGFayoEZP0Fx31YG4HnGUHt9wdxo9AQTWIT48UAQxzwmgaEW5BxNDzD4VDn8
FSOvB76/SLO36YTsUuOa+L5EGNhYTSqF3zhyRm5CWKVNUcJvYIGC5WjazJz/IGJOpat+bIDFO9qi
lu62oNwahyB0ovOnRaoryqDN3fEhjVuGalXp9wxke3T6yp3+4MFMwutUfYolZCvjp8eJPUiD7Vap
iNNBSk1LPLWNhIOCLEOb2vlEyRm9yiygLvIHT4vRi9+wieaoYZSxsfRIbkk0m3chpzMlXAL9AFnl
wN1N7Xv7K3Hc3f7cLS952hGPZ3tLVfqE74HyMn309Ni/vXKx+Y43TTGy5+xqOcvdwjmUM6nQ41Vj
QSE6S7w0J1l+6r+c0AOdY0ks+7+6hhBhwNEOOKs+DtE1ID0NUMHNqZdE/JW2FBV/R7tawmRJja+R
c+EelyHDbIxfLihWmsLX6ypTxBaDcTzjwpWP/GnEl7DkgZfYFccFXBIh9QOaH6oUCxepoQkKI2SU
J6qIZyxm1u9ZvbYyFQYtN0F+lb4TYIvDOL6MFwWlpIsK89za/Frk0FlP+HpdNNY/a/kgmrgUjbRh
30glpBnpJ7lF+LNXzaVN3zdDfgDTfRR1slvCHIbzmflFHMSdtT6Tz8BGRGJg9Fc4L790y6eRiz8X
EV2VxaqrzQY/+AGhpvvXE+vDEfFsrD5RWeSQzWXja2A2n8Yu2YfRcOpzZuh3Vna2MLIqepGLRmZ1
vPb7/VTCzgwWHpbnw5SxEy8WzNqMb2SfV1sJWyZA9SBiyamM24YNlrYRo8ipostk1qNxkbh1Xevf
/6pnnlpIt42IGjtg3GjL2f9Xa7RCmjKh5FyOHnz9O4sl+S4LtadrBU2iFRKvY6SLTff6FrFUPa+i
lys9DfKxEZOPRNiG8MB5WYaMViF3GFvZUXX8BaZeNFAuJg+v9GahtN571w+ytNdPQ7EFeZfbb10S
VvdSGj6gG667lAxwFnoT/s/Dm5Y89zg1AUF3uQFV5P50sZldlbSUZg9dou2O5Ij2eZQATeo4m9K6
0rvqwLDk4qnZQEpaJ8L7ZwGESuY8d/UL+9e1gU279FJXIMhWhW/1l9/anYMX/j4X/UZRJLIdBJkk
L8Q6fLvm0RmgBryi/9b2vddKMBKmmKL1i95XBRrPEmpdw1xBCiUUlVeye3RBw8lLDJKOWm3/niBQ
E11drIeZYWng+PwWo3MLOaQsGPqB9pMaSprr2e5hEt273gJcmtqoZ+J+gWHuvoWY+kBRa0g5VNfI
a4aR8b645VOlzsQGdtMQsjoMzOq2ioqavXImBql2iQzNgEbS5JAfn5JP0j3T2XVcrM5FPnR0sBpt
d2/JZkE+4LVw/7Xfc+GukOJbS0oLd56WqVk2IJzQgWokywSrO0fiYeVmhzddcLiLliwMPbPfpsgs
h4Gqbdewf2MVGRtWHFHmUDXV+yBzxmVNXCk01W97VF0YZDoSGGrj7CkbhcnZo/UoOokh95tlVTcn
38reAz57SSHghIbxT7nBXD9QISdOXDFMHLhSPKnIExiZhsOk77r5QPlJmngadkcwXz3lyP34jJ0C
Xm1C3pha/GmCU7FmIQPLH4IOJwGWaVY1iduMKiaMxRJM/WsV/KQorfbckxwJTjSRdd3i2oXfPHCq
E8EXSTvaU4wnwETVDgICQxdZYCUyb0h4IiZFlj69U72iIlH9ly5Dp/MeTE8DRPPWqWEvHQnhI5SO
agtr6sdEduxi9gETjtkbj+X/W5UZF0JOvgJ2z0pz2DYcvYvbFiwavWsQA6aWwJ8vxcwJ4dVPJmdt
7iVSAWAHAiZZ4oiTDPBFMeEw5wF2IXV00BR0gERbg3FUPAzPODWvuTUH+glKfXW20b76sqs+m0kr
B7nJglquVv0dQ3G4m/IicpDjhQnvx6MmEU3HT/YyQs3ABHmY6ZHg19Wr6lSOMNX+VP8z6yBxumz6
Il7dBKV5lIAyq1gl8VDUDoRiasBTHZkQWy4UWfBOjxBTiFs+QHWERrstfiyLh1RFWKj59IL3wF3J
m3jrRG5HQUhWewh5MrCCS+Ua7aM0+xHTyHQoXS/b6a1oF/HlAx6lTeSw6pMMvrG09cx/ljwKd8N+
resaopTdYmutXAy3gM6OHuOhR6GO07fzhKUmmKV1LzhtllOe+JgJCzlI39xrP59DeFiPeY6gA6MZ
l/VirIFJcoXd2KoHi/lqv+LlCNTCjvXcI8FPwl5a03O/ZG/kWRYUdnUuZ7jm+7XRx51xU1hPTBF/
HQxOTe64Lni4OYpS8zi26ijzAhENI80RBrN99+eIwqQPZxcr7KiQqN3NMCAJfviC3Cp33TJUDwIt
pB85ZBo/bDHycoleewi07MSFGDVHNhM6DT7bHC1yiBxJC8l6NpzVSWYmmShMGuRLKlxZIowwGUhp
5OSsOvLJEhyArqLWqE6Q3F+qlVSF06/5VMpGgPBqVnvJOTIFW8wSRTbLIWn0M+cPOyfvSwb7bj5b
U6nGze78krw8JQWowRMf9zKzqQ0vT2t6nQXkLNJcEOhJVccXdUNuT+MjzpIdyPwIJx5+9Tle7Kka
SYQK7J+FaD6ToF8Qdq2Qx+0EEScGjYsLMYxI3SYl2e0LEbVe3/QQKizHBulcjVYmqN071Zy/iMBg
hQJRiVWKfogPKC6RsrvBlmLwQv2Dop3+NRQLr6bUfow8zAEVS3Hoa2sYdX+l/PAuQXjzn3VU/ECZ
PUmG0rMjHmEf7K3dgFjxLb1reP2vDo6BeqjJD7mKw3i6YTlUM449dJ+6l/bjzJJV+l7ap/T9THky
992B6KnNOaZ/OKS1FmAXFvT0Xz4pP/1+m9QwvdrkI2uoWqlZ5w4uxXIQPR/lNcFJbl2ILdvz1gCb
jZCYf960CuaDRDczVubQghDYtyehnqPiEiORExtm6tjlxXmwhBxj1jLQ0TiuSgHXjQpWfDO/Q0/j
flLM9AsRRv6ryQREfVW8LOrBxLlnVFqY9+I5uY8ynNdByy81M6CZaQctoN7fluasxYap7zK0rU6c
Dpysu+ihUjLksaH7c5YfsxRVF7GNNd8gKWkhuY64ry8lnhD908VoKlbDWdcN22/vNuT+8yZZEUDE
o/vIg0X3mzkH4AAegLozb2fEkH9o0F9kKTTolI4+5OihMhEixMZVGRIXY0vUdxvapTAHcNpO5g8H
/webZq75/YqaYf4Yc3IWIe7KnIzOMApKmqnKjf512fK1EoVwbjPpV5QQ1ChYF0vRG4lBiQjkV5WJ
OPE/IEUGNc+ymP9SPfFktOiwbbLo4qNM6yHDxW0cThxlxqRRpa8ts8tyqwaawC6rU97KVzs+Af63
mYZvnem3xv/6Yy7j/AXhOTS8jBvqJGZo9RHYE2xgfHaYcdT5ItqQDZcntkBvkPExDoeSDXU8wKWv
iJOELxbabPg1I7cDuZqhPvxv6RXOuHDNItt0qEjafjdca7uAos6H6KVca8xrwmJfy/i5n1VsaccL
ha/BpjwJ5Q/INhxC91xK3RTyovdZZ6cf6g1D/PazeeAC7DtaHQb8+aNPxs3SbNMs6Xjte7yZIC76
j6lGlPOqLGRC8wuHBL/ul07TATsAfYKFb1Iej0S4VnoKe4A182OaUSwiazR+7aU+Ho+xgMEnWsX9
gMR+xecq7rXTrBm7wwOl9iM3wWStqEO3qGZHq0z3VqK4OYbIwUVmi3TqCmusJjvhN4pDp0t2ciT7
OgJfa/tfyz1DJzmOPg6Ja1JpklZiOvwYRHnENLBKD2kpO79ssFJjqb+lTMR/v76rUui5HeoeMLX/
DOX7M6VN2tsIVj6M+IlfNm03rQvgY4ziQ9kbQdMpR/qJUvcXsty7Rq385nwCCTvE54uPQO8S/wni
/EK/c92+zDuyiRO/HFkgIPHOUfXbST4e9wUVzAg7+BYQLc1opeJnSk1iEV7tXQcQNQv83IF74n8E
pzxAspeS9iVYbRDsqTHZzpRA7tezT7GyOlTJ8+W1a/wLw2IUAVP+v9G6QQtdm9aGc6bhW7OAfBw/
7by38II3NhO7s/qsLxG4saS5TrI6htLgOA4eFEcfDZw/ZMjaF8U3LVzZH3fDeL6VKO2LZKxsI0/A
u241IuovemyaXkTAqeUO2bUvo6Cjc2o+1Bb0O/4NnZMZsB7KoKN6SolvO4oEk5eULTCnKsqJPnt+
EtLPCSvN5S9oF8up3xgUpz1mSgziAUUCjxPY8bM8g5sNRcgI9p6G6Z8lSC+iZrcpEWUYHeIK7757
ZUwWPgEKzNP0SJvA7bLUG42yzDphZ+ttLf5C9xyD3LkjimYfDOj4ebXLik7UvyolMqJmWXq4gkr3
zgyrEqZxIsbWZh8oHVP68vw9xWY+8sTXiz/u53xVp597+/AvfQAe77nvv08uiiT4Riyprzh3NC42
hObLJt86heyqPYLOA+Cu6SuYhDia5/CyZYuyGjRkhnrxEAxapMQzAkUET9od6M1XkZruurKdjpvJ
UC03JNAZDuznNN5MKDLPH8XvtdFei4b2OBZnJfmvsMW0wA/91rh3ZeaDyVfd+dMiCov6Wj3iglT0
xYWmbBHHsAwjDLeOKg5cUpz5JnSTKJTuEcQxn9luLsu3JVyDIq3dt5rw5xVv3ZDsqN3o5A5eRlvg
uF7FNZ9qvy1lpaQbhF8dwZuirk5vms2SJef7UgpO4rPT/G5py3ogZvsDYly34qF1IfGPLsP1qwZX
pFC7Oy4zcMU4wxgOy+YX0NHxEaCzpBiNbttSf1/DYwBY2vrW4jpAEyG7rCFZJ1ovcKkwIXScbh//
APgQmYV/BPQk8i9GvechqZ7IeCQ9eX4QEd/XNpblXPquEdcXp7PmyiXj6dYHWMSJnp8LNkj9EM2Y
fMw/xG9xfer47Ew641tU0K51YZzMxekumOXiSaFVD+LM4r0fO1cqG2vL2zkjWiXG0yi1Gtth9G9v
IfHDXt1NzxRcXqcQnxzrftHu3eLAogBdzijIRj2BF8ChlYIbpIjL0Xz9ux1saxBByHSYcjbK6lap
/U6F3eOatWJLkVhgA5zx0Mv2DPHrUEYyHrw+kFRUMECsCD/k8OE3NPMZPOy+YxV9KNLED9iUMUm8
nyInUAi4N03y6MgUf8ifbeNGJjOOLsEjT47bO3a1F1dTWQfQLRzacvPzWujufWIIqnObTKZziAjB
sLfuf81j8boK9MNEzA186enEWN12nCtUputIILX9zo7sVaW/b4xqlk/M67XFvCS1jObj5stT+O4r
Ua7flG66QvSornQtm4txOc3XpawItt4kkcRrSxVG3KbZPz1JxLFE5Q0qPWPMEC0zE5wQ97Sifi0l
C+X/tDVfhJ6U6EpQYjGUVOcshgwhTOGbNHO4Z/k4zlhrEH0m2k0/nQBmajCBEclJkC1Y00rc3TQZ
C/RSxCdFmlj0O8R7cFek59lwWRYwHiV8DQzsn0+JAcPfC1ORUMi2Cvzig00KhHxmajeQMaz70IBm
Tk1c9yJ8TPcdj+APZ5JFVDIMdBOrPTCrMgLDBQqQy1OuDKIUNkAiDN03qOuTIXP32QPyufiUeZcv
hSGj4w5LZVwHhKier/jk/X0HBXxb864r41m2JYN23j46P6k5AXj8H7k9AnHxto4TfdXZ8S8S6UHn
tIV7A8/8XCEu+aEk5orCZ3qm39Qxde2nZrRu4TRGEKIP3qm65oNSsafvhZObEtnTcCY+b0N39NBb
Ft9P3tP7K+GTS6WWA0xUS65gUWUqEjNLGvYF9u2Sp4YdivXabxPbmNivuJ6QkBPzzUso1wyUaFFC
5+tjZMNji0J9uYNJOF5NfugKKyHWcDJJfF8b+/KB2a8GVEAe+83L1znrAjjMajlnazHn/bvy2SUe
7kEJlz+PmQHysBxTSnUxehpuy8XQW8uZKk6hVGNZJA4zmfqgjBF4CBSE4avQ+xjM5i6XQR3Jlzlr
5jNddgER46kCHofJATzliclZzLKzJS9C6Gqmz3YgP2bA+bTYRnCjxHVHMJhQt+lLWkRdNPgs6K7D
Dm7zk5BNvzd1Qa0ZJ/X585pz+H776y7wOUHoW+acPWeelwrRf/yz+JOXULnK7j6uCvCzvZROsKNl
NTmG37ajNw6q9iOR3mvlSrvRx8j4Ft7Ca4+8lXJPtwgmScF9o9trRZvKuyBMwn+yAWWPGlE4GUQ9
bsuTjmn7XnRIqGodXmZ/d6ir6Qy0oERnQXceG6t97xe5l/4ayaUFI4kzEhaB/sUcqxKNMx3+m6X3
4o06l4aBx4o2ue+OaSYYL9YjuJjcmxGSDhzk/flUq15/DaZ7XlN/bqAJn6xLXpqYm40qWcVA5+gx
4ga3259xBt1+x7ysnA4HaAbZcFZf54kNpOQ/MNbNKoBoMJMaurXeGD1jRFTWxZgJtSpaMltiffAw
faRVAAjLAXzSsIlQhahJiaUQmeliOZuu5d2UQy2AwlI8xQPx/f2xQoon60MFwut1lFBMJsDA/LH/
yXf/YXocDRFSLJZ/V0O80t0XJPKFXEwk0Ji++CAeXbjOnw/48A51E5u0hVFjcBLOwBdtqwFUFoQM
5bg5V8dYvdhDj81e/S4cBdP8yuKnVW7m5WHkYabbjkm+8+nCkzzHJOQCz3+DeE+9i0DF0C4801+T
5KX+/DQYTmMhoYumiMjl9fjQCP9fJcLfC7glau4Q9ROS2lGO676MUA3izvT9Ir7bfzIUBnS4JPzr
nJLriL/kZkm3Gi36lAFAZB37TaVKp/RDmHN68Me5aecEGNi5RusAwBAJtB805BxyCgo/9xkEjEGd
9o+K23rSNmZF/IFgynzcvh8bT/PqW9jOIUYr5UWMjMGRxqqwtpVRFckYpQILx9/ey8aQ+WNAV7/c
ezFsLq/zx8CJhw05jDZcjLYvFlpsWImk9cCmSODwmVux3HNbPOd+z9qegs/F/gae3FXqvEbisgeI
bM/IAAsDwpJdcoa3TCl024DWdAIcch9y1k3JPBDaBtoSej1pzjtNAayUwqQUYue7CbWv4njS0pZM
9ds6xAa9NLi/lhVKXwIXS1R4w5US6Vgy7Jh+v+QZdqaU61lM7JJ4nNMIgknzxgYXPFyt6LIxRO0d
p4PopWjTrHLkiBOrtSUE+L+9mSAKltQXzcq78g22aqraYK6hTn8RJcVTYnae/WIWAoGSkTS20kD1
i6ZmjwbQhzCm3LEo4Ak6oEKTI+dy2uv0d8T27W2p60Xol5Xa0e4DnkwzDIbdhuvDP83lZXEQ9V41
E6dkj/NFPB52K+CW+cnqpPmI5Fj/oVnCccanSPHu/cmK3YrSeWxTEnqoHShlj6FdRODncLmXqJWz
JBqH1ST4XBk9ATjSyFdRq4Jd92R3xNlIMzp2prIFTzJ4ZBLVlmYDyKJGVmh+TmSps+gcKorJ7Uae
EA7FEZ5hFxaa1hQeYBr4YyeU0G3HzdHzqAV8/xRjcPlwxZqz+MOZpChZ5NN6cBvWNQ+tc9AWPa3c
2v1/aGtEtDt0pDpphmaJe1bXtN+AXXTh/0gfGxW1ncFALMQ8U0W2ONhMYW3dv0LcDQnTv+V9IBg6
ztojQyU2UaflqmW4EiG3Q7NDClBiigQuyyNQ691sla62a2o756HLukYHc0gvr+H8GYBbG7mnzRpC
Q7uEiYmTdsRo0TjI6pOxKSGVw0EzizRYhvRKWQ68ZGia5Cgp9wdVHd4eahun2PS2wxrjIp1QgrSp
caq+HIyCmH9/ct93hptbqHmJacogRopTF72Mw14kl/Ju1IXk0KDPcjWDze4lhPNxWUn+XEi7U76l
GgZF/kw9KPaAPeFEZcjQ3GjIhcuCtyAvbMapqX2mg2iqTUSxXaEn3zWN/ck3xubzL4eku8kiGNS4
yj7n64W6lJ3gJRcKsHTz1AOUILlNfxbvkj4GwYWBmJKh6GgtftlLi8Tuns2y8zVu1E3rKTx0Uiip
Jyht3OUW0Nx+zBs6sltQvTSPvjtfx0pzUffMoja41VPxAAVKF+gZBm9Smkr87cxUMO6AGYhkP2uD
efuOH1j4qN+KYsZsBMRSQJPEj0hAF2RxY7fuMe0O6U0CHX0GZrpsJhPjITnEX5jLaGJs0q2zzpbf
aJHr72WJhRmD+sFZfyYOfKr6Mo6qqkHSUT2WQRbMES8BXT7eGl/fwVeS0JiCXCoQwHj1Gck4VEYi
q1AGX0EDqbOQYXpFzW6lfZR5z+8F7tGp0waLbjzcHuTLHC46wkHjsUJCY3VdJxPPWbWNYQipdgUQ
PP4CTRtb2e5UJfmH7TTTCdlu6oc2gWjIkiM50nXszqZVtm2mb3k9dvW0/fSdaHEU2QSx2shBnjP2
qcgXJQMssaEhgz7rw/OP2lk55iywI9vLwyHlixmMsH3lNPwMtfXE/RfYvrPX630g5UHtY/IEFvIw
gamD5klqlcVjtO/0biGUj38bPpfnK7cMmWK3hmavbzrGBOTVdSyFGFxzj+Eg1dv1DNd9/SE/SzAq
npmZuF29bRNjS3u8DH66CUw6Nmsiy3Q04KEXVYx200ipc0Z2iya5Wj4Ljtkxon/YkuU9E9ry9qSy
NFWyu9d/9GjajHvcwwEpvKJ/R1z4sI4XyQ49HoruTdKtO7DryJGgTGtdkm8Wqi+RTVby9nZZmPvJ
2yQEpLMHCq5w5a7xs6mS75Zqqb+8SkEDaTopWNqPo/sYipBs92eBYPwMD14Kwegt563MT4BPSq8T
XVt1PJgmpE+rrW1aMaJ3XiMPbXhzOa8Ih30LQcNqgAzXBb4o8m4Q3bTlI9jsevZcoRUiFQXZV1yN
vtyhfpriwYTFWee7ZCjfsp+7l6Q3Gu+bLhs0TROvfAFruUqxpEc/fhXhn7I9uN51yaOXsD8tFGQw
wPF1Udz2tGZ2ErOrAc0h+gq8WBhY8Qt5Dzp5wZQ8GFs8axOfo+kqDwLP3UZxIB+81DUWjyBglih0
AGwHffnKp10vZvo6d4vfYEwHFZPNgpwFavskIhBNgKc4Uf6hwdO/a8pz5dBFMyVjjs1dF10kccEL
gWpTNNqSy9fKFIv/YRP8as7hKt4OChd8/Jd0HMG8/vD+xrm3MQiaKW0O2SMhnDlCuMzjY/fjsh0K
ICwRkbpOyoelRy3GMnM8CZF3wPvMuKjORdP8u5Rbor4sWDGVh1CYroAVm35KgNjnKuMc1yhfbxDH
iD/yApSNg0DlRMYsuDVHWGtYxt4xq6P9Cqby+xpNlPbIi1RyzjxizQXaAi7K2MuZFKOWtMIdqRP5
dKlHhHCroEGOWZxLLb5X8/DzBMp1FHuiNblJQyA/9AVDxovFmy9YCLN1j4x1YEOxKWD+bj++znCY
fgfXW/N8zSrM3utC4DYCHa8Nh7EVb9/elQkuTwLDUesQKfHGeW7l6ihPEgBbVLU6SEp4H8OEglW/
ijSXSUZm7vT0PyzxbDLgISy5mYtdWa5/gQCb8GI+6zR8V5LY8hYcwe74swsk4kO2t46PnsCxbbsV
yIuWH1nRLUJIK/vgY2dlcmbLdaU+LlXQYRL3oYIrI4QIeCZasxQ6MXH+COjFnlwmTvB/+pLqN9WR
+eRwYLKK8+lmGNvGrLSz3fLPCPBrYMPGLynEwxCV0hxS7EqX8DQgiJxe9QXTrXbtCsIGMplDEWAv
cKVjvSGPGiL/QO6yi0rPB4RR8pDKPlVStiJKwugtQiLgIn+EmtXzRWHNiLPa3A2wjv0AdZugIlF8
FG+gqdqf0pxkeatGgqneJ2qMHTisikbPbjKYZdvHJqY67IEH/AKyvLC4nlk8t7I9+qC0lokDRI6Z
tfqo/1REGXttt4yRRcTRsBB3UbsVKLWxXOC7/NHBmKgyol2aNZT4iNF2GDPqXlV9oKDQ98Cj6nek
DtBfNhbc89oTn5e9fG6bBRn/M60VTx1iL6r3B2QVpKhtReWUTxBm568p6F2chqbPCRIHfU+GnxNP
wR73KSb1650bXBJsVAQJClav8G/UsJkQ8x2TrWns0CNs8o7DUk8eV8glaODV8/UmDrZA4MIk6X3c
rL2p7L92j7PX3sijjo23ODITy6uTPJj5jBcFwqdUaocys63077URfha+k8wSa8vfs8o0LxwsApnu
TmpNqg930tw8uiqLkg7rNZIdPNQOUXpk/6njknW7asCgxJLhmOOxsS0joO83H+K0d4TIqtaNIdyB
qzmG/zn5EPkUue8rAXV5pz/Mx+kmQ/lgiimYICtv46Lah2Fmx6iIDwhlyOgPiczee24mkyu9mKMt
6c7u6TANtxXuJmcLcMtYe7GPkq1xaE6kr5PHBVWmTXW7GySuKbilh2SgvtqF418eW9Gmgqrw3oLL
qgNypI0TU8hsyG3X0RhccP/CcePyqVbtskclRFUZz0YkMUvrFnWgdPwzA/tELseRfP29KOlyeWEk
Lsr7Q6tzKHtazatThC/jeJqjVoj98iiDjHlh24o89EWfnborfDkllE4lrLeR3UpzwxG6dMw6R1en
iwL6Z3LmuaP5gi5RIaC8Uh4B926dUWgoiS/iQkiLjItmfrPYxUbykK0rbfSfyA8QcfvE6MXbEjyC
plOYAYpYaSih5mj7uvmge5Vve6T2JiO6VuNeblw+p8PpZCzJot5hF7RCGrgaJz/+wrZp84AhQg8W
LVEBgSLS1ZScqG7R+2jgZIZn6GBqA0nTpj0wZtqMvjW8Y9CcveFso0TuvMAqwYXRXP4eGs4T1FQR
dke1zp2TNfh9uDuSHwidaGq8BDgEQ1WliEdkDCHEW5ZiCrcTIMB7fRZWTmPWfLAZNkEv7TJIjk0r
7eVEuE/UJIxi793vlSSFioSCcnbNbp3/kjqFOZxcBRKPo+YdZOkoJ8iQi2hWW8qop4htIuchXwID
W+cW12WfI6Lf3p/fJJ3OiOaKkpVedQ+VbAqxUrRhoeM8Qc8Mq0ikTH8Z2z275rI4IPDa/OR8VXrz
QqouvhL/3PRnsFgUrtzskdRVkN7Drcsf1YHCLyyiVOQoWO/3QiIzJBx6nWX2fuDu75aO5PPYTK4Q
wdjJnKdfbH9Nqt3bhPYfZleHxphMVs51WbQ3Ce6HFxRpZHtpvIkb14Sd4vNu8OY8EAzCbnfQDCtZ
k8v89niX+sSI7KdI2UF6GVo7CmiCnf1/C3cu7xSN1Tu/5lS5eE2oJ1kr3NmtySqBb32b83jxFvP4
p5qKH/4Uy5u0qwrCgkx21zjPYdb5LYPBRbcgZQ85i5IimIDM3dV4y9IvaYhWNDbpyKEVPslUkrnB
Y5YHVAzI4podPOcoE/xDKTBAPF2qCMRZCO4d9xnrJI5f073pqQ+yLPO3HJ3tvfuWH6pSRoCIVlRn
texIIu62Petj4y3sIlyOFqZTkfSLSyALwB2i5WqitJfE+moEHfsAF0QBkPkb/xFZPpdLjgnF5eJY
TQNGkfAfkE8xme4qI9uSO/an2YHhvtE5luHHR+nEhokSHi5GVWHG+ygcsmiTQN4f82b7vaLQUSON
+xXTAZX1U6q5t5mJPyGIzePF0v49NxNDxqo+T/fMxPIxvuu6m1UwZb5A37Iok0t2Hn5Cqv6+P78/
PObb7LXNQINrTfDFxtPJxhbLbDQKOf1T5A4lb3GHmNnivnKDTQA6zOFcX5ZBQ9YGq9IwZJ3ynDuW
OZ0b+vm/xTm3G2AKUXivlJUCsPkbEfql/zddtwqceTbpgn8lQOowBKxT/bCOx7ZnaLHDCr0M7fke
X3F9ML8/c9ciHrhLihNJnPHTGDDLI6o7IKdv4li9NyZYLP5viKlMXm2PUtn/UMWYz92AIgo6ofyM
S2d8N07uv/HKQiQnwR933a80QW426gbG0+DHkXHOZxgoN9vfV6cjjeCcCjrEBRArcAa74Dpa628m
85d+2KQHMT0UzLRsCHOD8DnZ+Z/9KuFfo4vzJxmM+CvdnJzJCOzVDXHDg4PSjfJIvXCObiP8d7cr
rgJBH9RIhcSiVgc0DnIx9bihDJRP3EVRecZVZFj3NK1iduEyD6IHFfytsrzTI0ibeexFdrX+tYD2
OfuNWebrb6yMZkK3JtxLmYshfiMznKY993ItCpQ/zH4qjyzjC8H7GTH8WIZ2tTzCINWKD5He9n5V
p0d1Ql9FdZD4aIjCNVj7YVq4Bc8/q00j6mnu2XyvlhAsOOkU77cno71jWyJUF6dp0IPRxxro5Hu/
BRC2Fqagd9cT5Lw73rh2CfXu0ETg3ndoNCc+9DKhBt0t++BG5T0q4qQLI7WEKglNUrMuviMnL/va
YiiWhOrpA8JPbvu3nFGkM+V46wHzv9bNWos2vIY1N37C4wJzOmBrinyqeiAjq6o8j1O486VSyunA
prELqbDk8b8vm9Ntxk55cUdgeWcYtQZmPLzEYLW6a8d+yCPb/hpRWrKC9hV8ktBrnTDHnYKm1dCE
20kHrxFKfvScNFLMePKB0emIE9EXc3kz4LjdTLxdsMmerPmAo/ZxwkixuiBROAJxgLqEnVeAj2Sf
lMN7yS2UhTmT0+t7JIiFWNWapc3ldTXJZekP4UIozd7JcdokK/AN8RGZZLEoMbSXNEXZOWDfE958
Ej9AC0FSJlyB4iu+sgY7/Gy135IazGnoKFACHXToj4hQeGqN+vm6t8IlFbXDqE4/05j1iWNkz33j
6fCPFXXuPTL0cxITh/8+jVVu1/MBDCV3Qym0Yr/E6349y9NPbDBeoJwOUUMWqF8C6fWMtgse9nRn
2ZeVu3yYUEAmY+OLpoOJK1DhCTs/QTCpEurY28Yex91laXp/lOXJ+FmsU/ihYFNBb6WJIthMKgpR
tsz6tFfkiPyqGm+xer9Q7k5o0kyjyHjkCJIsg6HwA0cpJN88Y6/McZ3sSMDnHHu38pRF9ZWWqazN
XCF4Kylt32A0BMECrPsUGSbvpwa2LCyXXYECIdingt4tqhT258pknqGu9en/ws/OpgH9eM5p7442
3V4JrwWfQJiM08XI5trHxLfkr2rLUp8zNWd0F+Kryg5WSXAyJNUuriB9PZ823gAG4W2Zea0gsbgO
4slNEI6fsKCuR/r0V23jxXYHgHeV3kzyBfvYSVtaUMes7t4qcx6VcnPhk8Nuihr47PSbP8ZujQZ1
VboHmSujI/RL7QnqgG+MDlfpzov1rHY5jgsxmquhBok+azzUO6DuXl+ePhkxKMjwgyyRj3Fko6DC
//O4wnTIiiijW17/gI764Sb1qJyPIcx6Z85LcD16/AF/XMymiCh+oufhVZ11cQ421lAFf4Dxwm+m
UceHIQT/Bm/8ExTJh6GH7RvME+0uoIr6z4ryAtEmdQ+FGnCwVXsPo+WpjpNwvfK+DXHGxeRs29Tf
a8Gs73tg1Laf8AYz38gD2HrsIjpsYBnsCbmFebPjN3aZJv7q+yA7mCW+BAYx5fb/IsXYGMSRaPUg
MSRMIPLJ8Ck/86TQjyhLrchh2S7uTzfjvRi1fJThC52KErcUnosuTUQqdRfti6d5XpYx9jpCjLLP
03roEVigfkRvghOvIi8iwlyLDunGk3x/Yp54K4IM10fS2Gqj+CZGNfQlnRjgydGFoWai2MULJaiu
XZJ+8VdHMW4etQArTmSE8TAdbSD94RvaQkaqHOmUx60+5zwuzft7QL4TJq6K0n+W6pN0C0Stxm0j
rMqafzPyBjMIVXjez+zekH/Yzu6a+R2Rt12AZCP8a/JDT+NoTxXwDnQ+C8o4mT3RT29lZlrOqtun
5x2U+dqJQfchJLr7Ioi8Khh4PphKOGkI8z8u54C4hYEq1hN8eTGViOk9pdnLrYmZ1MhGGAztYJo0
f0Jx7g/Zwu4xmCrwLLHk/c7mL+5WbWtB2pxMxmrJjsve2uUNvf1Gf3wpi02cacWxqjscF1UHeI+T
P/7kknjs3WrFtUn2kmn/4B3hxY+ZcplXQpACv8yGYkSFPB30wTe4Z/0rGeKXatzk9Y/XRoJgn8Wh
Xc+laQ6d97uhgZ064YGMCLzqQgHEmj0Ur/xGUSoaioC+PT8lI0+vcunCWfAetZHRShS0wczgFdSZ
BHNevc+wE0pQBdrZDtfcSL1As6t102q/lFIU0szYlnvhs6svDb1aRAj7NIMdQ47xLlie/oBpMD/Y
SdOm1zqCjUPXRlvzINY1/Oo4idwQlAewSloDd4XdESToO+CFXYj2OSa6vmqEo08EFQ6p8C7kWxQK
3MnPV7aDLkEagxk0VJctrxeqcZ95caqguxPPMFFbrc8TnII+erktIUN4vlkVvphFkrJjfwInt4RU
DwmFFK3+O/RBu7XZ14jqy1ireNzTI6dbhJOvGbWrS1IACqAEuc8a0O9PdcXulkJvUrzo2SwYFAW6
uePFOrcICmzZ/NTmVypkKAIxhPl/CrskpDBLreu735Ge5Fa4Q7k7pBT2avDnLfjW7sl7ArOdDMB+
3MA0l1NVZXr70nEi1Fes8IbW5M4w3pvqN4hLG2LXX3kxyUBbOOJJ3omLloGVIVHw0ohbRr1jDg76
5HhZ+/BjLH4YxJjPKO7i2xAuRtk14iWkjgqF3jAoHem2zFc5teWGTD2dPufmHhNUJZN7WwFp2AdK
nNfZO545cKRJaobpeT7AOo4CZp68hhxmxC+xnbOgr0qasVjQGncx+dMipUVlYJoCrr3ZSpPHpHsK
1wWzxMHMv3bimDx6jjRWfgu4JG4RNWuDs1uwJt7cU1GGdYxgvnFVXDN4ZjHBhkfqQzlkvPSYXrx1
Z2hqqrovv/B6NKx2x4YL0CdGWzNGX4Y9gpzAv7qPB2otXbpYhMqSAN4YtPIFkBYaOXh36xcmnV9k
do2NLi88fOkt7oIi9hPKDEl+87hGXc/YwLBs4I/pJg8cxYxMOLs3cqtTn0rPO5FvjvwXhho4bE8B
DvV81l9Ufmb9mF6Ogi06AYZRULwIA36yJTTQDjhVaJ6a1updfpA/5hqWv6qU+Gd2r2MFc4ilAyWl
SDsjFUXEV38Pxol1rZOt39cUM6kPJb6sCfhn3DcbVJT6fSl6RCWVxMA0DmS30oabV0FE8tJGUffb
vf0doepT9l12pAcMZ/pXjx1wyPevfRwW1CXZLji28m4HWeg+hC5EWO7gm6J0WOjGdkICSWFov1Fc
CfoekIlGCnMJ5sDBJV2TrKd9iwBGyRR+ZIN6jFIler1o1n/UyFrU/fz+B7SJ1WpmnE+XRH54kfVf
gpPYRSoPh588/ClT1ckqRI63j12y1TYqrGF8o9uKgGm0QNOmKjODPioBPeo7kX9Rw7RLrAUjdt1S
ME5CXk1zxx581NsBoqhhBBdxsNtLYrsWgoC0wp0vr4TliL6XD/zqjcwFdAVn485PbDkFnY+oZUSF
UptA2VWU46LYDZKgMoah5vNG201D5tIGCIBD1X1koa3Yei3JS6ZY7mrYxriZug0cXo6tf0SzL4SZ
jJPLKbS0NQQHdAuo7h31hZA11bTuID//1QdhZ5enALiuBwPCa8UUQmBAbAoDXjTj4knfl1Y5wE/c
l7+JlL0sO5W5OpDoCNkihRpuewl7P7hyrNjH8g/zvsG4El+LAGKMNsUbv+2i5crY02rrzQcvLE0q
2JtEoEiS3sS50Ra7uc5voGVKgeb5nsuk5+9sf2uYp29GI1FveJpSV8GsKXlm2w+MF6lGS6ZkUBmH
QYTKSd+3Nw/kzuAXvi88PnZdc54QVnXcJNVBgK3oWtQ1qbvY1ArEXzOYruok9G05Z9wm+oIEDwzk
WLL4/r+z9Ltbi/DOiiyVxWgVzKvXST10kKmgucI0qm8BQ90b3811UHscAd75GHh81CH7UPknrMVh
vfWxJzoyJ9UAX+pWqBSpVHsZtqCfEd/qZu2uityRZCRAUVW3RLTrnE2jCnA5tU2YiTmtdYCNfomd
6vYNr/+zp9NU3R+w17n2EuLqrHUDwnHhfsVsZ0QWljjrTw9Sv39VgDwRZmlpi/e8uIXpEo5JW3jD
UOgOAYGe3phZzqqswPzz9vhuRnTCzRVcTPGnXw08Qb0xpuZoP9ZK/TvfDQJCZlxclD+KeQTthl1I
YI/3Kf0QyqYBuAoss2vtjsfjuV4BORDgOjYPqlcALXwM/5aQ7GhLY3Eq2tSSyBo1FvnsI6UUDH7c
gIjvr9MAxtyMLRo2tnwSYJPhwCLAls33g4jAl76QgX8wwW5kFAGWz6bFxruEidV0l4PnV2C/BmFT
xtyHkhOQZpcSHXzh8q/ZP9HB0DxLujhMcxfMa63iycqQRapP+9xSSPNCoGjMnwyJvP+UAWqZXBjH
6d1G1YF6Y+x2gPYUBfpHsF6k7ybdf3AkBPxx5CpZWcGsIkFwsppQduaFNGODBBCQLUf3D1vzxBJr
wa4/Y/NxqeFfoTDS+vYF+71d4MIYHQoDQuQOvud08Xao85ZpHTFn+sWJCjzdxWt6PzKRX4YRPQBr
oE7ANG4TdMS3j0vLcf1i7TZWUxvXhB0vw6Pp460K0HzsEHgF8+1w8sCo7ltlFB5e3Hanf06Q4TGb
qB+6twLJhrjT/EP3R0jKTAPFhyE5BvVon0tPucuRLupMdDECzwdQPDG4lsp/uQEQo498n7Qx0Fmr
Abyu2R0zaT6TjdweSlvMEFqPlGywiZA+mwjfOItqM0tx+bC02SeQPFf1FFiPguvJb2P6wsoub1lc
JTgMEbQj40dJNsW6S29PyErhz2hWicRw1y0JOmkuolEjf1jfyB7jTQyIEAVPFG0Fmf2Nx7a3CIqB
awnknDqhxzjFicbNBUhuKwJd83tpCvaYJiRZoB6lhSczk/YUAHUqmml7Sh0maDpDAQUYKJsOi5dP
qf++RX/vSt3NT53QfkggIiR/lkL9yc9mHzeGodAKHp+CWPmXa2m83CpmxtMC3U3FhBF65C5ldMqn
DveM3NHSrtjUC53wJaGbZ3QFwrU8/AvjLjEDTWsRj+l5og1vDYxm8wpbd/hU9qH/2UsCMOWjgseK
CQd15gXp6WtF1H2WH/I+nDyVIAJ6HDdZbXzz3BMmmD3q8Rk7n098Kkg9hvc9MHXu5z7yKKTfW5ZN
p++bsNY21FAi3IxXed0yRR5Os62jxQXU4X9TwdrmhAFsgmr/IO9T0eoZKfdjF0EtK2cGLVtRbv5s
q25VUbC5XhBlv62rdjQbRRgp5hWAZAbrhTtjQTqSyfL3P3mYm3G/qxBroAWaaE9uEeWcnwjWnwai
LmL0InFNsUZFOTPrhuCgz84dAvtzb5g6FAh67IFN9Kaz0L1hY0tJMg115Fj9QYTliuNlYJvhAMho
Gzyt+IQ3M4tlBCcI36406qPh78IAlzIdO5vbbQ+jVjHigxTYlOz67uz0pG+JK9LXczDodRiJostR
1qVSH/hydMnGUNwje5ndjOSb2pR1f1pUq19cyvF1ZfXGlMZlQ5ALdFcAdM/AKkVvZP7/sBm4npMX
fJTuXVM56Kwn1sN7U7t4i1lnSgu1/BfgePrtdNZr0yDTZe9OrzKUG+OvnPHx/65XOo0sPuiCr5rX
1iwYIFON6JnwzAvogYaUPtBIMyB8iESz1Nwo4unf1H1LSmttF6DE9qZHc8wMR7TlTcrlyTJ8sN0/
zZCIh/jICuE5hf2b7ySVIJJGuveAZh/IyPp1T54rQ4SXymiOlehUt0TS50BYDZxOv7f68HF5jYaq
ZajLGXE7BTvF+B1ffdKXqQ/XlzwVFrfy2G3/6eM4jlqR+lMU5ZMaKNlo3daynMUu0GcZeiCrnQo3
TXGoYzgimkn/VkAna0/xm455aH6iHrTY2tQQkgGycFaPIrQNAOin6L6eZf0Rl0SadUf3G7RqKU2C
WbvrdkGcO9Acr/Zs0Stb6VzFAQQsvQNpBGIFzKMlef0JotcA2Zg/a5Lk0/13qBOwLC+8DpZ4cyvP
LZD9nemM9FGvlkSZ+nlMVdAvLTE58ZrHtsnO5sKfvkBh7ZK3hxELhB0CW6QHYqvb/uS4971ADlVS
W8GZpOcxa7hd1hrffhKzvKLkl/8TRQXuUmiWqRrMXpGEos6UpT7MOViI/M7onNqFz+zwMYS/rocB
9CzcfF2fyWLi29LuBJm8W8TklZNxHdnUDPk+3+njqsao55GEtbrrA22G2o8nfz0aBii94MxOLNCw
kGnfVBa89J4e5YfpJUwj64sx6L+Tpjvs6wymqLLweHjDIfXuMy7A6xHUMmoBFsghqJqpGIUG/O4u
nTeRhDtMqcPbA6pbmt3GZpBRSk4Z6BJshaFQIvuJN4wd3SsWAnFFhIC35aJyJhDNrk2zRPR/Wn6A
j0XT3JqO6ZRubmO0FVjrJMa+f+/x/cUkp/P0dCYOGF4ThkEFzTVoe0f14UXM5pyp348pRPE8C+lO
qn98Ldqux54ma2Lqr7KJ6MJsKfBad8MmbZTynRFJDEcsrDrigtQ1O7wFz5ktNfJMcd1pP+iMOviG
/ZNlQ0QHobKNHzSdjtpBB0dwAPIlHWEt92mgkpGcUpcStiSjscugrYhj4rf75uDHpdzRAO2dOW/e
Qnr5vGDtCpcuo2qPflXjFntbf6Jp8my308wWdeRqxwEy8LCtoAWV9uhSWJX492nRf3JvU+a94ULU
uUV2RBBTQz7SG4L5F/FkYjy/ZExN3GO09I5abVkaibPQyx6Qi2G0Rp2UngJRm3GrC/8XTLdLdPRE
mAE1PQEC65Zo5bqpQnujueGoLlcyWagiTnO0G6zee3bHPcrKnlHcV1E7D8MtX//3dRZUPupg/+J5
zBxDiUtFxdjGMneRNZmCR/UsPhQypHMb6qWYR2McMNN4x9HBlwSgkSMwODJC6+cr1vbw5ETUlJLD
jIFz1kPWXz7bvNrsZ9fNrn2pLKLUgNtUmJIK3pFN7g+eI5QTFIEWn0SOGsunJyH943Tia904zGD4
1vGL42o85Oud5FCwinfOj+oeGQfZTSRUXuNtMljwQYuKSWhZKOPxFKD6LgHi2TxPJkogsno3ipiw
uH7h03Hi00EfYq9bktQuN3d8wmzdQinJGReTA+bwBDRTGXHpiyWcLAkzK3lZoZ0zQoktbE8K6Fhw
JzuEocMxGPvPvoHIB9pagzCNGcN74axcmXwnzu5428jAFPw++bi3LJGn9F8hSAnH32VPwJ1B1Dub
mLSLBnCYZWsgJALPy6rfyqBkPRyWCKue9bkncMXsyYbVj5ds1KVBKUijkGRz/jJ3PebaVV71Xczv
nT1FwqaWlg9onGm/ZunFm+BI4oqlW98b8rM26hCFM6nTf8aY4qnVkTpwHKwvTlX55k3BTvzH5GJn
n3xnevAPpJq9D4JeCHZmzjDgYJvNrCuHSbpjO3vbdsAXTPeZv8SMtvnOhxnVNC+Udv+z2ba0GO9d
4aQdeWdjFxPg2XvWxeCjzW23e3jcV7mKVtf46C9RbgCJBnQ5lbMkk0/pkgiVLrCXzJi8DxX10MMn
r5iBkXgXIb+gy2dtQPLr63+3xt4SR8rdW/aQ8Wrm7mo30AqECRXTj8c7OUl4ebgrwM1QdpIh17t6
kIGO+hkEHFUrbw8/Qm2E3rFx814fpbeXU5vFNQgW4DGtzHhJjBcvvEkcYLw9bjvpfiaZLcYDzseo
s0HfCG2ZGk/xtQkhecajfsvEteoFRt42yjpe8TFUQs8WZR1CvrJmEoIlALvTI93UmXZtHYnrKnkb
EQV3Oz93eayDUl2KxZkClbhLJooSf/0HNnNoBcnrtcp5xmW4i7v3hNfdW+N/v1cWKs8ybfwphZ7S
cToc7N9Y++6cUG0d+AVhUXibmJEkHsbBR49oXZtLabugKIgqxkWNxKYqHj55peBto1whp2ytCjNt
SNewHhAfKtDZR4RtO8TJ6ONVtSNuOTUiibghUF1fIpd0iViObrp1462rz+bftLIHE/oUF20mv2Mo
cmqviN0LXFEefY0i7Kd0IJ3hA6/kWloES08G4QnFDmIbC4uXWucuxMdXu+6lFYMluXxspPmO27NO
0MKRDw8E90upvUGdS9wHZcQaCxjYWIl6G8Za/SZJFLWNi5gzK4fBOBDcJU+MOIr7igckdFxv3CQp
QK5+V3xqBsFiRZJYZjYcSZjoJ/O1vT7vc97P1idK8xff94vNdXOZ1k0UZqZF7iJEbtAcARHh9Ts4
IgLC14FHuOQmPLTIpd+qMlVkziI0NMhLJ5Al7xJusOhNtn8mBZaKE9Myf3P5NKZ5J1L8E8dVC8lf
YBfIBMgD2hEXuikMPwm68pzdInCCVa/dd9SkebLHyGzikH2zSSjJolGdbsIIA832J/h7WyOpAA6s
VQ/ENFvBiecAkSq8m1x0AcRDDMCrmYPciPNNwuopFdmnG8Gv0OmThVpDXP2ALK08ja1H/nqHFzLX
hBb07mIMZGngzr36SK3gceav+S+Ed954KVC1326NJ27aP4B27RY6jlk/Io6zp5eb+9h4t6WjYMvm
iDyfGLRUtGaZNILj0Yopq8jCmoc7lv1B/1/kgkkUFk7pYv7Fw5jySfbaXLgcP+lrWzAYWEVW94O6
f44p+sjGQ9kXluvx5IGuLbA33/WM4p0zygizGwM+2BKK23LMlw8p1cQ9BhRJ+korfR1mCf90+Adz
M4EHknk3zq29zAsJIssgssleREm/4TZ5jt3TqNUkiu8ApmvIBeSBkr5BKc6uAiokWE0+DhH89jdi
KKFE3AVCj40ZFriatKVUgotuWk61f6ydf15kxJMhpFQtEGt1phUexQEOvrwZqdcOZieMPb26XTTa
zipKw1Ys73X4V/g+JGatCGd1u3cvsL4mSB3BhN0Jq9Dmy0RaJws61518GOoYoxKLJBWuKsIeK1yj
FOWyOHiUUcu7cVBo9repdn2FoUvTub2pLa4cZugHnFznpP03WZujmhPV0wp5CvNJDnjdM0DDVuEp
bCIqnzPXnUeplW5jg4VhuiFG/Ey3dY14BN2IE3ch/QohPPc7TJI/uH7lbhuf6ap+oiuded5zeMMz
9PrcpQ/CG4lW57wMAkEs+CImdnLioWQ/eoLx+rcDT+iRsUJOmYegG8+16Hc/4jqQZFHLdeiB2jn/
/vH4fEp1TtRgid5MzwQYs5Yi8n0wFTlEJoBW20oZEWfe+YC7Rt1R3bCPyKU7zYvVodZkhELzo3ra
rw62Qasdr7CQ4NfgXfqRN51bntN1SiybTu8DAVtXDd7/oxQn3cbzNs+DBzJTsJmllwP8HPnSQDGE
FteydUXox8s9Jnc0Ck0jZ5Ph/K++j1fX2H6xDmUlo3Wd9w/kdBsD+2jHy2VVppROe5s1zksbkngV
4qlD7e5dYLeHVD8rH1Dx2B/xpm6CM+9MscJRJ5m/C/WN3Vd5zoFWoEMiS+tlC4iqOtfDm6eZuzm9
zprBTVmFIHitBUlThzTDrG8oqUQe9B/rG6C6ey98iLQwcifccbuEQ2gA4ncAVmZUubsf1SxmHEDZ
IszhyiLhZjQ7jj7dekd679UuxAmoGdmASJ06h+2IlLRvBLaRVy9g5ox6wfJqiD2yTI4BT/jmkOwh
d8hxFZoA+0QywKiscR/OvqA5BPIQ6RLSz5+/IRWIrRKmOq7P5AV/8tOcpzJ6x+X8sN87grmY1/9D
Wm4Dtk8+hmJpU7dPrLvLwcM0tVAvh1GxNxlYjIQJl97FDUwxb3lTAJln5TvRPxEDcFFnACx9qWum
0KFEpAqNuK2IVIcc0SvgQiUXB5P4DumRMj61/BmyvPy0wn736XWvoMe+RoKYuO89n4xiskjYtTih
dQle4XofzE6KnAQGASGhT3xI8p6xZJrKAiMI8TIe6hgp+4uY88JrMHjTs30dgXf+Ir+jmc/rWpF8
hxOn3y3ecwTtU1Ui6Dx+dE+Vep7oIfb9lIuZXKbrqDiDI1FiRqmJapEmA0vYCXtWxXQYXJmXDw8z
JsFF5mmna4EEBZSQVw3xJsLdHg7hy9HpBptoObYDfquuvv0M7KB66bwPewLCNynRNJEpMjP03laR
jr9Qa1t0+3EmFKFQL/U9D2w8loEuLzByBMQhxS8Qb+p4N7DfQWtQFhJisk/Epf/XwcC2gJ2JF4Z8
RtFLPnt6D/Gk+muwCKiSqYp5UIfazT++z+OfgDzlWHcoDdlMaTd6DkD28TNCYFLO8y9g3v/cABDl
F2knJLpeycIIKkPaL3h8KNSmAbaIf2YmsEDoSkql+s32sK41sk1pkv7ldWV76qGXmB0tvLvL9Y2P
C3B0eBvdWQxSzuMyPAyJ5UxiC18AsL1SuSUK5b73ZdzO2v3qQMjOTjvvg1AVw6RcO4SXz7ABw9ub
r0ESbAOHNM9Wzx9LHL5/b/P3yOT6glXS5QXrO1wwM9rYP8egwwNtdxdV3/3xAhhcCet8dH1wLtiz
K2t4O0m9JCLhUNbbB1UA32yoxkNsXHYBX3Xj6Rweqhmhxi11Im5DpBJIcUvrIeoQy0NpPtesy9ul
8v4tmjdYWcewrwjwuriPk3Jp5Uk4uHGaNCBqJZqjwnKMw7LXpTfCaJgloZW47Xsxs20Is9KCPIOt
DyVuXG/53Sc8KPtAicEo4Q1QqZ7/lu1DfGbzssigfa2NBqs+kBXs0ZvBGqZ74UjCAYxZJ4foEINQ
RKvOXCyyImq25eHqpL88HLuq7YB2pR+USSA/NfRtViBg6fFb0kxKNdD2mO/DE357010P720Qclzv
zqeZFBmljl013/78XsaObJR+VHYJ170BRJKLvhZkA4RtNTi8A3aLiSfNFav+1fK48wbXAhq/fXlg
P/w7pvGSa9JPacLgi1ZAwPYWlUDFB8nxD0i82GUQDKTQV/pwiEHyJnyEWLDrO2u3KkwVsVy+tR2B
GQQgQLH5HBSqiOF4OiKqmpZfiZpnIxyfgakneCJvPNU8lUC8iLQwEw7JKJwCPz/viC4Tam5//HeV
54Y/1iHz6t9Tr+j8iU25usEmR5ddZoNSfaOU7rd4AhjUzgNCdpCh4/Ht1WUQXwtfRIpdZZw/gRdL
N0JxAo4AP587yKLuX39JVrr2sb+YPFzw/obw/PcdIQTEK1BG5seHkS6SV0lW45seC3YauUlJkF2B
RETmeFe9InW8x6Lvp7Ux7XyX5+atLtdxh6jmoDwdDGCHdusQnyPuHrJrQ4Fj2n08H6SYNXSJk/mK
EOnbLmd6j/5/BDJm0dFJ+SYzSsZu6YKuzJPPqw02J9HtKhkhjpfOw4wlRL69L1/469vaXnOuREVD
LJNke6r0nRbOVuNjUvAqievnx0GoiHVSzQ5FQDk12U2qzP8enQdv+Qb4jAG6AVlWJhxLShXL6Ldb
NVTmojd/sBcxCUUjnip0mEMT/enD/csvHMGfX42Jbh62C7+43M+qOzT4m0wYuM4CuoTmg++Vb6kk
zy24ppsY2LpD2I+PjB0yTFD1VdVnNUPiiQfG6/66aB8oQ/W4XXaxY00/ZbdhxqRaOf2xIsEiAykl
L1GjzEffrwPFZq2iE3pXvXcY9VgEwAxPIUHvHf8ymG5KFQaFFZcnNsJxHk9a3Qvwpjtdcy2GH6Zt
ciipG7eE7OZAU4aGkMzirtcF+2evc96uLoVNQ/mOxGrPa1FNFb8qnHftuJZ8AHklyR9xjZXsJCCE
Ma+dVqvbD06Vl2U7QIkyKRqoi4n3eSnCVZxaiC3v6IrdTpGsYuJk7+v5jEKAXPoekF4q/CMYKdR7
bFXe8SQXDQsC9FT4Qxsqf/mN4pVSJ6Oh9rP/lZwAJRv7/YfPEmciHtIGgFi2b4jVXymxSCVAQ9Sw
PZ5VoOUpu4p4yLqrDM2r4a2iXZF2u4hpvw84pO+rNNIXaskONX3GeUKkhr7Y/05ZG4Uj8QkAcuT7
pmPuxwXvEA1RVGWBlP5IKl5BjIfml68WfpD8tsnHCb6tsPdJzLYVGf9R8b7sXVs6486hMexVFSjy
IvSoIEtLyuJY11rsdEj+18Bf4+tY5du0tEP7bTCV/uMaft3hA/WEEdmD1ceUy5NVopBbDBlR9gE4
8xQbMvFf/LPUIlFpgRm6HZXgeecQm5cjvAWzQ3fPYm5M6pZDU8O2Eb9TUUO0HWxn0KMizus554b/
1+kbPjEz9/OzBtRCEXRmQ7O7ZqmNkO5AHJoVnFVykhHkDIu5jP4ch2Swqxg104LubLBg2t580cXD
os/GBh5GF8wnHtJuAT8DJ1ymdI1HiYJPyX8EIoWUG/74Pq4+aqFMJsDSHrRUQfSDc+ZmXY8cJ9I/
HZ0BCsBiYM7FL9a+g04savI26q5qJGSX73Db9XWykXIRyHfDDwmkX3IHTaKXW+CUdMTDXVSUxG7N
W1H9W0Y5CyfiSQaXae+7a/ylsFNIlcWKaKA0cYDdDxW8oJaaeZRowttjva0VisjZRiQ1KIqEYn83
QNxC7UC1XY64DIxEN+xcco5hDDdnKK7fRGCuOOAk+iNZWJcA3wajeJp1sDxeZB5NLjj4Qs1dfyjP
krroSI1JZ+wfEYSEklTQa/efsWPKrY7VgAnaki+3jJAffpc8SlQVhH59iXn6TBAqySwvBYiehGSA
j4iIHUAYnwYOzIu3xwhg6ujguZ8iiJHqY2g2lydGerghpOn85t0OoP6q1dhN1yiKG0FGIRW8Z0J8
vwc63iXsNh+qjl5H33ScffHO+CjGWEpRc3SBB8pCW+5XlMDiOuOLu2jq41yC0dpnv2ZljoCkeHNw
mHWFUL2aGZSRVT9eaGyeR2WGCPLIRTOfhV/0uC4sV1/fYPIetuxyQ8aEoOnaVd4HLDtsijyCPcnx
XQbE5xOvxqDEp4ZFBs3cpDzI0wU1+LWDbGp2oj9nrQm53TMcE9AzwewKBcbb2ge4MxWynzrhWCGj
GIuDkD7kaBxZIvDAJqk01+5LM+jK3G/Hb8obv786oLxTYC8oF55skfFXSoF+a/X806ZEGJeizcDE
Efx464SSU141D1lRjD1ujNOieLvG+bT6yz8V3ctSdBlfsWxqtc+MmXXg6omr0vfGqzlPyXDQu+0F
7p7CjdkeOBn+CYJNRhyYWPgjCgk0BL4Dd5PDY0ck5q4M/Vr1Wj6wykQuP7KYTDUq66ywogsv9CVJ
Hsoc3uQm5PTP1cTaFWOsp3MYgHU+OEKj+NP9w2GMZnrczjRSANSeceowD2KVVRmSN9ua+T2hIFPT
7qgGKAeHJMot6uEvwxbbtfOh0XbGq9SO4d5bEW1Tv7tBnmn58uOUi+vCVGSWubfXR8hGB5HxeboV
ILzv43CTpzlT9063IWIbVQfX15vbypkTfSN9Q1CpDKRwGNpQCU7b5ZH+iILNBYxowHH9j3+IoL+8
mTCkTB69Op4oTaC3BUcKTVxdyY75LGtKEP45DR9Cp47t4Y6FA5TshviyFLikJJnkqmMu/qRbtS+Z
3wI4bL+Tk3e40TJWHTNQ4Um8camQxm+XXbYmGmHCk9F7PnBm1QJE761GZmchRnQHKO469iKIWl+L
UBU1HqXtk+GB9t2MYJZZ4vGgJpUr05uShEdkUr+957+GBnoKi63I3oOlCsy+gEJjywQ2PrZuQifd
Bw0hiL94INyUjG0+XdqFRJdeiNsP3oYSOz1XybtZ2bx+Tc0vV5eq+qM5l3P3EEHvlprjOvgKjsa9
fFxguSIwIydeQkrWp+hIfhlTAFVAG70ncQF6X/I7onYlUF6jgSYUntMKmw67i2+F7sKc2vbfTFdq
xxB9wnnmIg8nAunU+T7pQiaGn1SWlPKOPF7eajJxOOHLB5m6yDSF0G3nL17kAuFIKG+PKNBEQAhZ
vtFpcDAMQI0TqAj40bvKRnXC5o+xwTYLAFQKhadIFmuscRHDiNJYdms6PFD1cwnrqmuvswsGBVPB
KuIAVbysPUqGl4d0g1d8L0Ih3rP8DR3Ik+pnDfgP+qfA38WrMbe1HgVbRp1rkR6JMrUuBoJEkM6f
UIzoqch6BFeaz7wItUCa+4Mj9kVdwGqkgVRCk2urIHXcAxOd5jkOXykifcEvMim1PzP7hmgUmLPX
gEEcoGCtcAubVMcHGXC9Ug5/WyDTtfMyNfqqp0tAhtJ2ZSdVhQ5BimAdHGxDb5G+ZhwJsVuslOzZ
LP+9gAnWzh0ZYRsTRo389tnn6zgwTC2viVr12heYO+WnBc9Wo+eBM3IZkXnNjublMWdv6jZbOAN7
M+xWkHTrmjpwt9SK2jN+ona2xH/nAR/jeX11xzLiqijIy+hc9rmFvXJDJOqMAVvHah16odM3VvDt
p++qOTKVVN1Yw+1ju/4XbJ1l1S5N30DmD/picXiaBMUWRNW3EtAAlhKnuJ1SUFhy4t3EnDBFO73l
GJa/7hPfaTMjxWhiKcgDdmBpbbQCDVduJXPAZ9HftLPmdh57KEwLAfppY1lnigvf1Yd2Kn2pExLb
lsYIgm7ZfNk1RAL+pJt0M2kq9MqYIzyx3A49UsSdnjR+6012cOWwARTGoRIumayzuVuk3PJsgBYd
b8Msl1sdA59APz03bKX8Omr5oncsgSD/sRnSn1t+fFUI8Z/66MrTNhfY6mRW2T1tGz4sB6JeCABw
QJgc7/ZwIC8AYgLcWO4cwrzSKlPgv9+/SDF+8VCtLm2c2LKCjRlPzRuBoZlYwsunpkLSoHAGBBk+
/Fgy9ftPWkcT7AYAN9/eN+Wxa2itX7mB7mrqyY75GOrkyODjfA+tk/53521Ppo16C1u3JZ+0xTAz
Xebns6GhsqdrzutA6pwWbTtSYHRT0GJCsBrxXdQmKv3PO1srca0NUPrsDIXVJYD9vl6vVqu4RhaA
esLxUO0OICrjLD0lffboCALOPHXA4xjMpiTOZ6aVrvSg8XNHKowczqnMRQ62DUrksKi1RKWfclJB
+ZrdV6GiFCECuC/gI4S3UwZUSjs5p3c1K7D+vgtwa4wmSz4KAyOwWjBsed81iLXc9SChw9u6JQzf
aPAH6o3Wn6i1cgzWj04PCqJ6KYI7oo5NLD58kPg9kr+kD9yxNpGvy/4/dkqtO7GZAwK5QiKrtdgO
5czakzxlxYCd5LzpJclh5xb0g9Fq3vWBd0PUp10OFBlnRveSMHJJ8l7gXxHJzPoTrmss2zEI8wJY
itzlk5I2m/ET0dnKpEuVmHqkWE/zIKDW9FT60aLSLKjMypOndHucqPuug7FgYpYXF+0pl0hD5lCS
xVQKuW0nz0aYchMnfhAn84QiklgdfwX1ds690DkvuxFEhjouR2D3SLmbf0jplqLYt1zEuqDUoEvm
w4STM83y8xUys36aNa2exeqo9gLCgDMDysRR7HU6YX+Incgj29FEixy6jRiAJJjHhf7X7yP3rF42
YReUmwiCjRIsBV0cg6lwegBQ3HUNEDnBG3Fqwu8At3xchkaftMNIQnNoICJBICUxjJOicDPlyV+0
MI2VB22VRxGpKz39eMPduNqK1NnzGByKjpY3BqjE2KquBsTGBESfAqJKBaz7/3dRuQRv6daIIhBC
xXVQIm+Ngq5M5VtmtYdUCUa3WLPUiNgKEDXlLdYLPPBqgvzMSzDRsG8MDLRapY0UFlJg6lAFvUv3
q5YnSYpBhZ1ITgq/YoeoKdXJ8pUz4AjJnz7DG8S1aRJcFl11c/Oyi5XOBlZ3LrIoL2QpmoZsZqlQ
NODhFQ9JnLwN4PUnoM0ZsC2TFwuBNyde0X+jBfucHgXgAMcqBDRfVKrUQaPOIk65R55zeBprmzcR
dDnq16vn0CVe4zplyIOTmD86VLG78w+ju67VV5W9h3sbLZwqeVGFsZoP5fvNsMtrYPH+DQj/KdOs
46N/+zEV7r+3Yk0DIx2C98+nysSoEiRYC1moRrVdkHnrwV2GnUdv3o9En8KRzsSDvQwk4Da9UxLU
OxCzdixW4Y9FdyDpgKBgTbkkK+sFcv6GhvYglHp6b5T284imv7CBBgEjXUudXNUr9+krmlxtMjyE
BIwldU7+12+NFdki1137sy6wmYiNgXbVgP/YJPWSnzNZX80lAZQ3O9uI+4ZLoqPs1915MhHOUP42
2ZDRvcWqhphb6NHAbQsn5TtxcYhM181QKuO/XzOiy1R7mELbwfKTo+BbP7mchjve1jLLzDPaZUEe
6hFZCD6iHZF9km95bgg5G+7ZCdZy2YpQJn6tG8sNP3G1WPJJARk7fDWtSq0mMAcoYimY0Q5m8CPk
JWVp+HqBR35TnhoNESL7mtPbZZ+tSGE9WIZuUyhfyRheT98DUNSmUJDRQlyOhqtNpTs4l6LF9cBw
sIAnYYo3/nHaqMMNKYko9oqPyfpHvUbifPuqb1dZbPyY8plUH1PKMoczLcmuMzQGCCxV9iV4QBCu
/aYSYuDeohKwTLr9ItGxK2HgLq95COggQx2nRhmKjMeImdta+CA2X1GGh+bQvkt8Nr0BKXwnzfA8
RLOgOrrnCShmIZdIsmRWrt3EtkV6SVlbPqegmLCIk7G+7LxcWmGcT0KttVM3tB/059FDCAbetO25
x4ODcSIi8o9RJu9dMb82yIGlkVCNCO1XHyScv3qHyrwfMRdZqh/Ro8DOjNTiqcdNmYstUyGBGrc+
Fnz+HBaylL0ppfrCs2GN7AnASlWVOMtB1VjeYxbcXhvmyejoot6GPcsS78weRDc5/9EqqAE1uhrY
ApX23fRtKEt22L7CLg/Bv6+NNScg+p/Zoe6MPhfVng6X/KfgeJX6+vSr+llVavCE/wh2XKC50PCa
dF3VhYq5IYyyNqA4wkF58l+/WAE87H5qXuyXG0gWKd4FLLaJXnb4wwep5WPYY5a7+01NCPnOUYm3
Qfbkxwuj07sA9xA4AoorO9ggdB05uxoHxnr1bVHT/G+2hgWbn289CVmOlYs6IZZH1d6FLsUIfOR0
HrFlLgAZaBzAXr8PnRYvitkB9wDkXabzMyJ6oabd8a+7JmZS7jl9Rsia1zCsmA+E3jUmS8cTr2rf
DgBg4NlTFcTcaKizGJi9FprKiA8POw5AVdnueH5uhbrJaiwP1caGYvxWPz0Oe0ffng4V2xgBMgAP
+G0sOG/+XkHuJaVAxn4iTrgLeNYjOlMhZD/77EG/ZB4X8pqBUfxerZ83+oPiLO/nsTPFOBAV9GZk
7p6t1ohyad8LRUsh4YVOYC0JgJ1rJrZfmfQU/EMLhek8yDggOLr/Rwd2BPvvcyfxWRqMXoMS+LMh
gsPY316Gx2nSDljSKKZVOrWA4QnSc/XbcCs2mtsY3KCl2IeSB247Q8zbyi1w1ERLOz0JnmN4E0UV
uNYQrbWWILka25+Yp48bJBBZCeIOxMOuudRGxkWjDYpAhAdE8D/HgB25WzwOxpTKIRrlpC/JCT7V
BAlgs6e68EaOfB4hXnpJcPXTRZwgEsUWRnBcG1YpoDyFr2XZg1mv51IjMan/lrDY65mNK6Gp2Gnh
UwD1n5V+SSzLJdUcygdhT0TuqBpfaA8E+11MMTIURJmIxTJz+XykAsEuSATUvrWhB3hFgZCsiCA0
3k4oPPtFQYPa0n/jWsLyfnlvAM8/u+LjNqLWjXvwsM66rMXEV/5ww2NxM1ybDbQc3SiNug93kzsg
d3An+8wC7/SlMbpKx/fKsq7HOa533ZMiddlaKyLYmOO31lgeK/tRI2uggENpifSYIydb+cBZgtFt
FTc+OQg6bUAx6Vi5i1fwn0ckFgjSmSJcHKeLUf2LOYAvG1gxm5fQupuKj0HbVz0cbBnxTGiVspoq
3JUeOYzrBqesNqJTkgbXYQPDyhE5znSc3YFsqnhbIGlQ8mCl+1aZErESrOiBOhi/cdv5w94ZEzq0
feG2M8Ar+8ZUTJZz5U+Gyv//kilPH8yg+DP/ZDJhJw2iN6Djf7qCmizy+3UTjf7nRQpgU/3IfQmP
IWrppCjWmFuRWOoEzZOxwjvsCJQbqEFU9DkGn8eZYA1S1gwl5Ib13RjvoSekh8B3FyokP8yBIrkI
VWKC9wS2rcAPA8RwybBqCML0GjuLgxZLpLd0bco5hnLKSyGhwHcRLABY2cHgsdJcKbvCHy0lkZWp
IMXoXx8cR7bbJ7CILbznwJ3VP9aLp/hrVTstzS938Aqdq+sjIqk5dvTH722J3PfvUBiZD2T3G23q
+LudzyEqnt4AZF75lGEsRSu6pWYY7P6Vx9gOMn5NP166r3df1/g0+k+6jEG43SkdvGiISKVY62HF
Q208AEq924CMyd+KnO4NNQgnxCGdZNv/PchNgnMS2zDQpm+qYFO1lQrFIFNuEa8rNO+D4k2WJ4Hd
CAOYJUtdOZK4uGELtoQZGM+pWu4LHHeTYeGeZNIp8ohDZy65fYpivBe+qbds0fwSYuocSfCNeQVR
U/zlnXsrlHbrumZq3fM9zQ4DZ6VJu61dlGdZdEIxC0ccxPU71fpr8O/SvvU1VAORz6vmzc0Cm22o
eBaUT/uicwST4t7SmVnyvRSXvJ+NDQStK2SgiG83/MWiLuXZPRl9OBffKBKuzyAhCIAFZ0Ph+Po6
rGE1S3ALb/SZ9UmDzA27y1G4sM7M8rx1ho+h7rKzsx0g3KjC56xnsdqoorfcNRHUS803VO5wYLDF
FKz8wRNkTANuO7jF3hmCYvRTWTqZCUk0O3luDz5tINuixQJc9XtpK6ue/yY/H1YuCkqQJTmcPnop
dBXA1PnutvwMLJbCbbY9NRbrp5SuPkFiBxbFbzSApps5pUF8CH9nYp4e5J6hrOnMWEO5BKmnyeWS
h42UGEGBJOij0yK8F7XtcphACf3DXlWtMOKzAsCpIAEFSKI0tHEaM9Jv/4fG19g+Kjs3rGWiRSiR
6McFxVmyLKYo60S1zWRk+ZohGb3R7qCdYFlnq97fKncVbMf1En4KgNGiFmH9Z3XEcGv5boIE0fXu
tduWBP1P9ha3B/+zE73lATpRVubhcXlyMXtFLTZVIjWMtWPszh6qT3q1PUEo+lRjNGuRJwYpgRkp
7daaTAQoiY+IkpoIOkHvmiJ6Kax9mgfp+/kpAhYaA9poztmY4BkS/P1ShFTvGG6scVx3QN9Tv0Fe
Ha1y8dqvnJvsKFAcOiyrZbwgj1QiCtU4MQMCs32Uu/QltkoSELkikmpWvvs6QjzNxA+mbrTIVKyT
lW9SFZvTYq3U0QtrJTmc+4Gy1X2Rf7KUMjTSXPCemB9cw4W6a7RJzFAl15Xw6aLmlaoJa3ta6BO2
n5tdtE+/GDVYSsTtsskUGft66T5ZA+yqpipcPy8WGgfLfkntjFwoNGvp1HD8YlmjnpKq1/AwDtoq
2lgcB7a3b9rgzkcxh6rY7c1GsJhnYRhcmQA8uiGae2NofDMZMeRFe5rEY6ad6Jq3Ysyhmq2NsD9c
iWXHWgXRYBWsb6RCRSKjjHdGXZJhxQYpjwZtHdFJs8HUnRxtMNtlyu3iV8phHLMy3yruxDMieKZo
PemXY/hhrdQWAV0W4OLP5CTs9jc+g284uUqlw21HYNMxlUReeay8LI/q8sx7w2QdX8AvEWisBcPm
BGIlj+nWkQYBUd4UgoFb7erj98qkiDargQkDeiUHktGBuzGd/ZiRlrR3mj2YOAcbOacP9BPeP8Pk
yGzN4wfGG2cGGccUytyiMhNYIIkzuup0+4bbyFbBrYrnm5p+kWmOF0ooDIOP3DB65ACTxjKjEKN3
WbjbVJmeh5Fwq5bJOJ8hGt4fgYP177zruH8Is9jepEbsewPCfngjsCeUnmHb44GWr3gVrHRMnH2W
4HzIXcoKKI1EFmKkxteJDr7Fl4lqXkwxRdgZpGfGbSwMQfcEAJT+noMtDTjBh81on5PG1IdQHW/F
GXOQ1tFT3KZqzvlem/d236dO2d21v737Hzne0Y82pnnxUaCB0L0iISIKAu7MTegQwWafpaP0tqEh
YXBbWjgpLm8F1ijPkr1VdU9qTIaW0fKPVPOd3LGvaUYVPJXYOO4/TvhfSV52aNo8u4QDFdNf3KTm
GSSjQeQpbnRZISYnay5uaoynFk88Wl4bW5ONMueVQGf/J5wNRcke46srFDYaq00TKgn3hMfghXMX
I62YhN5oUn40HfA517XJSBJubfoWrtV369pdmXzpcXofEkCjbefN137byaKPmcJKC3HuhDSR/KFs
pOB953GwG8f2gNgHFoXSxhJgkJ6rvD8Z6ES3Wa9LQSKRbzBAa0pWz730GS6X/asVJmpzFPymVSOB
fYdq4H/Ii35yJZmoyNwoKEBEoMbk14otVjceFiqIaY5LJ7BgOUz/cZOGhHjCibSS+nVE1PCAJBlo
sDUr/9fuV5ccLZrGn+HBLGVFfsBgXSCsr/WZ8lMUp8PYVTfk5nB0z8qlKvKmBQHuxmKUyisXAs72
1tUd0MsSScbpLjfy3/VyOVh/AQMJnDRNbNjhuliUJw/N4ImeEjQTsB3IZDKe1YQE/HnfifhEzAXc
GFwJ3VJRcOyQRY9H4H4iaZ7lYoH/fUPq0U4a59sBDEk8Y9/8aHFCWHRQW+Cfi/JLc7V94cB8mu/y
sf66rIC0hryiWF+9Q48KhRrcF43Dq9DC/7HfLOl4la/P2LUFa2823sDsjj0JeJanNsPmBSwYWWCB
L7aLX3JXvVlONjQ4EDlv15qldiouVIrtNQMhMu66RZPxmHlHxDwQBtsTE6L3IX6XPDIxUIOXJMjf
08vSAHT2qx12ADEdltWYjObp8gT0qg67N2DuGVWuo1B5jLxcTCjEwg5LjLYxiuBpLuJGLRagbsAF
sbMYjzY0QsZoX9htdXLbyX7J/mCIbrNwkYAjLtL7LqFpNTseFN1BOQ12sHK2ng0kLHBZUjzBUUC6
D2173CrbSaq4/i+Jr+YHoYBd0+LNIVvD7k9mb9AypO0osPNnIclAAg4IWGZ32r5CkBbru7AKQGRL
i63k+hArnodznRSdUHXAogo1Bi21SPb2Ucn7/80n1U8MFAXmlTji1d1IIFOHNHkmot3nqKclabcL
TIsLavHDJXOGZqVgtTM+nqw47xS5+KxO3Qm37wBmd/R2qov1+V1JzxgmXFZHrPM4enXSNXfSlyYt
/tFIuWcTYJ+OuooZo6c9ieDbziiwXRuvdJthmjd2IijCSPdTEpXZA0nkQO1m3p/pQfa57gtPRoCh
H9dIZWV301vGHToCWZUYVbn62w8Rs3o9W4+QOKRBPuOTd5GiiGhnWG2Vn7pZIHYzNVU5pPRDB80Z
uXBJRjDfdSC+vBlardUyi64n+WUjpY3DlERbkYeaUZBVEPvbglDzZY/j/sgd7g9w0jzxnTAlrFek
uP5Y8hnMArf8LhFeEfq90iNHuDAAPFWLdV9jhrl1RtlgMIMbKyDik9tit2cG0aGAvnUpJjEIKn7q
TlY8EZI+GlRBfWWzpRMnx38SvAna9oPYCqcljtPgryK6nv9mZF/kP9sDnnpvo2r/QmMVaRxjcMcd
DxIxfNfFHj6bOr4mmTbANfnrbfIfV76TxlJuCCLRc8cxEgG5ZdmAWkYxoc6cDGcWSiXl9/B0zh6L
rcAYC8U+uDZQ2skM1XLoBIE4U7dG8NKvMj0FeLZ9QnIc1b0ka4SdZKxx3vrJWzIK2B1nZ3OAd/qa
+KqtlIDCh2zt7qsxA1R47BMKlyBpmFM1xgI9BcUJrXWGZv7uHtP+hMK1YBYtQ1Dmrlt4wX+q0rj1
7rHikJ27UiYuRi1Xlk159QvVv1qKYi0fdPjNLTFP0QQoMG5Hfa09dYXTaytpXom42Vo5vrol+ZpE
57jk/LNRW7l68/P2UTrj6dxB6eu9i9IzbOHvORBH1eh/0fb78hAP8iaOjt6hyb638Q7uq+JMH6kV
mA6/rmmUUxjHZgMvK+XQHLpKB1Me5KNSqylfKYJO+09Xl9cp2dO9ApMX2nIYKmMq1QNkIZoMeOpO
MTALNDVAyYLJyZe0puR4g5ICED4XIKK4BJhMqnuPysiZeVkqcpsUTtRm2LWeiQvwBcLRrSd0Awkq
oeFnvuTCmzC3DM/DVOHIm7ZYuMBEFoPtNTFYqneL3jjCAugsraqdzTXXHGYrshtfWy+FaGKYcwHK
hDoHzLcNRJ+pRjZdZcPLcZ3s395nGEK8wNaLnACs9oK2d7sxvLGg4sKwjh0a/+CWvz2fz3xle+2g
XQgOfTuQAJPIkIaqxo6XMnYxbgpVoZW1/8kMdW5gNauqCTElCBaIHwpciNtjLBbhaLt++VEBebJy
LkEWWC2Afn9Mchu0OPEOpkK37cjSiHE31b84px16C6rduVDqDHmQVDCkjtCrOS0UnpopN0EfWPil
RbL17MI/zTrRWSsOi9lBiwax4MnzDH5ng3mu8xWWs7I0coLRxjGZ8+N2DQhWB3iESwi1cLZGcjXU
2SX3WdZS3u6F3HgF1CRVKBclbxnWxiTNSkhjZ/zx/lIl1yt2pWuQXMPupU6PazyGxzlq8oQggpLa
w21svkQ1veL7ntRKy/eFwitinL1TnFHYbXmYC0J0S/wbLkU+v+luBxfaTGSTR4jn4cCRFDJYsEaj
Chj8cuKXGyxXOWuzjzj/dqspgUoIpZPdRaZbPkyDGNzxxBg0cPBW+bOe+oqaVZRPK9IS5X0NYSN+
vtaH5PNaNTBeugpNGf4X10uqE75Q85Jxzu23mKU8/WfzD5iWYZbfD0D8RfHzvPVNtUcKqzyyIaGQ
bd4el9PpSN4Lz7p0onl9AO9ZdDu+HAiVnv0Ooc2tHLAojJRjhruz9rrqVGhFNrtE+3hbtynhFC3C
krNHKEMRbw8WwIqEGsfodr9q3arzWSFXHplyzLXeiHak41Udv3LBw7VTRqTm6AbSPOxJ4tlwIQip
9Jb0OH7APyccdqyzQhtwjQAWf31F6fiGfwFCEIinC6aOMYErtpxcpsC9MLOhCbCOnEdmoitsZAyN
eIE8KsrQtcRr6sHK/ejaNXtf/Dxz5Ge1CQV/7D4ZO0UJgeAv37nAJP0P5VN3zyrlS78S9eHmgm2x
HsJ5YxzTXrd8vVktA96W4yD3ZvwXQBxPORohrx7zphf9WQveS2idckiBHMO1UiEBXhxBUvr9D6Uv
xauNePfI/vM8W9NjxZIjdkneHab4Q7JvMYRRT7QFVL1vZ/kgLUHHjyR2juHM5dMG+RVJUk1pMhWL
OpENrn6QbSYK9sqrgln7MZ4b04AH7KI2uLEHzAhatAYjKb7pWA6eLckbAba4GTWB4XqSi/RbeC28
iKbLOZaZQjVt+1wSBZGJHTv+ozmUSLCtNH91ei0BCjSozZ+APgtMjLKclFB4H01kV6pQQ0xWh2uD
v8sLbEfgXpxEJU8xAO4AeVHMHtaM/6gQ+gHuSgBWPRZnHpePj20YSVMM29nD+LO/v+59pSbRSVga
XKlXl1vbVLh7s97zkHgSopsHZ4tEY1U3KllYH8pdgpj4cZ/JmmM5JBN+KeaDyumRA3qL5d75FwvR
1pMPiEhje1jUwYGli0168YVIcxyoHs0dXr40+fjaa2y0t6Q/dl+DcSw3H6oF6Rs9G9G+DbiJzcxm
awzW1mcNqrIHuD8rZ3STmhX5vIPmgo/EasmFIFceJcWCs4Mj88CPAJuHZo/blCx06jnqH3GFl1Kp
KMEEaF8gJzrX0iuMIYuyuN9WMclnByYzS6mW2OZ6CSIhSFu5f7OlGb7c63uQUDBTtTe0NEYPb5Ov
dQ7WRcx/zdceqIUlSXzmp7dqprugaWK9hlX2dxjl9maWq9UMbJXeAIVP070lp6BaN5soH2PVMang
Vumtm91MMRp6OOe2p9A4EfEmx9uVPjnaIs8pJy1rdBS9a9Yu5n8HNrNNvZF1oyO+fcVQHI06cQ8j
sS1dC/+aXaEAbp/zAKdHrEaSb8FdQ3c/qQifkNV2AHoIGeoJHxQkUMh9cgCqX2f6LvnjKNBNSveU
y6fZh5RPLBO+RI6EdmYn63HDJvtLmdeVzhz83o6h5TBMFKj0uiin5G4TK+q0xWL7MLjlca8tXe0j
J4a+29IdGYY5TCPamVN5Gcx9PMPVv9c47/6ZmrS6SyR23MpolpmQmbYLznX+Z496HtpY3tww0RZE
lB6Pa+v9fSkfPzVAGgSrMQ1XE97z52W82aGM2lnlqcAtVtWHZNx+qJkYh2T0wFf9NSSMrzNFg5We
4O/XY/TAEbOLH9UYjeNyK97yfLUCgUz8oxhG/cF/D9yBOVEdqhzRS2LAOzQ0fzgxhfKpTHtZS+6c
/Ky6D6CkaFQgYsMr1OJLtIaQwzXoYXzoP1TiDe0QYc8dx7bEk53kxxwHeJMYJg+LTkETkPCiAZ4P
L6yQu8kNjIVUiMaIm8pt7F2ySVdRl32vSZeltJCABopH5mktTJibZ+6tObAQA4Hl+fv3RQOMgwxO
uegCV5mFQab1Lwhsb3PDTsUK2uERM9biRspJ0T7PVxAIXaqTyIbEd0ZHnjws0U7+Zf7dgbd7yktX
+I3BWVvGzwT5Yml6mtxUX/xE40e1kyzsNElHu4plzyHk0nyzdrzEYCCX/88wUi2yC9+pesaOrLUI
odaS7MSzg/hnF1nZKaTQFbMjwoe5XoAwbMTBaEeQJ1yTSy6oRAYFBC7MGAZkj9uD8chzNvwD9GtN
HFkEHZvw3swVJQ9c6RZpqPZ3PbCEy1TT/nmMh5pJDJS8ywWp6BAgJOKmz+OpQA9eK/hqUMsWt8r4
OqC783Z8CBc6JUHQlFzYs9trytn0HGnAuyNlmpCRagKY0aZgJmvE9XOeXIMG+Eq9D/Zk4uMHj3fq
UnsLesyPnEDF6aCWmpubXaZP7GjkPyRA5JD2hsmdXyFDVMm1u1cJGDNJwEbErzmFUvKW0HvZ3VTT
Tbur0wrqNAFq6p/vbUxpRkqB/23espDTLJoHH8tXzhhxcoINTkHysLpB2iLWM+rmlBMsaPBeIw8r
VKGEkI9jjFZh6f72J7g8Za89AcqZmFAmnjqZ582CUNbHo1uVnbW/vRxXLeXKxNEoeUFeXcb4G8rp
ZIZstt0xnqPbj8KmR6fhJ7dgNlJ+zWZSGuxx2CodFjok3xsvL8aa+erb1OOGEk7Kvczxjies5+Lo
njUqMrajvM5cY0Vs0RrHy5Hpnd4kr7dwwFuknrcx7taTN7NhUs5Pb5kTIk7bJ2MoDzjAiaSdCGVe
OWXNF+/HSUJb3tTM+scZl6Z2abQJzZjyE4/AOqnEz8siH7H/B5JTdwHCfhCJI02ythlAxNDkQ9hJ
8ts7tlmzFeqwI9Ih2/TVWkKYKrnR5scFd78KqNL5TOGBGX6zs1ZTNO9xfwMPjDoP2UmfCDma0e3P
sD58cy5d0TKQrD9ETYO7b3KD/SD5YKuCvjZhadQPUXVuORP0aadYviGum9CGW/fPL+/INZeGjcu6
HQKPsjxZv5zw1zJwOGnkK+U8HkQKl/E406rRkYOHv49eWTPthS3O3IJ48SU7rLO0dKPsQLfJJvhl
ObuytITJ5ToWbJplb2s5LZGv7N4/w8vgRO1TV4XpAODb9sMxtpMPu5cJVIccab4ulONJnvQfMm2d
MDWYxM0PtP57lPwlpRRoKr1CBgr7BRRtjKZJh/P3AmZc8r6NnDrZbC626bTGZwaWZ2SA9QVpCs+U
K5bVva/Ci5iL5Icqu4ZNepGIL6F2d57k2BiahrS7CVFiV4Ax+OVp1eNds/C8SqSGevZjDaZgtvHa
8rF2uPk744d/1s31KprxjiAMokLCH4YC17lrtFztEPLyCugPqL3m/QoIh4Pet3v64GUXG3lyOKyL
VXwKK6CcjXqqGrS99p6eKje0Bx7z2Q2Z6xXIXsRK/4w99/DgLgDQLzPsXXlilo2Tbz52VdxHh5VV
uLqjBx1ybde0MNqFIWxzYqow4ZgS39fcQYPFrgtceSLPUbK/eZs8L/jg3RQ5X0QdDCmuSgT3CoK/
6jo9tePNLHTtGfHsRZduyIkFWvhz44IU/Us4jiqbVEFz3H5E7mKbgnhrjDvHPEKKMzy8b8juU3Rn
XYFMTWuYxw1QU1SzgreZ1ITHIYz1W8Z06yqy3DbwQSj3WIQRUi8LNmhgR1SqG8ZF/Ad4QcQnPx5G
So4v6j0jykZZ3gLjGF8j/cpRCHc01q6VfFRzrmb/kuqnPO8H/C+5ECmMOtAfLspgIAgEhsg++ku6
WgUg6WUHzkfdnRKJeGj4dc5BtXTo4e1ATlUzLl+WA0sXeOQLbrAXH/aNeQNOCMvc2woPzX/HjXsd
di3AFeTbDBUEgS0mrVc97zK6KHQyzU+myienYZRQzhEsoWmm9pVGGIMDOrw2yQyp3nFq7Qltfr2/
+cv9/aiWkbwbjsczUMbUmAYIN3Io4RRtaJ+2plkHj0T9O00dX/ASGE9MveF1khkKssHGWPIu6y41
QOpK9src16L7FVfNiD+TGblp2LmBUoo5u2SzYzSJJXmm3pNxka/DjU5QjsrzZPvfre1dtvs9J6cF
0ioUSCxUjD+qIchdYxsH658L+L+pQUAMPFA1yLH84NqRasKY1iszQQBkAQo2RjDfNIfbTud98lmW
tfXwF92gA26hK0j1T1hg8VPHyoCf95770FmfH/alTOfnErMf6g3uQQk7y/FCTH5FxXAdjiegthap
TXk7+l+Tz4J2hATW8yGLzr2LRLNYwFxMJX0JXmvBqht15NykcyEgb9LnTW691QJ/z5szZqHJHdYi
NRpz4AmwrNqc+s3n7XCQzuB6dxpOqVq7d6c/CPbaBxj7TzZOdmnHlnbN/uN2r8YuVVBKIB6PM6sZ
Z1kxDmADsX/YyBjivP33UixEhuHg5n/QZUlSKAOVGGy67m3X2EME1kxrDrFsE5LJoHvUrRsn4a8/
ZlWRDDNPkRzjOQZfZPTHZ0/IKNZxUQohN/ad2v7tAEpR5YqaCb2z2CY8OSDQNP/xXig1MeaMP9+8
Wqs/qxVkEUCOLJTdcuElA9JVZv4MB/CRMvafqRubRdAUksLXkXhm1aXiSqsTBcogAjF/lQyKihvx
HzuuAq0YBXREX00nOjKVE4C8evRUUTF9Di59TRw/hh74tMN5I0OA8dqUVpv3v8DropXGVsqdWyW9
7hB3oxnxSt/lN3EUXjkb90dN7IpURJDgUeSp+ifINH0nXSyvZxf4yk8X5lSjXkHAatXIjLWxs0WC
DO5ZP/KXpXiLCR+dBkpSoSTvEBhLDnOY13IliqtVTAsgpDVIlBYcZdYWuFOTLzuQ01X+6XF3w3/j
096uFwFT78z3CuAnAJ2PL9mWfLJTMcIBHHDj5AGJA5deeGUtgFefhkS+dbJj9YPrxCVKpHzlCE3d
ZjdEE5Y3ITCgtqf6IM9geCJKZh4o327IUSNGvfz9XcmhNKibEPjNE+sxyGbzTlNCkG9ctByU96sl
+7qAou/W9rIDjT1sE5Ahi5UV+gn1uun8FCrULPJFHtWdstGQx8JKXdd152LQlJrXbJWdZ6gm0reo
6FeXENdy7wB2KM6FCtnbF1mau+dFCx+pST7Fj491V7PuUsVOOyeERW1UdG3mUMLAsvulND4EsQeR
6bxHUmS5JnSazt81d14VEKdntQzA/CGv2r8jXyRrWt5Q8VTs695rKS4rsFT1ywHHwN510vv7WhAt
gbEMB0Hzy6YE4AACgnS8GXeSZyJc8NZig6dxsoQyI4GJHG/5yfUcfW364FlxjFPKYgUoeqoymn51
+PSMxbcO7/FVjPTC8lcm8idyq9Q9ZDLYooI/PwQPzYXDdnkloSbjdEQIeLjQr/4GRj6fzaFIUDAq
X/90gkEHfm4DtJj1UP/bfMVrmoGAEKEcZYjK/VRMJp/eomOZYSMLX1RuUY3Tev6EDNCsLp3RU5/W
iu+6ZoHJioCRJSeBegSv3HBbhWi8B3epDDY5IaBDmSg5hka72FPdLuDJltStQC5zl7wM95SRDzPq
zLt1rLLcf9fncGQEImSc7WI+GKRK3a+YkETlpitiKlLDiu3++VhD2LP73oZnmMJZ4vIB9wwOq5vs
NouN/GRYjmabPo1SE6svkv63RjzKsDozOOfbVyFGx0Hrgy6WbB3ibvRXOtzMHZo9uQsYOeBRVIY7
Xq3KT0OqskfZRkq9iCS8oQ+WjxuDmE+saH08pPstidxt6C9r+YaBxA3w8HjIqcS1dGYkoyTkQOnm
Gqs7uqYekxFsBy3Re9Xtks4W+a1NtGEMl4hkiOTq8efJtzEAj5gyhcYIOagpEZXUU4EDlxfNvY8/
5xZmjhQD5kDlwNsnALI1mZIly1qhO/cS7hc5XnWMVYLrkERJtA5IPV3+1ffEgGrPIDklDloBGTE5
dC8rWzpoQiKMVlivtdhDKLrCT7iqbVtNqXbcxyAM9jfUjkFA3IOUNnakmXo/11IBidN7srCTGd4M
g/B2DVXuvJcbNlkibOw3b5KiDEtNv1h4SpXUBSZD/LMVHB6yh7wR3veR4qRUsoM1BJ8P9gyYEZMK
S37jPtVI04T51CeuSDboz8CCgNnzRV48qjIhE+U5ayieDoEa5bmwQRLDBFqoffoSkmXfDJbTbQzw
y/tYyj4ro7vb52qLbZqP+Ic1I3+RsL52HVwTEw9suNBgrWcXxpl74LhZfzWqweSvJdrWCxJNFRFJ
F9FJhlPwsxgS4Fl04eTuyQMvAA4Nk54fl303KG3yB8f4IA5GMwUuO5xbjwOXBpdJWVZ7ogPPxH2H
0rLkMe669SXnfMWJzkz4r8OlBCGy7qKhJAAg2wQnRQJH0rHVvN2IbtV5ye0m/BK4+im3M0fUruOg
c82zePWTEXDBnHa5pPxB/IregsgA/VviTx1xFqP+dK/kn3ryYmaTIrFFyghgRvOi25E2vGfnCKYm
x7Zq37hhry76M09yRjrvXLJncpaVk4jVB38q02kxuZySm6LctbBBI7B6Tg802E+c/nwOwek2ymC+
hMzks+PbAemrKsn1/XyZpOz5XFYd9Z+ArgfplHr5Lggaor0Cle9PnnSD4DmHdIe9pUb6CJDSbbpz
nsMQymvOvLDypdk0sFn4Zyh20NQohhBV3uM7QNKe6g+wU4SrstiGB+b8OOFNGvGQXRh8jYt2atxa
InZzm1+/MSaw2qaKDXYS7az2xlVts7z9wLdHow1PQMA6yLuTeOhpSQXrywxVKIfvFkEyLD+8LOTI
vqXw487k+NqkPvvtZltG2T3et4gZqPbTUqvT+zBXG5yXlnU0u/kDU5nxEE29VBxYkXC5FxJpLdsH
mCCeclKW4nTwicLY3Od85Ma58V1F9kQd463bQ3Pi6/xHndO/qrnLPsqeustJLFIAV3Q63k1LCmSh
pg9CQm+JSO2TNgcyAy2A4ILzT+pSssWl88hV6z1H7prHBzVseVCnLxk78CZxeq3Ecmm7eg4i4+xg
2DC3mSwDQ6rNAB2UGyBzb65Jt+3dE6bK0q12enMZm9phnjqMo0XsFSrjm/VQ1ubZHtJwM0dOMGOB
pd6fuL+BV7ztAkn7PLf0aLHQ6ULCBgh/jmvxYHLGYlwEysf3pVehKwYH2BC5rFROMnJX4bKhge3E
q0V5gjVkepaNOVF7R8rZKWvARAr0zLLl2w4I4LPXT5M/RKY0FAzsPjg/bW3KUpeeeW8Bsu5DzIBN
3f7s77mVfiKyAEN+8uxU3huHJv+mQhhwG5u1l0xBBrCnFG1NDWPeQbbJT8h8HAIHKAVdMgAEetWK
iYvB81t34Cnu+xVUDM593eRrCoCwIeW8euxXwzkuKrEb+2U9n41tDqXPXIH+LBlMo9imU31WK2Rw
H3FY1SYLoGaxF0x/1BVzQ2a9+xL2MsbQQtGvh9urVyrjcUryotV55DDBQPyS+vzjQLL+QijUMS9b
NrHuUSAedPb/lusxG0x+jaP3exFepJdwuP9BWtQEQDshsKex9qjaFU5MjI3m6CHW/VskUPh26OQb
W1ZyT8dvpJduDWBKYR4Sp+C15uR+ZHOmaubq78Hqex9LVA438c279DjOwT1vk8STKmnMhlI+c31h
kCVbx6s3fdzzUIEq37Eo0z7lhELq8WmFosD4f3cclHm+R3jmVmLoyNt6/3ma0u36YqNp+5PfxVZi
MjkunWbFABisbsjd07f5ImThtJfbBGn88c/+aep31VkWBimZyXnx2BOxKcC8Vi7+HR9FcIfufS21
w9n9W1187lSbhZyejP7+rSnG6LtIhPf7utR0rXULEY2Ao3zcO0KT9G1df/YlEEKHZ3rVLwOwX85Y
DZrBrhoyvcAVXzaSAff4gjNGc52HPUSiLZqNchuA6WF/EMorpIxLhNSiBb6heHZuSxfFDCQ1SNX3
m1DqYXEMGud7iZ7LuFl/qaAE7x+nC+3Y5H36ef/IXQci6g5cFighpHtFWljSYucM8P+TKKIgf+up
IgxK0Nzkds4H0m3GJe+Ah5hHxY8e8+YDvFqZee0CBU47jXFstgHLI6eDn+SW0wPKWKx4FcyxKIAd
qikXp0vq0wUcIIRUxCAmx5lkYnncXMOZsBm/EoPuX7lCAJculhr57BF9ri81TSxXKJ8UiVrLx3xm
C7t/TVDgpFEMwPiIsTCPwdChXvBqJ3cXzcwmvnKshPH+HtKABRtfE/rpjE82EgZNLKKC4/1380lp
I31nTHyBCpsDC2uGpiN4hWRccXw2sVwJv5ctNEFvPial8lDPhYUmTpQvgDHL8PVjowal+sooEXdi
EtpMcWYK63OicCjcw1m85IU3DDr0BqU0CbaDZ0jyHlUdCAJn2fNk+zuywy4kFTrEAKxMXq1Tqr4/
+yxoG3lQAYVTPLGoqPv/QyM9pTxiFX02LBk6/TUSvN7ox4zmcXZ1NmYbBbz/qIfIfrLP6bgGMk5p
SqbH5hFgsGqLKbwfRQMiabr9Ud12CQGmGnGcXnXs2ue3xf98RW92LRkwFjWC48bksK69pcyemuPm
i1ML1NAR60rVE1xttMODKWmR6ck/u+YenJxj0hYDPgLaQBbNyH72Jkbxsg5aQYlHgoZ5wCQHFj+M
XXc8lMR+Oh52QiGx2EVCagxxzV+zDAMRfaFSHlrv69KYYBIqSeoT89VD6sw2Q2hCJCkSwsteqypC
0d3gPi8zLiblBMGerj1DXToHLabP7wiGiSVieZKIB0wIwmDYA0w2kcWtlnvtjQrNpZ578zEFkJ86
aL8kG9sJAk9XlIWEmqOGvcSqTxPXM6tCkhFS5sWDGL/iRWCIt0GPrDxmhfpuxid68BY6uFvYlX6R
7Xkonytr4SlSqhK2Hiq8xDoEPtekqcXXIpHCo5XJTGBhpngK6SIG8ssEHwxyjjKM8zfzNQoIdfuL
+tS4d/THXVALghznRKQC+qw9+3wXIF+r1Ey9LitGJT7ODwmkj0x3F2Yvack46XzIh35/iP2EKpxD
EWcOJuUGFfAAF9wFffisf+WXze0C9VMX+O9/octYsMV+FUHTEo4TyxmPUBvxWH+kT/D1wE2ug62X
/L9HfbiEYa2OT9FP/pqKaopgFMB/sur9gxTfcTFe4c591goojrPow5+IYFc0SW9WuKcdY/XpTZES
GvSjBa9mVfM0yGEsoipv0NzDBT3xkQMnjbD4xUTFpb2jwqVooyTQLweccoaPC8IxyIGUpXzkVHpq
9j9p+pc5OMnas/i9fQOSERywIgbEnPK0MFyekWMxKhxr3JLJI9nxXE4UXwFxYegjLfDFedSmslGK
lFSZznUTP+ByJ/lP9Tuy9bph6vMAs2NWT3CmKN/r46A2oMqaYnDDvlR7FZaHfz7VlECckCT3EOX/
OJURq5dei17l7O2Fv/r/oQWJe5wrxFBm6oQ/0lIcOHZ18NByueDmhk5Mo8aYH0u58rxRrGWKQ5HM
x9ORwomBUxPluERslncpKHHtG6kR/E7uletC2j+AevlSwuO0lgxUDr9VXlPRZwZHaAtIazyDUbPY
Xc4ZbppymOCd1VDiSv03DLODndSBNSEkWKaCj0nQvm7OPXDd2gPrzw7yUOMYHtyiAspGnizYUbIq
njGrCFGS82rVt14jVHM6vwo4FxinaVh9bJagKXqMTf6oFMk66AtY5s4NxlA6Sv3xQeCbUrM7hvIC
IiUxzYmTfRKB0+CmAbqsVoCaVDBY/q59p/yzFEoMuJOheDCVTWTmHq4kcg3ji2NcP2oAchTG//im
wP9qpRplFp/mJKgMnPzG0WmZkthbkrIYl2CXxPqW7oEygO3AdgXP5W/4qGV6fbJj7MLbXOcOs8x5
CzQWMv5/xyDmx+jPhstrHjoQfXq/oWI+Vh/RFuEGBjkexciVZqxRAyQrm7FeNP7Ru8IHx//9XuZn
pC2PCNCxCeUz6GHruEh0tcwionLjio87LlZRs4sSfHfdjdGrMZfu+AqTN6G9jjDsxkKG5jxTmDvj
PzDdnowQeKo0MewothMGCKEFdikX6smOMcGevMhGFiD6NYKx30kSNYHLH/0/cYjGe7zpQ+o/CS6U
YcB+0zAItqRfTGya3DMNDxOHStukExmWtd7zyfyEHGgewtTXTDcl9cSDVubpLXBFGd13x0EXCgLq
tddy6Oqj7bMkbFhN0tmSN/t8nW9Q5mYswyvSkHbIEMg3n7WXTfvZQavatq0nd/9onVGzLo0KvcuD
P9j2ogPgrVgBl+/NGOk0frhpgNxK5OUucW2iszCf8zBLj2eiy8X4yF2U0DyQr5ykY+WIpI0D31mi
iIMu4B8fZvk4X3/yKMcXuj1KtyYozhfRd774/ht703i4K4ApoH9OHn1hXoaeWhehchEqo4SxtyZb
xVkKfj8wUmCMXdlU9Kw2vaXzJNT/p5CnBrfCVUA8Gk/76lRT6OejBe/yrnZx1PNZjxhf5QqlZX/x
w4mkG7vvMJVavv8wxMChqdzQp/FofXVFLYU+7G85xKIsggquLv8pAqGxmkjJhJkDlaiNwR4l2D2P
TumZ4bsSPWGL+GZ5+RfKsHHh0aKcxPL22Pnx4XbYSyMXSnsTsN5vhUAfptgjwCyL9E9jGRH4+5OT
q/HvfpCn+kkCaEc1EIEBjpqdTCBbxXkEyenuXKUw8zrTK/vyjHUCOjMX0BO5Fq1rZinfBPQPL0Sr
Sxk2jSz5yh0YLlhtdywkaygzaeLke4wf/cKP70hm0VrXX/pWsn3r7Fqtp2Fg9zexoeE07ChPPb8J
J60SmM60/aUdkPJRVKB99rzLinrrsdIy+PonKWkLp41gDSRRHjJVi9N5eNDsqB5kCvWy7BMnHY29
8HTby/i+ctRafPTGynjMBK4y4nJK+BAVbscmcDm5cjBE4odL6IwTti7D6rx5K08rE51O+RsFDNwf
yO4M8AlGRhv3CXYqlrdQz3QK8vtmWtIe9cVZ5ZPtiP8aJLpCZ6cmd7dY75l2lsy9ubfEYAhbEAS5
zTFPPiyHjhRPTyJjmiCHBcMlfLCODltmmeAqzcyTiYc6I7Tw/KrZ4FBnsiOcR+66TLJqLgjdTR/E
J+5TYrjPbHBh6q/YBD/yWSv/GEuHrgIqFTh9v36ChSqOhpGCeFXxVeIS8kY57HGr3mIksCcBzZYV
dAIQtSwZF9SpSE9JqDgEjG1/0UDxQX56QxYZSun+/Zxd5KmEOBhYTKOHknckhi/bNaZnVFQQTQcf
g2f1wCMMoj1gsG8AUS0kK/cx0FrKPSDNX1nppx1xMT6VRf+ebtoUpoZRU962ve4lz9hA4X8D24zV
f60CL13tBsKKeReBu8e7JqPZnDRfdUlUcPhiifUIhopQfAcD0phCnEgFYQqlCWxCCdhHprT/C0Px
gL+8k6lWusxWMOXuuX+P1GDI8pM3VyBvESksTgA/XlVIxSOVi0xw5pmfVMU7/kvVJ1+mn6nfxbFn
CE8i5vmKy7zJlpAi2jxTcJy0B5vH8xbHP8Uqa8msv9T0pbsuAHZTphn4Q8S1BTWy9MwvAJA/N9za
AkyaXjJYgpZ+SjgePv/t1syZKelyCRpJ2XdpJSsGPewTCJ0xaSZ5wXfT7t3iRa4E+6VrjMCdA1g+
Rr7Mh3ZWmnov3TYxIzfuI3w28I3WCmjmMNQXobLdqgV7rNQ4HH1o+v+FRr9XeWOdHL78spwo7tec
6S60hnWgmFBdhcdvpmiKxslTNNYH0RMdAMOVzuJjSbauERWVT4Qoe36yTxMR+GEqihO1cCpvu74t
xbrn/moWtxaFVfJiWIEAT+KMfgbKH45DOenqtHkFRCtZP0nCNWkvKc2fxYv/fakme/qAtx7FyIe7
8wLDXWv0ydperWlXkzXmTuK/K1qUh3o48oreS9iafKvuWnPt6eez/XJG54x1fO8BHMkZ8/LAxDQq
3LVEgNbAdaO7+58WqZkbkurO8EVPeZ1wgPvHX9w3FuCffSvzjvZd7Xf/oGFuur/EiDu62fVnIxzG
5vlJ9eOOPpY1muOcRFAy5ultaw1MPAtOiWXe+mdkZkjabDplM17mbutysjLYvwFDdXZnG4kQZWLl
WPc+poCXDWaa2EFPT411lB+bELA65oB4J6hyhqXBywWQY6T7cZVOpTyw8M+yOrtaqmT7oZxm9bYd
9hVrAzFDEFTHpZsYGf9eLfsNQDO57hIE/TLLJLZmoOtvtOHysgN+EBsx6hXWS9BoK8GCT6/48SDm
75BBgu7QPTEX3AHfWY+HzX9lh5JpRJO9yqL2RhO1jN3febflmgxVtRGT5TTfqacJ/f8DH+b8b/hr
VmWF84Fb78LLE7qWFK4vtNmUjmhj5XACyUa7lWQDoHk4IPwjeRE/oHtnFYVinZu0NZSsYIqi40kd
2aoK5HnDpbfIbB91GINqZp5579deiO9Ei9qRrabkiG+23zdjGnsIS+Wmip7O0ptEctcoNjEX2Dto
3deWN3FsjFfIhmb+sUWCmB+nfibKlbdSTwJIyC5w1gNBxlZyrwvJcvckTisFe4Pg8KDBH9fEV2qy
fJKbuYBb5d0YcWsgiYVGQeywSaq0b6uAP3vFC+lgaMMSza/Rks8Vlq6pKmW8SXFv7xhtyZI2QNDO
XQnRwu5gpWqz+xPyHXUct9GjX0pOS287v7/2xgCyXyblyfgicyPfxKVLacyRC/Dj0mjCmmYFWR+/
1PcgtkvvNWj7E5FZdz3onbLQjrRDQfS8Yn4WqjuZ3KLX31PHBONQjh0ChRSy0L9JX6JlKVyobbkv
fpuTtg0pA6J1/3Tjj4Hx6yyEePk/oz9ar3cIbZFHnO8zdkFN+71gTA/GQibDjjUgXiEKGnUSWrJK
/o3Hq7ErU4yxp8NZhjCDPjifGRJ5RYUyvva8JQp7QU5DTOKSpUDJhfR2CezQiRLD8oIbO+ecOTqX
M3s0QzmQcM+90bB55X683XPzLph4sykwQggXtM8MgzyJAyilVLb2d/CzbLXbd41J0/3Gtt9lha0S
NXl9QR6P0fKwG7NCjbFvSrOX4ajxwzgLIUpBPXldF/VEMn3i11iR1ewqDj7kt1EWRUAwShB6CMdV
O//+DV5VcdpSsvTu5bpbQ7lACZn6pPYS06n+RA7pMmQvKX2wAMeK+vAI/Lf8vrVBeOjiOzmZS9zY
QpJAo+wscyDAYkT4qMqNFQt+9UqwJwWGAdI5qfX8zidu2fVfD9d9dJjq5pINj4vaFSQUu8ENjkSM
x42LBZn2JrN1fht0n4aZZxwdzsE9eqnAcKEj1IM0dT8OSMR6I+Mp7Za2j2W6Yf1x/khCBjNzP+yi
KOtp6uL5D6dDVOMkCNuQanaGMsmcPlBzcknmlvVy5tRDv9vxdN90mKpdh+2yn8H/V8IaKHK7eab0
BbcOIkR45BBl+nE9klV3Iwp6m1Yz9AHRJqeaNpKq+sCgNZAnBnotbQGlVktHe4cCgjLMfvLQnSgd
PRUlqbNK3GBg8mC+sngBmRPK0OcZSi9Y8HkaZF0MK9Nkp4e5LTikY8ADCD9acttFUsdEcEPrylT9
tQw1ewf+bgqY8RHHl387fmsVAomWAeZkNzlh6moMhPeyFruUV68uFuovlA+T7C3fyWVHDvFKBeIY
4ZdqD+N2hi5/gYhxGWscPe9rLZcLomFFinpLO9dIn+ibCgBmNBPuTN5c5faYBO+9qhpf8t8/FFdl
rdLVwg6kXzyK9i4ae+5cqwuZa3gRP6KPxsimnGb/fLSLfpn3k2ubd/5H4hAoCmYui4oQgeStOi3z
lE4nf2hrBuRLXcMmis3Kf/xyHdgroNeaZTpZ0OhUGeQkRXfQSoKA5kWSaBX/btOzVd9D/0ZvlZL2
Roh1HZBCAG2T+ts118zNKzrl9d9qjoSmB8BFLLpNZ/3CQrdJ9hyZCqC2sFjb5y7oAhGqDk1c4bxt
hGSd8j02ud1OY2bNV0eUvcnAYFjesoNHCkHEl9e2xCY0/qapT3fkFMX1UgljSF6HAfl7FuvxUKC5
XwpYcpt2V5OYwDsqIcmX98UuVUwCr2yaV5MQIAGgE+MJvmV4WCP3NXGE/KAtEMjhW/eWACkXFAXW
7Y7zIdDzoqokOZNbFDjB1lAtCjYgYDxjqOR/rc0w5bqUk/zumU4uoYDkTOhnvs9XLhwbCbNB6jcy
ObFLAZAQbyNa8ZXn5Lg1Pqza/ns7xgFUWvweijP0BiczGTkrydpGNj6ssxaEQ91HloudT49MGPYf
GhFdPvGtKCKqOnDXW14bR86L02CAN/5ZB8pZs/RwH6xtOtyaq7S1Hv45DPi+bFnsNIHGtnk9I2dc
NLYzQOpzAcMk+cekoR+A9Nf4MReITC9tpO6GMpZcAyD/LXMh1mpbxKYtsGdNO0HzknyuB0nmYYTt
1nU0j/zZaQ8qGUGeDo/YYROsTU4wBh6m2Zl0xQhH88VTluA/AYDa0NDTEJanmyofXIQZqtFctNlH
fUk/MTHz39zuAn1mBnzS5VL2IlpJJz9KpQnBGj6cqJpbvvHg2toAipVFEN/us7kP7BS6ybNckGSJ
aWfzEW051y1cTzkErsZZbtFw89xvkUrr1ZOPCKezekP3tT6WGkco+x1XWQfqlcOo7aqpB8KKgftd
ZL/oeF/F4p1wlI5fQkKzve00zmxaRPrmPru+ze4vBcVoTPXLnqv1KyLTmOyulyMlUPj4QXZ7846E
OxWLlRbKDLk3Kq8dirZutZQW0YSBNxpbLIbqcXn5VkFCblpFPSALaoPYqV6kwLU57U4qevaO0174
5NLt3bdC9DrR47OQif9dfkdupI0YLW8QCZC/wa5sr1GGzwNtNJU/PLmJ1EIva2XwmvLfWkRz1xRv
H0bBJ3lWHaH4OrbiaVgL3KLTtvRBubS7BpPV4+UYYuVDiN/PJ6mazJvdp1OpZy7hCjQL0TMQp0UD
RW5fTNQ0qcqXGb/vriafZzkKaj5Dzlf30oJdRLAD3D4fzhDDVSJvAwOo/VCmQT+JirG9KHPDLgsO
FxfiL6ZUCaQYa+BqckKCJl8KO3s7muKqTOhwTDKDhxPmEGM49GF/DxjufneqOjGkgIXL8AEuanGx
t/CEbJFW3L2bJ9VOW0wd/6NMynYR5QgDWhVLkMjcpbKvKGSx7xgV01jiQosbQreRzqgkwx7NDrNz
GJzubRHZMLZpZx+o9LU12+EJKIJHekAw+rAuQcqSBiW93vhKvCYqB90IGbu+9OVmo6C//gZch5J8
MyLI0YVIXHKUjdy+JcH8opXo7rCtZ5+3D0wUtqeiGqf/6pbJC/kpTKg0SrDiiXrcl0J7pQAjtbkw
6HNBXegHZM6nM3da4T0P4OCIGPmSI5fxEw4UdzVmOnGxBSsO2KmffvCNbe6RIsd3XxJQLItqEMCv
qQJWULlqjR50Ytbngtp+TW7dwLMGRMXn6GyIOCaC1rH00lACYoxUrkZhq4WSz+mM0vQuH38hAxxY
KdSR8P40fviDFLbEsCDb0yWr2alCK39p+OALvR9bsu9m87s0jozoX2/L8voeHYS9S4/FM1RvKnS3
48yVCQ9FZzL1sx6gkzl4aAYe61JT+4J280mXZIsB0xkBpEC0vNTZp15RTTQTqQLiIkcmdunuYvUU
9O0sSlN4Brhjw/n4kkJexSF4fPjfAV648GvyLKMB5NbUzTVzX80xV9ZET7+vPoDFVycMOhSx0EJY
dajdEA6CdmK/5B1eBKXVcOshv6kF7QlAXMt8DIj7khLgG0e9O93E+Lc3nBFzR1gIZq+chwVsg72K
GGpXs5NOx4Jv/6LUH7135hxOby8A8FuwqnNOv1EXeXY3Go9ptaEFQAR1DFqmLz51VmlhFIsC67LN
oBBTPvrGdfoMIsYyNcIiHLZnhtmVCEOMc/oW5b0GCCzwLhIcfNDJhyO2YyNHS4e7Oc7LPPadlff0
IaB3zewL2YLil2pUqVidtmQrg3H12wo1voDNIf/DaywyreN1VNz3UW30V1erFZKHJ8LcmRDx1U1I
fs8byJurn/LmYdMDuAEBZ8RR+veUJMMFMf+Fh7PoTz64ijdkcF+3g8welOfqC1NkGVCS5X/M6sZ8
URw+eThizkrS10YCrAGZF033wd+zIr8Y1kYkEcj0ZwjzTufZK53peMggiMIr29Zph09J07w0kLyL
w6iAfLMBAl1bzTL/mpvSDp8PnbcQhLCnv7P40OX7C1gVRRcbVMgMYZ62qshXQ3Bjx4ifsy+uWAOh
jUtLgY/sTVPwEpD1WdbakQPwaMfr9MS17mHcxDMj7slrRjfMG60Ut4f19Bm39eRDIlz0C3Ab9jFz
wafoBhSEi3a/x37T2ThUxPrmLqPqi9qZVFC/F7rHqRfESo3UQXqfTqtePw3/2gVgSWGLGCvzq15R
kj4QdC0vVMKIQ5OlfwZILrK1yjJSY4qn326CY3JGKbgneEpE+DkNFIYmATQYgGFaC44mVW1caRy/
+BLcdC9wL/ktwfEdiV/L0PdDmJbSkrQemnpQb50i4bDgCInnhbKUb89vLupcm4wmi5gI85aaN6qO
KNOqLrQtNEE8bH/waBwgl1tuW3ROGfDpyPMx5cefEDzfsGB09nnxRsekv0uJC6RISPZ2ujDo3Oc6
vne7zaKvgfanYTiA++pSPM0Si4dGR3UHZPkVgBG8Y33NHbG9JjUCQc2Qn5zRx8ngREw6pitS1/rn
1gfo1G/aBSC5kndvOIkZimtf4464OX7ADvU3DexwsyOpCiLA0BlBbo/+heNHuBRBqqWEK8HQ7apl
4kdSRdlE1RaWdIzL1QTS030bSYaj8zq6pE6iiQ5gLuzNnR8qsVBf98RxSQm+XrWMRxt5VHGioQFk
5mHFWKZ/Sw+QPzeW7p/kt/eSG1OjtLSXWtUzY4nC9KrF1GNit3FMTGk0KKXt6lm3I0+a3A+JS0SG
edrINDZDRNWcjq8Yt7Rz8tleTdQUfWMNpXpuzxJhSU6Ppo77h2u2RPT8mi7wJmmuHCh/sICXpidx
NzQf6u9WOgfynoD9+UZaQS53GquOm0Rb+nt7yXbczESNpDxqiRni0v32c3NzBofWyzPFOCWxI8+K
wrKPAZawGLgN3eJ5LJjMVSQAp/NG/OZMfyq4CbRG65t+tDCiYRqIXv3+EuZutdqMUQEXMDKtXyWC
338XkJUfdoZZgCma3d0Lkj1cQZXax+MdUCuLzVFaLe+q1cV9A8pc4i+MdQkAUTypwqO7J1w6qlr7
a73DediSkSMMWSU7C/MUDuEi3+mRMN0W6Cfp8z0KPlh6q3UBgXtRWo8Zc7EX5dG68Q1d4BSjrYmm
vFH3lD03omr008CbzURds0EfjECdHNbPV2Y2vukIkxsqUlbzig3HPNZczaYT4X2ZRJk05ltXd550
Lb0z1nssCsRBgbYb97uP8Cl4o+066vw3uH7c0YO5o2kLcIxXEb46F7USZfV4IvWaH9YyOPRx7Vee
s5W5vY0k+Qjad5JvQVqySZtx19DYnNRqD0tvh+ocT8JHL+S9LZDWvIrN5mZwrO02PqVngMjGKumL
YfbI+fwrcZGfv7n6GQ9Tiv2SRrR9YyLpBZEvZ1X3FwoN/nYDpY7rT21deg+OHWuCPl3I57kkuWX4
DPCW3FVsVnPHt3yH/72kSe1Y8R5Uv367zRVSH8sxYDfIhgwr7wecfT0R1uP0HTRSYrN5O6qSy07W
L03q6g7m9DcCPRCnr/tx3Ga1RupyjOwFW2mt2i2tXw5GNUhpE9opBkJwd5asw8DpTbXeYcMweKbP
FSx0/YymUFODtiedIFipRIa0EKGjA/drhL/oq3OW2Pj7zO33mE/STPpDn8vjY+ZgILbrr1RXvQuU
6VZAo2nQSD34pSBNDKyTfKidbPpV/2g2ajFdPOlVvrDs5OF/uzBrpo7rR76imIoidNX8T/Rbtdle
2VgpMjuY140ThTruERK/cYg/z2TLj6Pmv+lqOsbEKW66CUYNLwCsr+XLXUr4qYjwEiluJkiYmXhT
ZFEuseCarwhzArL+TdS6PgylYmL2DF5U1pM/yjWrxXQGYzWQiQbdqT9CJdlkysx6c4XIEuVtq4JV
YydU4FeCqXK+JCRzbtT6ev0bsB8TMJFgMmXRyeWhEd6X2yEHCM/kpHVr/rrF0vAP/iR3VODhieBc
tJLMyW1RPpkWLXwXLmm8ce37QyRkjgsLBtKuxzbC4S+tg6+xyxDso8EtZnes6nT+YV2Jdfu1RWMd
ulHCmEtQLsp7i9Jrh/8CyXoN0tjFWlJptnlVCHxk+UhP2bU7r1IPC/p6j3Fiqf7yttXrcNI2ugYG
m3o0zrnmC39xPgB3N2rULdrG+v8h/lrp16yZk3YjN4HrMExVAQw4GjCqqVJVbGz/dKO2Bvn3vAdE
ujjtWYg0Ne0PG3ppC76yE0JlXVi7qu5RKUnbBfZwu098RzMS+6fp9YxWiQUl1AVaowInFArOUCR9
D8LLHkOFxOr42LqlqNnZX5szoAYWbI4HkJtoIEDLR6pwDuT+7n7DY8q1Z7O0Z8ERWF+/Wwx1sfrF
O1+/TIAO1vVV1JcQ6PkZGEU4T28+FSrUZ0Cf0oCVOaoG8xweymUdTMtTpFGveXxbuexPYmK36lpV
9erVK+ePo7ub8Rd79Eb99FTYZdzK5YllcbcCWD3LgwSDHJKAuY8lE5FDAvRPZSJHMvbSj/7ofCqT
3zwXKdxJ8szbVscuDFSTrwgxAq9tjlPkAXyBRJj8XipCxScIPos1vi8qLnWbj3UxFmdq07yhT3IX
BnirNSyjJ1iXE8QrWyBz6RJ6/VHbg8HKQ9qoaSQw22ZzHUZuaDT3y60PvUHQ/3c9b0oPMORh+s8n
r7HyArXEm6mj/IbBMQtLApmU1WseVxHbPW8stTD9t7QngJBGLhwwipXzukqiifNOAJOefeSCxfzl
xZkJVO/EoGlIIjiK70xxl7r60jm4Hs/oHCGs95Rq63Q/Yot7TNVesxyzTeSG6wa684i87JQWeLIE
IY0W+Ftowcu/cHIP3tCacLwm9r+pPoeF5I4TowQtitXJLD+ZM4oyw+PWItNwnc3ChEIj98HS2Obj
CS7jS7/s/sBJcGUwqz0sQhYgd+rLlosI7xD9Kb07gCWaaEVXPBVUisb+G8SwRj8aopDNqRX0MT0U
EZZKwvdX2GoE3bQoGyN/CLUbsdObsl9zP2GdPa6Olfx3fynzOGWGL2/CAvUJxEIs8la4YRbrmI2A
Z2i2MjoU7ObMCm281QA/Szj4oVD2T9TDuBpuVw/cZJz96I2uMap31F76/YFxwEIJqew8lWk7M5U2
JxM/4tel7Fef+GWbX+zTlwxv9PUXlrh9WTSqLhkTjrAKUmGEVG0igdBvo1ZHZVh1xztMD6Tk3aJQ
DG3ZJqaCOtyhZvIM/jHvfuI1Rab5Y9IU4rBvQc8ay10tEmch/PSuXNiun8v/0zQs9yKWxebdxNL6
v2qbEHUha5Fh2KIRMpYoAfFOJIbamyOjs60oufIqmsexk08Dz7Zkt2Y8xtadyd19+LVI0gca2vnl
ezir8J2X6JYpI+2phnPZ+dn21InT3cVMgidg0trZZqXM7rfSNaiOZfq/tE+99gQ9I56AnbBvcuCF
0XV22vjG73FxkjL4142wVMgtmf4RFAL+sHPgoVhWPk3lk4YStoA4iW6evXsxMckdVylWNQ2q6VgQ
JK+Cnqvn39HBzSQIZBdqTB0GHNGrxwaWyut04WmoTjb25Ee0AJlLgBkTKSJAcqs53YcED8tfUZrk
wVYt3L+i4KVsLjG7GijxHau5gGJBjmchIsc7k1tLkpUjIDjLkr46v9U1wgDMjq6YdFT/Xw8z1db2
qCkRNm4d0kMIzxApb+a47fzGeEc5/BSCdD7rHaDMlOlWesu3ZoMeBxIawBMUQPBbdVeJL0v7mcLB
skEihsdCjGq8qEeFVIjh1zL53nLF23lzR5HYPK0uMP1TRVRPnb6afrd8mo9S/ytT+kFlRkFO0OGx
oKsEnSiN7eJ/4oNv8OY4bmt6tmCwILESho0rv8et1VkmpQijtFgiBNxwlF/nHtsxlvCGHZkXTsXg
Y8QrPAwRHEbt0CREOfG8iZIK7BtmKvQxbeaQaYJczvgAAXYvLYfBzIIhbGcP4lY+uVLRv5ddqU1e
gF+jsdD1qVWhqcjwSv84puD4LsWyBKDforKjMMk2MJfsvAzkgjsOmLISsF7KzuzD/Np+aLS5pmw9
VaQXEvqact38A2kAzOinICFupm5tF8R536VD7dETLRLGWSt+L3WyNc/HHQDPvc92v2uLziEHFdat
pytrrcDOPs7PJu7vsaM759+smulW9x5CJ8hv7GTBdD4gKSmQ87m0w0GI2O6H2ngVSsIxp6MeF95p
QMFGmAhYZkzbJVOa/fup7A7uPrhQMPzp+/juQU9PVRdQFx73cfYwGpw2rPkOk+anmHFNXHNi8eNs
ELUtHaBXcJLsXP3rBVsF2R1wMgNfFsqDVBQxuRTNQMq8BvUtiMcDXz6AcmwtKE9zYoJAHiqkfJjH
vU8We7C1CPMBGRbaipL2wMdnxYOOhLR65FrinbF6cOMAOGPnRXBpYIGbHeFpgAY17W6pbacyRzxY
KAqst28oGcYAva24Fld0mgZrmk8KtYrYgl1sNipNa9CFGLC0W2u8bRlT3S/nLoL5hoDWw3GxI264
n6iNyFlovPCGPu5rI7eagMJa84P6LIin6GAtsZqETJ9sQ/ef4X/NPNjoVaGb/hm6dMzJzU17DOyJ
R40Qfkb67ZF8Uw4Y0c5eqDQaDvSEg8EyiOZQ8Rftq6AyUVfH0mIwxUHMWCJ16ZFm9r59NOoZ2oLV
nu7anXaz0EZvSPkxD0y8V5OKMT6taBOeVB4Qb6fLG5oG68/NshHPIWtFA0u56qBrW0tZbHP5FmEL
6NYtf2VduPDg7Isp6Uwao7RN1psInmdtba+2xSU1DLfLb00orR792NI+f8jl1B+O12xw0A053Vku
mnVBFk4UfIJhJ1cB49TMS4MFwskW1hli+jtAUIVgM9K0xwhdEZ34rti5cB4DrD42AIyVDKf9FzhL
mAF0Vi4AbIfUwyRRPiFr6Ot3jas4BLFiLBAe42/lA6iVFeAQSh0jeAkjG7GSwCzBE3HNNWQBvd0j
u14e7yRQro3e03OUkkJMZUufhiBHLqIt+O+n1NM+8tfLcmSxo/IS82vyZnhWIIjTlFZFd+69zlhg
ERtboyQRn2Wvu/x1F55zdMsjTecwe1Ntw+4zAn6YLE6FjECG+KfcuVWLLkgyacAAd1nUGD0/UIjO
dFFJqweTY4+cL8X7RlagnJpW69SYP+uoiVS8R0GCvxHy9vLhgFW9zySDU3GZTxhKVeTMhQBbHN0h
WHvV8cOm1rvdimNZlO6XC74iSf1sNaz1jqbcXI6LPm7zQM4R/SGsIU8H2UgELDJdQvw2TkEEPBmt
Di4wKgi8CdmInj3gavMrrEiauxLn+luzyMD6lmxGe+53yWf8eurN5OQhE9wdp+7bsc1Fy5WJGwT4
Kx0kU0KTeEJ+xDiUJmGug6M2yCaqvTnCPw4JE3HtMQWVqDGdhTv3YoRQDLmsAS72Gy1uKGjXI1Kx
qG/dX9JW4PjHGwlL4i5fJhUIgxR1/lb+MWHD3pVAJavslPpguT/svqrmY/wIPC7ylA+ciLmB2gLq
kHPcSHa6fthf9dNSA6DNGb1CtYkXcfXX61rQJcuvjnB2ikCL6cWZ1zKYUXx+FxyPy9b0wUDTJzuY
g3pUDnORS5uppQUxMtnJDqLFSFJu7d64NR+VAxOJCrI5vzVBDYw/EPPtzuvmbBL9dMgu+sFFO7Ii
LosJx5kopoxEDOAX8Xm5ZNjCPZxa6PjkRsrv+v54S++Sk+Z/Juga1XBkHGv2AgpzhU6vNjuqJx88
pWDarDJgLVTq0Sy5F55ic68WtL5VDw/42RQM2LPKKMEIcUbojHxGoEc/GzimSh9bxMc8IfTB1nym
J6V3uQj3jQIt54cEumsm3XwHgWrgE4sdl40Cfxy3nyLL9BcmDA8nxmqGKSWY2rPVT4Yz3Zizdi8c
F/qD/Vn7vjb8J8taRGJqWfxTlcx65x0u90RmarWPT8IB2yLWi27ccGTjthMdgaKOSDXayUWpoLoj
FpM2CagP6i6WMdQEvTLn2pnVx7hZiiLSy5T0GDZ6/HNKeKkVIfDoqU9XhADiKjXyQIXj02+lwsqW
9f//GiZd5XW+YUdiAu/RHJTmx9WPQIWWj6ON8D7jjDQUox3E/Zm9lbRy2izRMwVjIqiOQ/QLQWig
5LTtTsJjyzJtCrVWxod66YkIOptP+h8EbwoH4EY51cp3Z7cQ8TzyDKQ6dv9iul2DXaqj/B0+xn0K
PQBeBml3aXkry+i/1cnmEBQc1KFlUXeYwS2gSiIKjAFmjuNQd5thz5zkdJY9Rc85olL5pptyj9q6
fCfPgOaZIjMU8TbAbQwsA6Dh6lWZUw9ou4KasMW4dQs9bUrwE1S+ueqaWCmNIv/wNmgO6GqTVslm
5GP4+zaAwh6kdfQYEtq8kvFU848lUZ51Hrly1keOvcd6fnrxC0aoL0mP6P50ojqcXzJzMJ9HeQyM
MsTLOYk8FGTxxtSbIQmYgqosmJyuXE/KHnc4LOuFrwfQUInmVJ47jdPooe7bJH/fdq1AwBfNF01z
boCVyWkbeztCzN5xe2cCk3BAdfgOgnOjd1k/uk/t6yAk7Kj+RDR32Q+p1jYKyMBnHvJdjNXxFBWq
wIeMO6bihZjY96ARhcSh1JqI+2iNa9nDo5OO39p9z75abtSwBX8hKKeWTJObDbbbb9kF5alPapnW
XokoJKQwYe89dwJIJH6XtfyV/767uhBcblLS8pjY+4HH0BkUnWgtmSKgPZTJ1Ec1g+F0jrqodU/3
1w39rmAW85bZLX2HC6Li0d7ltWuKIP7o1xmOQZn/f67yUvQcuR9iiDWa7E48DVM46O0CKG+ew60A
qV17iuKTOc/ds8iCq0X9nFI/1sZY0HyiwqE01/c7M6DuC+zA1FY/rocRTZh9oMnj0DqQ+sKk3fYt
w143/q5d50uRYfc2XEjKybmrmOGj5DqOrdjrEnrVqqENuOmyFlZ6gxLtnbkUomupgFUJoE4VKAlt
71yBfX85RVpWN0+dfZ/HnNy9Bmy4Gza/1NSyfUPqOMOMeolgNokT+0NQ/FLIHcUJTRgx0XVIWzEh
V7uGAGe2nf8E3eJrnw++BrxsY1vVBS+nFVrswoY7kz09PoJvpF2h3zN59dA9DFLW54T5nOTkyZFU
LXBkvTJ54LOwZxIp2Ib/aSuHNcqj1AwMWta4/Za/gZQXVZxdfJxfC7+lJy4kajrzIR3XedtVf9s4
KAvN3v9Tjq2gnc+K9CqCic8i9uZdgwK9xsEpuUmtQXHCYgKp5ZVBVyWLWgyt3sLT1lJDuY3Jt9Hn
gN4uGVDQTTQmUJNUiTWNOsnOHXOgNBJuEJPryRfTuO1vRkwWZ1k8uh7nkz3LFOiclOBeAyERH3x8
LQR/G7y5+m9nWFUGEM57/OWyVGXeYEgn82xvlHWLw8C3Filb59n21YovZy7n/Ng6AT2aK48ovMT4
gflDsxs/BBDSpFDHrnVr3VYtDbYjFb9FuFTCEJu44EVauOJbBMTpkoCSbAiMmlbt79aGy5tCJOni
sPquZI/HMdn6VN9R3Q30UWqkaJYHF2TumRd/l2jvyDekjLM/Rhey2uSpDIKspP8mJhEjH9uG4Zxo
WO0T+lHLWLzsGAqvHA2S6bRihWvvPScUFe8X2ZfBI/c0q+bfFloTQac6lhZNCqz7v9b9hYfDb3kW
Km7ebSEaslr3lFSeaTY3RbjC7LUJRzuiIGdXRDV2r7Da7KUJoZi/MA11IL/AWOwr+40kPPd+3xSs
pTPxqcgwmuiQlGKk545Bro9CeGsNLiHTb6UkJaHHGYHmD+Pu5CzxGyCNsmRS+0bbHhT4SRXtM3j/
dts1m1CU6izHxZDjAOwc8yRpjkzLgXHJjVLkowa1VvkBCyWn5BEGDY8kYNpX1or1/3karRIYwixn
EG4dQQkIs3pJdnfE91CwuXeWFKKz91Q3AHBrjTUTDRNTOWlibzFe216p9uUVPb1FBJzG2HXw1i/k
HbHiovPQiIpOKEiA/ZkJV7mJnWO37ovMYNTskkOkbrfjeISARSYTvlZJNOI0MP+gLVVpCTscXW8C
gSOmBwCMP/NKBKlIH1GoAGASNtq05iHtEjeunA+vNiIgAzVvmfnqk/HPMq2DYw4kj+FC5gZgsm4R
IKPPAoIlBKeV2wJ0w6cli1pm1xhx+JvQBZRQBG3/Ehn5NdcEQyrpSnZBGhO83CGeXcl/5YEuUSml
M2dr5pcN9FlqtrhP3eL0KlNkYEhtOSsKwcNbHk+aWNa8TVn5eo4EARz+JUrV+6y7PGUCjno37pG5
h3KnYoHeh9HIeeG3jLXznojBTmS8xCKQ4/8yGJRZc8mrvFC75DUzzRK+SqsYL5Y6qN5Iag4Fj+Iq
Jd0xLgdzGqX2Fkbw51wGpj2aAR+xNuFynN2kX2io4hoC11n/eBXCOzdU4E+GERg++btbiBbMs4jq
0KHLS0OCQLgOteZSTl8IHbi1Ebrs0a3oyVMSNSVGP/BLIJSur+Ol3awZuSKrWHk5q+BCjPJ6UPg8
AIZeNOxqmL+PvlP4Kctewfwkik+VZs2IpzZaYxLl8aOD5xiZ8PglWvaEjLtw+PRKb1jKL7bhQnPd
I8Y7Tq0ZTOUnbSLFgxNymEKPymGfP82rOmtL2REL8R0nyJ7aFKvyGS+UdSc6dJoNrY2QZFfXlBm+
+wq539PIXLHITwH3P1LoVhABmF+vkohz2/Wih7V7eSK6BBAwADcFWhwTuhWn8FS+UaYjQNqqatYl
uj7/MCl/LoupqLZpCeLncHp282DCutxE9uNRpucN4EgpHHmhPK/QqsUQ+yGS1hl7VXH0XzHPEarG
y6oEkEznueTN482JcTZ/v8XUd81bxiXSozdR0pGSXscAYsBY4NtFb60mrY3OL8VdGmpjc/AOXblu
f4A5hhHPTu+xavDWbwvkoXoeB+u5ZWWWblyGjcIdEr1iQhe3IkGLQ/wLbDfi6ojZQmdP2XBjBt61
r1DPrgh4S/nitJx5reinfv8GAoDnSNzj5e5yYBpqXqtbuAOefsPyz9lRFWb6VUXCcHWBOQkVbeBG
SMtDBRcv3tr4dozSf8UZ9cz6X5iYz6SFEsicnbeCqqEi9NIRUd1MXQquNrgzhaNR9/nHAk37GCdI
I/VYCTxWRvh5/pBUZNLMoDZssQeK32VNBKylpZ8MuJ7TpKU5vSbosJdSjN/VMaQQMz3HHFtpP0LI
Huk9vklK9Cdp4MgVQb4s1sMeZ82u37mm8geCeZ4RU7Ht+eQtn/j/3xHp9R3N/kqyopXuTh78vn4D
F/ewVvMpViAoq9CseRk+5zDuTeSNddkKzUKiOYQjAr4mJGjO3nks1S4y0QdLrDlyIpmgReQj76+e
usNCCwdRsdPVZF1yBQAqZmcJi2RU4UfZwtKsYlFKrkf3U+MMecOhcGPitAmGtSACKSDDLNEcU/Ku
ludcBLGwp6xqi3wa9EtAo4QieaxNZI/ml7q7GurELyPk6A4QG2d4Wj9KW4QrCkvm8PJ5JXHaN+PI
f32EJTtGlDufhTF4zIiiOYQ8rm7Jllox4L2KnKq90wz5wQJJ+Kr4P9vcVIwdgODfZ0GCcXutUbIy
Kp1AtRb6omVPv9lb48bCFwLq8iqKhhqbqay0+2tqeT3Y+iJ9LPaiZjjLAJdgediRsD5ATEN1y2S+
8oC80sxbr2Z3lE+uZH8Q1r6REMpzdxehkiC0ALbfoAfmvUl2UkiNx/5N0ujMG4qEkmVsNlRS9Kog
lqQSSoKI6uPfbAEJ3II+cCiUpyUVJSZdzFIrmkYWTNPOXJQ2J007VQ6FdyoODPRbwo7JSj/HbrHx
KloE+IPFPcdBsw7uzQeT4hF+PMqkvzf/+CvbH/67mX37oSl2ko7aeJ6eU5q3fLI1LwjL18s12Ncc
bNm42WinhwoFy9ceSNPOS+0pX1/3fTEacWdcT+YiAVnvCr0iEfMg4SHB1Vd9IZAOlkxnbbJsVz/g
ofg3QDZ1dRcg27IwmuMqu63FoWEZUXbyLmSRaqnpVh+7r2SYaQs14RanNPd5b6FuRSw69HZtuw4y
PJOyjeSCWs6PQTEjM8qt44flU/wL4mYV+0qGdqRJKTnU4AO4LYhMPDmtZzv04dpUXuuE6np7Pz6p
7tjFKfgX+Bg+vtC/YqyXRUY08PKByCXlKYg/6hbdgQHzJglH/GgCQ0p/M0T74T5uCh95w61Q8/T2
iH4Mu+DG1+bX5rIdMhmylhpCAcKjnDMXdDCjtlf6Iv2e4xnMRrYlj2JpD4TZpgk9pqPXSYylSNaw
lwzc1OZypYighOJ59SRVEwkvsO3m88XwVK3qYJV5Z8gew0DdXcEKyUdd5SUjR//udL964VDGhQoK
rKKnD1Xc0N9AevLHQU9WuXb/7oM1bDVzTFr/T2CGxSi/oZdqkn8vEEeIbpwKqhiqmCJ4QcOmCuIM
wpP4+euRLnFC/xQ8Vv43qn2A1EJKm0wEHSmtm0fL/hbldgG78V2RpsomyopP22bWFY2Bi8GSWxJ1
ZDXbTdDLLF2TOoR4UewmJGZXzLKSMKdNZsm1rzIbgCwlM/J5dWMqgtQbRICsnuDEMnAioYK2hi7B
g3ZRqWqNfcwl2KBIGDhxj53/TmQL2+tpg/CXSUMb67Ot+3xUBiUJU/KEwYzBJBiiPdUMFRBULO8n
wXAzTVilfXwuvxwoIIB6PwmrF/32gHbpbPuqmEBfhlPitJhhv4YzmC6+QpePq7YamG4NQu2D6ZeW
yWj0LGeTrbCiq4kDvJCFPrAm4BlYxfI4gLPv2enUYXaQPjmrC56bv6lUaVRYV3owT8FSjjkjl5sj
yhXewGSiCDT/IVZZj7F9wDhdNo4/bZIvrUxMjETWNPHg21/8UcgzawPFzCuux1lQL0tpC89tAFH8
0E5U64x/CBzjVBbqtMRtlgdOgQr5TwJxY8HxZHkw1nMrF5ZFRIBFc1u3RxwNMbODkpohTe2f+TVX
Zz0djLVZVLJ+qAnbMgONP5DWw5IntFkTenrDR0KrKqFstKCIhBPsuzqnkCjxRpMOF6d7WCJPxUI/
F0lOgPCUj9PGyDfTyz/li0duOjoRamOgPdYdguVkHlUcVmPzKIiRlrzVKO4vLln75/hZAQmhfUN9
gTzGJjsNwfJm64jsE/ocd/iMQ9AnfDN+69acKsmaIaZF/K9b6VhRB9KYlzNoysE95MKmlLxuxlpV
6zbtC+7Tw9Ucs+aNCOAUQaeZ6d4ItTOeLBYZqRj2GicpW4ccr9x5VAAGixvL2nbKTpxtHogXdv2o
zzs81HbsQsNyFz/Lrsl6Sgo0OGgfcGqF6uV9Y3csdQnOCIHLLL3SYy9X3z97zgEU2E3wSIMlgaDD
/4DALkoWhjWhcwBSaBZxxLfzToCcz5ghVPcL1M0RIL1fay7rt5w8esCrx+9RumZ71pJdhThzzxUj
SjLYqMq3Y2nb308J7Z1JL43ftk397LINzNGuKVKe1T+9970Hwh1X/BFWwVTQWhFy07FoDhUwZLst
tsTCSCmlPZvhSkSa2HuJM4kAeuQBMHLjoQMmUldcMNP9Ju1PyRm4L1SG7yMft0d8U6OwKcNoU7/u
RJaYShs7jnM3Q7VAWnLtEZK7sMzrlr8v5rwvlO5pWkx8YPDoDb84pgb5f6Gfw2x4ycmXLEGmk3QB
lkx0YEDe98z9IVLofOPjPvNtCyHYI2un0SokombfU+15O59att0xlZL8g/FDpT9dl2dFaZrO9JEq
M8ldTdbV2QnXV1WCZDrwJJIlLj198MkGTEeZP4Otra8A0wjMz+woUNumBbwXLFbmw7evG4Ucl/vK
Jl/rxqNvMxFP6Alh+drPiIS1/q7cQ0ZjPc9RdQsYPZ15wWcvbj33k3qKPivxNly2ufAoicFYrIUN
6HgGoJiFpYmcTdtdAxr8IpwFT9UHb7x4zmM12bOk+qQcK4xtiQs5yp6mdI5K4gQisfuJ1bY/CU3m
33979e5n4arAkdk7eO7PAMRmt03/8IdedC/7F44WP+9jXsZe2N2gaGAC0hry4gqXv3Bh9qoaDAXH
5cgV6b9hEW3R6KqiW4KdQz/TZAZaygNau31mQGdhJXCx7q9p89eo1cBDtxbD3G+gzg4K9GIVSlAj
itYMf858p+Xto9NU7Z4wqhmEBbzThywc7ZvcWV1lZJiU/PHOfAUorc6rkndiLeLTksdBfaL0Lapx
P4vx0MOmOnhWvEgQ83xsZZd4PzVf0SMmCZZoMX21U0JYuG53pUgvEhqSz7D2Vmji+XqKjvB0fG97
XUnloQCq5tkNG9kd/nV5/qajVLPnXEKTbXvCRyapnkYYy6vfYeosGUuKd+zG0uSwFYUqfnbht7AX
gaW8z6YrcS9aDR7PjaJddXsku4/x/X88rAD2nLeUS6fn0O30db0vuR/IYZoydY+RsJFEl5ohSlKU
pF7vmk368SPzmFVivz4SJ8yCAqdtOnwgSfPQ8D/LUIl7uRYkH3ReVWHDdWjX50ni9MLN0gi5TqXK
stDlT4hBBPrk941WjdA8px5q1SrhrXKrgiBE+HqaWtjeG++m2T0x3hRb+E2I1Fa6FMkNVgAaz9TR
tinNvArwo1PlNXWg6tN0/wH5zI+K9vrqPgDJQ8sfSJW8NtjoZH/CQwjFJr5wmLydTU1ACdkx0VsE
15ZaQC1rk66gulbn/OuMnuiEcDf1kL8yTWbzI5zAAKs35ge/C88UesPAMTZF4FIlJ5FSfzIoBynX
2YG5efYKBNWHT5ifTpRHaE0HOpOhvW6KJsq4GadbZ7wdS84pwxQWfwRiFaqZLa8HLR9dbxedhzpD
2qNcxlQHDQ1cVI81dWKrYP7q+H201Dil42ym3pPYmq0Pormh9RgeXlRL60/rYYno7Ij3o0RXw2Eh
HuoFarbmh9cFxzsDEzQIdpDiCDDwwaxU9EIW6wQEjGqZa0talBzAK9zE/s91IojbXu/xcAtL4AME
NU9MhvdwIoX/ZbL+7pRSjj4Qh99hsnWXYXcwA+shncTnJ1YH/g1NBM12TIBh2OrAhDNKVXPG2e68
ui1+rbd1FstDj8tqXiFl7qHkgAms1cHDxSa/iXndeEKdPOTI1mUXAOyIa+jmjrxx6rI4uqCeDG6p
Zs3w+3dqPzrpVydwoouL2dR8q176oapTcDTjU4CsjBR1rFpx53bxtmGEfUbPMRaQiiSZ6+rnPM1z
+I9rmJs1mkLcThdCnBKsm3vdxoSyEyj0c1j3jxjk0rkbhwNkUPsEIx4FXKxv02oGmWaTXCK6nAut
9dCqYSUyXucUa0m93UxD9juSBiJ6/l+sfYAfEKohAGQuGeYlViwutjBYNO6izI/BG6+3dLDU+JiD
1HfgaaysJJufEX7C8uCsXx8yFaCTWAFldAzo17ooUvH9MH38L2LLneHUIje/fevrTQdqRZLoEqOC
nlzWBgkkAOGq2TzHnyrddU1hAetP3HCJS1gTK8I3ZDvxkg0jDNNrNzZ0YG4CYz5lLTV1VAJZ9Ezn
IzcAOtOCyk1j6nKRSLtUhvpXGPvr8s/LcIw9zNc2HlCu08hEYbbkvFY6shCF8kzJqqD8Xkid5LdM
XqTXtXyBojXnObChQrZP+p5Y5RGydHcRdLJGpQ3e6PYTaXHk6b7Gd89F1GvPPDSZK834yXYSdkBi
nhXIC7LUlcUwntSgoGlyv84DjyUYsG91clEBniCIOHYo8kgXffePkJDSKK5ogRjcH3bdGnvLLnnr
JpXnWE6gBS7g30FBX8MiyrWX2uAAopmxl5RKSkeTEpFyrM++iIXrQOAvRBk6VOvDT2WFV3sV3tPS
ztdQtlsQ7NpWl1yS0lQMaRbENRUkVE31rQj53xmayDDCnflIFBRYHWb2IkiJMW5CIZLhkRJ8TaNH
npj+OrnFIVdAjrPhh6Hoybw9JOCJV0vBsjQY2CJhdmWmLq9zCGjy1CUO1OSd4RtDfWdZOzQNoqfI
UkfS6WS74B8ni6lZ9NQiMXtywy8nSz0KkZqVHHnye475F/3VmrlEUWuN6Bn5TjDLzd8C4ijHmkyv
IsUNW4JJcIneQuGqph/Os5wWo2fMD9VKMkHkHbfe5O2GyJOPbjHMyVO/RKMzledQqDcBiAGc+7Be
aecL3qzPVyM8R88UVzfYMXW1RMMlNxssx8eeEdlSGZPe1rnxo9AZaETKuW3HRZRHJjYPu+uKODnq
N6p9sxSIFUyulEhJjYI6Sa26LQOszxRh9MUCCVpNbhAVrH0sMNvWo175Z5O2kJw+QLbAjbwa8y0Q
9Nky+ZyA35uEAGftgezAmo/M0DQCfhTUjM76PPYk2jUGvoigo9wW1luD/daje6Rhd9JluEDObncz
QXGUfqLaHg0KatfSYCcOSX+Kr/my5Sl+1XqmrozDUgdMsfHUQ1KhbHsh9QAgubKVOCDWlbaZA+Mc
QmXN8kVSFLI6TklDZL3VVa4NlNb5Mkm0w2QeV0QS5w5ZEnSxTAVYDWq9ttiMpWlsP0lxamTE4wKs
lY/LPRt19mBoUXrGCq4Iox8BugONa2oKvyrK9qWQr0pGEAdra0qUxdT0hOcTFpPqNz+7Z50guWcY
yzhE614SKfD2F4ZDxr2taV8yHIHiYFhJ/Mvtl1XlhMLtjZ84Ho1RVXQys9JvVf2loT5ua0SfOiEq
IvweN1jmIDQZ3lrYD79yVhPZ9dr6vNqVONO3qXeTGiyUE6FqkyG9EWCH9wY+hqThhnZ1AW/4krMr
wlupW+btHBO7oTWGCXjnLOeVrRXyz64YRKp0iQocvWSm+aIP8a/grBnaxEuhmk1pRO4fe6MjAax2
cB6mWNjFwWd8JHsU/lDXEjWVacqJItYECLfadnW065S2PuMwV3xoJlfCdIV2antvVPbIPPjQfajZ
3MAvftKlSsGC37xyY/gTXJcnVKgwzvd7w7MRSGQGGZvJCQlBwv7QnSxRvWLVpMaoecfwXZSwG5P5
E4DYYXGF8dDs+KRGE5wVIH/zG39ECqPyJjLy6UqxTlbWb8YTVpsqZ7XxV9Td3lpLb+2x8urQYdfA
v6LZNx/G40wZxXUNkaUSUKCJJQvKioe6IJuiFgoCuDURKi4CCLRaGMsrFmu9+GkDwnQtGdUIhDIb
wdydPWwc9KMV8E97BR/fNecAr0QQSEIXHBXwagQ5rP/7KcrAZzqmfepSm3HKuZohVipoErej55SF
usuHdtmaJuLxpljNmICkQeDzoLuCfvSoGwsJgzq7nGLxMnq5E2CiSrq831DVChPcPoFghnojYZSb
OvnGeFM6fPndXkuvVDqR/+Y2UbFqWo6as2TVTbLoG0QRsp4YETY7sV/vOZ5dvdhaAwNYkjmJRF1X
7k7QzMVIjXRKiCzoX+iFfeF6vUHm+LHhSOnR1IXSC55FLZbri7AmHp7rprz9c1iYt75TP4+VleH5
Foa4/DQIHQ4FK2mqvYyRkUU7VTGj9xXikYNczvwMa80tEmFywmlrBZpwxqp1/bsfPvg/rdZYKFjA
L4vF+RxHycWd0f+FTt72poDZNi8thJ7gOqKt2yW4aP/LzTOJLmgrVI1Rm9dGnhoyySUOzAidDtjx
rw7zh53Hb6cqISE4U+oJNPIW3oWou4iKBfj5+jROHqiACySCsiY7P4cMwrOnrQ90NLmF5GnRgxC4
WBKo5cFD14kQj87268O+0F6RN62xAPaFPIodtMbGfWgHIE/vdlW8ZolIZI6kL+jY4bgl2pQTbDrJ
CBOhEAWiaa3Bsgvu5rn69EBzsevGydTS+dQ4ifz33yxcnv6dkHrhGnV6ukDhbBW38M/9v3/gdBo+
hQepQ60JxGfFlxDlknTqkBJl6XF3k9QD4OOM1w4xaBHnNgcVIBE6FL1wsGK80pwxZcWg7nHGSFxv
RRSRftVmTXuk2m2n7JZwqneYfUIH3ddcdq5iZFYhWFZxUWPiOxj9+27zdg1geKPWOiouTJqoWRtB
g0hMAscDGEjmJrTnnKTuADm7T7clt47RkJJFD9cuKx5CVKy4I3gBoZHkpufbByd4tFSUgErak+7q
Vje3Pc6G/P5GB48wDeuwZCFJ66wILYWO/dVPHjx0v6e+sBeJF1Mel5OUT9jZq1ufLg+8YyEOFSxA
HzadO290remVn/QL8O537LT1gHcf18jW5cr4goRiYhdCAj4WkuX5pl/o2gaeUFkUYX1iPNXvE9nY
0LyGJiE+6wclT7BPyrBq70uIs9pi9thlEKlIhgfMLuBO7eGr9SwBoWQegxW/t3uFIdErQrsOKjgp
63fX7gcn3wb94u13EH0pk9Db+3jWW+BBFRevyHaKw+DzFJVobpL20bsI3bt9tG09ozLBmfnwFfW3
+WRqnhgbCzE4HVcckJtElJTLsPNxbbz6V/KRkgR/Y6LvP+heF/KCYOKULYHLe9KzrvR4kelIJRHl
PB0xhSsZdbEwP53zjx6di9ivEbrn3pnxkxXSHdvRseMOuMS+Tk98w9zVAhMpsQHmLT4m5NM+5hS8
ZX25Oca9SFQMwIoKkLUgWbzOzs4BSOw6ilXSs7T6IGMF3XGHbwE8PFtdcd2PhWLY+SRbJCTNn0Ab
HDAENP6EmwUZBt/EPOnXt73wZ2O9jgfSuBDCnpczj+ISOXQcBsNR5nLd/4LfaVilQntSJ5jXRYen
2IA33MwxXTGVsVlYklOP562XZALQdqVMKBtu3zZyGdxxPooP6XrIYJ4HEMMZCxrmjBL3KpwK458V
Iwfp0LQ5qmawQXNn0I7cx2QyOO0oqQQQxWWerWoyMDHxBXOckP7jqNJDY0tAGrWqWaOhuHoh+5c4
OUw3uMMXl6JGMp7EZjMUyeMkCBxcYtayHtmcMMQXD9n1JCCVQ/pputfhfmlfGsE2pe19T4XvlXnh
bpVCaIlcG/esN5EBwgfaToJRcIpxIGXTXRVlWaXHNCwZzzftEu7gjrcfdXaGReNghDQcf4bppK4+
1c03Emzq7JCN21+2Si0lN1wKn4Xt+D1hwMg0aKcmzHYJ1JfyIATcYFA/vERUWcIFUIY2UaiO/E0b
yaJIm5ReLoqHHYDtd4bQy29A7VlK75wR/mnVQvQPSvPdYc7fG5+9HJ/MmPbEWrku9IXL95PgNRkl
iHkE5lq5+dqZTqglB512dPSm6agPqz7xPmsdtTR3Rpq6LbB7VRSjdcBMrAabUh3ojo61L702dUYW
T3S79MQPVo62bQdmPNvJst0cxzR/ENZLQhHsPQObgaoK4BiaEp8/SUDCXpXt8Ef/qCTnLS0b/fW8
wSVxA5qiRfa5v+K9pnF5A1pZ9vPBMJLV0Y2BEZg/9VoDS4L5XaPfeduz1VLpYitphUe3rE+CvoVt
FEfndLdhkTKgUx2vZXxaSRQXACT95ss14Ht9x9JsE9QmxtfjMAy0NBOoekrejHOgZ1ZsnkiGr92d
FOhGasO1ag9ci3calAiskpR/8zkpRIF9QDiPjVt9sa2MQsUKEqNm+rRixmx/jz/CEWv73tfi1OCC
ZLDmJRlbhk5vgWgRvXB9hiPNZs0Q4Bj2nB867mrys80G45FNXMg3jFWCnZM9Yt89cdb/9ot8yIYH
lCJ8oaBC0VjkMBNYQGZp9E7daCb1yDbF+u3DeyJr6woj9+6VAaTMUwb8ksLtGb4uyhIg8F7achRg
jvCTQUvT3eH7ny+jBo0SKl44SdrcrtIkpakYcVAediwqGHNt0loTKuuS19lvgVfzx60/nwRj04Ts
OJL7Kv9GyHn7aGmvwM3ilfD3x4yFOK66M1V7CNndfkCWCpe7gG+utlAEIzn+salB/tEijIiuynqy
QcX+JJBK7SQzYRekfhPhkHWgwgUZY+8/7rMdFJKFH3BLcvzc+lwWUrvUxnk0Dxac8ek+asoocGTa
5N0wtBR6q44migxh6vOi6GQF3bpnYa5NzcsfRAgl2wjg4FyBbPUCUcs7kHn0Tpy84EC/H5N2FLSx
XbRmTFBr1IKLJSBc3FPkJpQnd/HgH2zBZ8dPtjaZBwHW7SIzQl7YFd8PBvr4BK4MbgXF/B5zEH2C
NeUwVm6RKe4SUhMosq7uZVpmbjrKC8ZNlYR39sKD6htSMVqcDHlP1LFE8ZfTDI9oeNFEFcqjPMJg
Jcanip/TBxiBjoJ8AwYD6WYKapFwMubaDY+rI22BSv6MuJn6P9QOM2iocTQxGd8+TuDY7fi+gJt+
pGagDO6x/hqYqrahQ3WyspuI9POAh6XS2JCyOuhuvfu63DwpZEqQB5bF7XhHN2wdJbK1JxVrnpqd
lyFGhsA157rlGBmowuu7nGJGMQhAJ460HjO9FonVKmI2eWQ6qkgi6CjG7N3KljbDlrkwD4BkwJZJ
HI0u0Adz5ZwB7Zwve8HP2Bsx69ry4evxBDFuVBAAVQxqhQNijFDkCOhpUzYXnXrSp6iOCrwzh+T+
O/QvU0wyBsRvmGps0yhKEgXxst9KGUVO1hhbkEczS8+D2bwlzPxIV6K9S6GMNz1es3+PhgcknwQh
nw0Vb5bob5d+JpWKmLxIgx4xgj+wW2xfUJZmTqJUJrwGrSMYVYVhyy4iGWO0yC1f8v+WrbGrQLe/
xdfKoanJ9VLXUjGl4Ujpdi2cuZjdyQ0dM/xeBT3H1JqTuwURi8Nd/514IhCk6oF0LlOyFV1EsI2G
LJrgTcwFS5ZOMJGIZX8uiFmES6fLmZK2ckx4+5iKf4bvGUy3hG4Pq+4usPSVoVgUE/o2xUerkF8K
ktGFyN3Mf1QigOke5KgEWmnP6pCDBsrNnvsbi2Z9iVOIZ5EGdxgNQ/LGI9x1WYLhGOeRAFPrK0WF
Du6WMQbxjTIzjhEFYyvnBFAREjJ0yv5mZVZVLSvWJ5U3izCb8Wvz7Y9DzSG9emp7ucqB4cQ2yTNy
jC/OAjL9K58h7wrWvaHQpPuXVPT//hWTC7ByZRQaD0T7zQ3EEodYTpvwCWEXDi8IDMinFBQPIpJk
zUUZJEd6TERXJevVdpcLDND/rzXf6E709gmXR5hHpPlSnRRAYJdHwYRxvW4pX4nX8hOREdz0zdZY
XFKO/yEVEqZhshF7Rdc/SiGuuiucgHgSoytimDe7iKvcyQyLOmhE6ewbc4/AbyhaeEF1K5TnYj/u
wrakc74odG2YYX+Zg3Q+8c+3HTjiHYdrli7n12bvMzIbBy4keTHq2y1W//dprufacshOZOtvc1uL
qOqfB1G1RDN42LF77F5ZS7L175rQmgNvgPmZlDRrO4ChyE8qU0eCXNECquAnnw4SjefAoiZujniX
RkYBb9uKX7zczYliryzoOtF3IWUZMSmfliPnW/2gGC6XNH692QdzydzJz1lc6hK6KSY1G9HyaifQ
5k5GgeNw6r6wE9VMcJ3KjEc3V35Nx1mdJTj3Cu27rE3w1MebN0+BHkBtnnhF+rG12cIgWqJmHDjv
K6w6kmr1OMf8cZSV3tvWAVxQv+7oDHtiStXXI+5W2Utj6BleeWny6x0nuj9hGQZcDP01ZD4ff5JT
Qe++eykCTWS45Sr5pP/I/YIH62lmV4WP16dx0je5KqURkez5aFWtCMBsEysvFktuFegK1U/9DNQv
8IoXL+PIpQ65E2EGbM8WLaNPWTOnS/6JuFif5a2uv3lNmnQyunvA3yOLNtZ7dbZFB4ww7RxgW7Pj
0L0m+fLpi9kZCkYr1rg/N4hFTYVJKpB6yTjVGPLaBFADAR7Ca+HH2X1MU3h1W3wEup4PRGKY+XIg
T0YTCf6Hajhbamka78BlfONag6glevKpC1QMMLK+rsWYeJmLYaXZxhsLsjXF8FLBVRdTCIts3Fen
72LZHx/SuPqijIi2wTXhu9F1y0KkpjqAPc0w+MDFaXsZOYcmGM/kWE1uhxEJk7NhEOjvHDOHN0Uj
Vn00SicVBB/fLvZkaFJ5x1uMOV16crDS1tmoeKuNetSgBtpLKY+RlHEocWty4kBlkmi/6w9oYaoz
mSl2GiTIRwZYejLkBS33ypkcqND7M77Kf85nK8ZdeVtLmWNI0C+bLTV1dupWGrVTA0w4qV2uXCis
/FS77+VyZyrEO8qTSrw+6AJrw3XXpXfsDSFb4Onl90SmBheqDQa1PcYmSmZ5+ShkEtdzn3+BRxPL
8lYAQjCFFM7k4w66EhY0JfUhDWmGfY8+Dy3IevSkPM06k2TQPE74EHVWDgHR5FxBG+ZrqPw968+k
Uksups2weYl+2yfQ2WaAYT/EUrO0Vf12FNxeu0svTwOZrNLv6L+Z7G2/jVjWn0Oi8FYmumf+UJa1
3dCBuZAxl8Fj922uTmFm/qv0dAE8DqPU3nuwjPzZQEO2/dOjFIDrnNvr9vpcNbvk4RKnhlulJYaJ
s4+gQ5D1Y543p9kCBjcsYPnsTY5oY9slb6Zg2lLY8cAQ2LgaCU99d6ALteqHIRwkD8YG4IJo77hl
cPKz4NzJbHqkWZRSmABuB/tqMLE93zRR6gCcUUUEgQQtxHkQxYc2KJxhuU172EQGalp+IDdSuFD9
+SXfkukACAtPmwE+m2Baje3F5heyD/5I/RXnJePxjDIkk74WUn4M5yAGLR0/X6YGDoOAeKAJwoke
30J0/nJu9r9/E2RwuLYW6/nZ0BwdUmbT5APvBOYvpFFJ2g5m4GP8Qq7en4cLCUs7c7EqjRmtQVts
wXscvpL0tJAQmm2d5nfo2kH4GT7rqNelU1QTYIm181IgT6PEzmVX9DRLKKmFyVu43QDKd+WUJpuc
7Z9YoAyveGhP/jk9OYHKOLE65IuT3W4BYbNhL9NDs9eIzk5LEsljWYGSqbh694tLICTTyxS5UGnj
w8K1q+2APTN9CQ3d6WJe2hPQ9d3v8eWu8MzudgfYmdHj0LXPbhuIDBNXamTFM4gRiXpbcarFSxva
DJG8QG9TpYha9OBEvtsApFFFFEDe+/VM0YiuLdUy0GUwjDOuaitoqb9z2Y7il598n12qnp33CVZi
zxspaZLLtfmtxiTsrymhkr8nluiqPMNb5LW0SCY6m/R3764IyY/9OKalCAXze/kRi/ZRWWU1JIhG
0x2E/bRkrUEQCXx3VY3GxRZ54w33p7FP8eOqX12dDW24e9JbqKSjCUwcTCTo2vPGq37ncd1Bt/R+
Bea6UoOpCjsQqLWhAI1YcBeHmMb6PSLMUGj2uN/u49PQxYM9ql6Ol4vBueafbCIrBhaSDUz/tA4v
NQy752z23emN8QXfgQ81i9GBSi3WBqcy2wQDsEHHuxV0PowVtp3A2AHplVNSMvh212NqPWs2s7wn
nHJljpKXdP/TRK6AFQwTbsUY6ELvqUxv/XwSFagXCUSV5xD7gZSK7ksf8PJL30yBNgqWKutoxla3
PWS0ZgAM3ZrlXLZ3HYRY7L1HpclvGvRIbbxpWK422fTw90YZgwkz9gPxeL0CIMLSvlInSHr4sQXX
oGd5aF8kyKDiNT4TAuj2vjgkhq2UpKcWPjUNJwqMCpYWZmUiC38n7gjST8nlKRRYTxdeaz3r/HjP
vDXhLoh5owbarp2ppwwnYvOlDOZ38yg7LJc3op52t1Elel6EkLx5v26zmF4wJmYGszs4jbG2l/Bp
HkZGLkOmkSLdTM5NxQi/x3ZoO/8lEoOB2ORTiyaML2nwS13mhslOZeYjXhvmn87JYKKmE2rC+kMX
/I2IgBEVNUKFgJqDXQvBRuh3x4WzvdVKAzzwiDKQDdQ89kRzXhO5BK2LJNamOW67w8wdUVq3dHF0
0CsSN7oQg4aFs15q32qQd38BB/peHwlD/nkkPrQf0xDMvEUbWRfpzqxtfLXgHyeutpjSYFStH0hb
qmg70TohOn1gTcrn9teI7hFVDuu4Ymm4XCPNO5yXcfhrDMk6sbloBohFlWFwGvkJttgS+sghzb4H
KSPZ6blz3Jlka1KWQxbhfE58vBq1Tkxi6qS9Z3FSuSu4TnSIjpBEKRNWTvPTi8FugWOR6K/0Zuar
LOrBywvOVnTGdtL1rhPUYAfLWdUtGQtVW8wo1L45OVXBakWLEZug1s4u/6ZRQYkibOPS+8Xx0ynD
/KhMM6z5vlsmeEN4cWTLkiC//HvKrdbrHL5UEAuhxZG6hCAZLY9a5sxzkwRTUGkj1YbBgnTKsTV7
bePUlCaEhSyw9FmvhCVx2DGz3h1O5jgQEcNTFyLkuWLvCMFQR7G0W/vDwup7TDIjH5rqXqiLjjOM
MaeO7LjLjwmUNZ4PSHy1Fmi3xLIqLFnE++5m5zTjn6luuu5dJmsjb3tNB7pIFUINu+6v5uPcvtg5
Ti8YInuo8F0ZIDaS3686Gvq//HXhgCp7icTg+VqFROATmHe+AfDp9sPgpeWwLyZb+ruXvPm+np8R
Bj7EZjJpfvCS/ZUsIPLHeQIKcqN4WWnc42oufaGDWqtXBiofkdLW2LrKPay9wiTjtRbdMZFMbKvU
jcq/UhtgZupyzgcoHYgne88KPKfwJegXk4MZQZ3ug0ePjEvWMMn8mdaTKTb2w0KN/IlxCn9f+SQ9
NlAwSwi/GWqDRKOjkSMUvoGMDbdXiU6+TirOJCwsaiLpOKxwRU8lDnfZVGEL8kYqEYaAFeVUWnqq
2hsFy/tSQs5BkHBlrkNojmtOmkU+qStL/65oaK05jQQFbm+PcV0tZS+dH3vRb6Nru3L/5hfF1Mve
OOpNJ46CS+P5BpIMO1xB9yIahn6wa4eST8XdEw7XXh+XwxNSnOSidO6JCL2QXFP3oua4+QCn0b/Q
LH/6HGpAgqAPx2eaPsIxYYOfvR7cj04YIP+nAzN3A0ww73qr6+XhqluRCuwwKDiqrmfQE56+pF+X
jUDV9ZmLNfrgFmhWkYZ04dh4e0kI3ANGvVI7bpf1KnS1s0scAE112mmJ6Zhrh2Kk5S2NYWVsCf9J
QDnpASklE+RRDSIv5ebYhtD5Zv6LZLiVsiQrsQjTAsUcz7UHIaAwbQOpR42AeQZbQwcsI2xD5eDx
9vrWtQdbzafGZ4biLSFQmLjYVtHg3LM1bSefFIBLKk87K5vdUsWHivs/9+ZZjNR+TF638D87zWxG
tGNECfc8C9T6BpXqnPwCuhhFptFtTbN9XqYW4MzpHCWMI6TMETeZZ9dTeNi3E+RtKNdRfTkon3F5
IHsvsAUGgtjzk/dUCSWQUCTk1R2ah1ytoSDFMFPcr8mBY0Imx1s/Kgt+KMhw39H70r/M/g9dL02F
OSvHHAPlEUEpo/MT7a3i7bdD58HLkt0i1BtnRwcp7KbWWhHv1wphsMOIhdRXv1MNSiJbiQZ36nH+
bBTrCLmCtX2JGIsCg4NIQaFIq2YHb9T7aO2xKGdL9e2T6vLXHkvt2Xu9PMEMELDCk0raQa8NhKHF
xhL34mC5yVmLl9lu01nJZQnE+PHLW5XhuyVzPgA4QBzkqJ84+jixz7ViBGEyVsbZ8BuHooeUELBg
Gjpm6llngRlFGnWnmcDWJgC+fBjfp8EJ+3MkrnGrYXtzrkI26Vyzrrb4bnNawgOTWUK9biqwythp
lZW9+IfKPjAqBIFINQXM5bfPRauiCDma5wtltWBpA8JTtfnqF+N35jjH+JFv6/2Ha8OZFQEDe9A5
0EN/Q2CeePSV6wdoGxPb2wlgvjVIAy7MXJBEq4oeGFXZeAsGuIJXQ7ZsWnWM9NSfn9y/bDEsZ5U4
+G0UQvxEoyQLbxiP3tD1G7CH26lvkviENk7POR7u7AeBmyhao3ffZW/oVdy66aaeKK/RwwZolWj8
OHK5bzK+TB5VRc45h9dbX9GM9Hp4L4wADeVSWm+8dpfiM49Mk+c8pHdD8wguR4I9il8ssHwfniA4
C4PAujT7spTXR/u6E+tnwAfaJ/hA4iHupHgE9CPT3YV9f/oT3NV0lYUrvBNXEMyvBvGBeaPNPMv2
5JHlqgD7SruEJdh2V/IbyYXQbfG2e5Zh8g+XoRHJfh6ORWu++Zexnv57T0B9IQtfQeMlK5w8oces
bWztMeNg2zFR173EZMwaMy5tzBUtU+ndMlqu9YlT11BfVow++503kJJbw0Ad0dQF3T0BuyyUaXkF
Tkv7ZlYNnLDXLxrDydfINENAYXLvRqD9ONVD9sa75Mu8Qlk04RaFGhmR6ZvGsSG46nxTthJ3NSm2
DbcS3bSe11kXiN2MtVblYJtUlYm5qXYF8IZNOZ2PG+qHC1DAUZH8pbidEptlvO2eKN6NeHzGg3DQ
kSObOMOveG1bRibg+0JBgvNBdI9FbfuWxq2QxZC8L82sd6f6gKUmzXeDwPWaqI0SMOxxb67nxI87
g2T+9TPy148TT44kTXVs/txh4eCSrUo60475yicK/9d1ilbODupH4kyZu17zbfnJJOwRtrDFmDT8
7dZXwVi4qxCx6/HqpJ3bEyvtclVKZIt1MjavouVtEaR5eaKL3w7s11a6eUwod3dSM0dwpuGo9UKo
09o601C4jD21VM+fVC0zBfoK32j6vIRVRTtrd2PGGMhpWBlHvz8l9k+ACsXSfP9Nwf3WuGNXqxL/
Lkl5QgjOQ9vgwW6ukmoEcBIiEGlU8upXHajkuiYOPzpbKq3K7IOWrVBJKRwz+KMVg2hcmPVbNhP4
vzqRzrEKe4KS76oiYiY2gVmGdfyYnqXk+1oe8P2+3W5yJNOLAkwPud66n+knQRz0Qkz7s3t4vAdD
v/+iKGLgnrBlC8ef4K3C5jiSZoFBNq6Yc/BtNWJzleRFAB+bH7yxRryUqyvyDTVHaDjsbjd+55Im
N/O42VoMoss6lHrLnVqUXM7+/TFBKL/qTPgH2/7bLZ1e9vY2NP+9903MnWwEW3M8rTZQXQbi3q7m
FiBwB8BOTbKJgAUk21c93Wv77yHxon6VV2Nj9FlnmmOmbgROLXRcQVr2rqdOhxy0GDWMdcZE7V6U
W+6vzcpgdqopcwQiCSY5UcpkxfwKFIQMuqWwLIc7fDkLgjGbs1xwg5t5HhElkfD7U2us+aqAjuv2
SnyOZbueE4wodZfgriWSbuyNPf/AW1kTpJ5h01IK1TA55aF7iihtNYd04XzG1LIAGIyu6JdRBpZZ
iCi1esbijiSUXqihTpiiwViS+LVxJoGPSs55XPUsWbrr8fHWcUvczMaEXJHtNux8B8A7KBGbapuk
iW5LqfyketR+R8UOMWXwPD/myZnNq+cSa8yRRcVXS1kBugA8FMyAU30bM4YSgChOw9+6hBdAkves
BdHX3wdYN+jW2i9ZUsVq9ql8/utEAP/RfcxABL2w9gJA+XB3BMHLW9eltt5AyeERpNzZ0vrw6Ksn
wCRJJ4BZ7tsB1YsnQRCm7KLAAxDlA3LJg7dd23d22LTtEihVwRX1AMHmWG78H1o9fUkKdiAkNZlf
CdX7sdjGbXlBYv8PZ7hLOpFhK4vhgEfpOmk3rA4SK6vJtb8KLG3uqBEtkCxfhXFTXBq2sIG/vBvR
QPNBcp7njVVyXZJTo8h+lzt334kkKWKI5DQQDCJVlg27S5gU1y+5LXmTbW0024HcGcPPVOkYtdGh
ckENmJW+oGvaCzfq485xoixF7S+ml7s/9MJwARIbUx7CsFOERGMhyyK3JQRRoSGED30uTbA+JfKa
EhoZtm+0XHtTRNNzkoH2y94MVKw+57+zzh4MIxqKJWcSjyHjav6vaS5lR0zpg1Xa/84EWjHJCSfZ
SDboae4RdUQP0mk7gaxlS1GbLRvLdPhpXYga4HIPadnowo/ZkafIkKIj0qka/jETDzyvGNrhbONG
G7LK9deZXhDHs5yg8CaRrg33YzJqMihgNExN/hdEZRlfyHCpgbS5nK+BtmxMd3Q+qjhubdKAvCJf
EJc99QeQeLzetAKk7KtnqcqkUF7bMFYlFdJNH5Yz8dthZ2pSXSGQDXmLAMhRvLcRmVGpb050lnP8
rUEYOsaw9BynlJQY9MYsmTYJTFXiLoqYR3jDaJ09Ze4yHr3RUnoxHbA0povpxrG84mvthhKdifjk
auOdX+Yr3fQQfUkUd1zCUn4y1pBz+HP8jmJ2oQtxQvNXH3hXZFcdJxp198y53jE40VaG65Ux/7/e
ae6tvNJ+SNjQyV/PxNXBO9yaktLbHjLkgFpMUrVeOZGJ9YNCjGR9BZQ7NH/uksuwhyF4yhvLxqEt
LThAlBkOciWQS2wHxPNE/dNQ55nW1QBt6BtefWerbLbXj4ccn3WB7puJEjGrThePI85gY7Lm4IAF
5lGsuo4gj2UYYe3mks2vrT8KOfzPFOyJkU2ScetwS4WRvzm0FzgkN0Bw8yKCwBHsZI51NhcOu23d
QY50tu0MG4kbXAa/WfdF1/gedsstiPi8b0vTKbsv3dcazdTtASp7pppeaF5H6shmd92On/rr7Cwo
Ig13PbyVT7tmQxbkCbKs4Wet9w6RwKbQcQCjM6KqmbCR/ehjtY9kCIzdmKWbq3gRFxAmHGtwuB7j
lrMto6lKUSjL+WVo49FyU+N/G4w/gWlfsJHMJqJk7z+NENeu62GogvwCti8zQ/8F4DGLPbBWh5p9
pZgs19rpbV43XeZd9yXrzh0SxFWibZ0REtvS+3po/rsazIWwxqAnCXWvacKbLN8HWXS/OkwVh+OS
k23oqtlNujha4DtC4Y3ad3nn1sV2gVwTN9Ya3ZS/DcyZDWwTCMUiLEESCvp252cSkIS7PpByK103
vdvFcB6z7wNyqKLa83A7C2+q7lo/vbp/y53YKrWOhmV8Cyo4sIITimMgxXk27xKfotjRZaxne1PX
Fjw2BUz8EAKMI/E57Y7otgI0MOKoTlogfntpq9ZJskOXD9eW/xSzWbg8QGTBwJUfA8z7Fe//UIMz
xJqOenebZVPpYAKCkLrl079IIf/bAjDckAvNhw+aaysIhz0TALHaNOTnM8m4SbZQyZLIadTih7Ni
0mcDB3SvbsU/cZfTI84yqehbQd72SQz6vONT98k6Kr0V2nAVhZM8Nj5isOs/DV+GJyfLmSUr6BUC
X4W7FyOqQnhkUKUWksPPU5ZQe6oeA9jZrQowfPtLj00nG6/1aLnUtcX6lp18rUU/qAN8M1krPArK
dRlmst2aPix+aoPu92Lin0uyGqweufsbalVNp1p3amusQ1IzF9kggKyCnyuurV+HkClelCz2LPd0
S7ByXq3uYI+3gZkUkxKD2e6kyxHznkDKMJ864XSgD3FwbxTB9VPJQSIvGc333OBSuKs7q+Grf424
nfk6u7CHED7RmI/2L08pILtCS8AyrHljolVf0GYEQKyn+1x8Tz1iBUvr4eSLWcchMuDzT+HpQ1x8
IuWJCAJ0VChV231XYq7seoF/GrNvnTyp7RDdwhcZ7oDtFl7B0KxbmFzwHLCqDuW6Dku9aiE01Zvc
8cswvfDSOWCFwu+USiIS8NKDaVC0jxGHDK0A/ba4IcOghxQvTy58fWkSrzrjdn4v1L4kg0wuvJ+t
5NZUJT8jzZAcmv6YJbEgzZeLDJjUfWKPEZFIDh/0Yf1YhDA3R90v+wmVlGZwalcn7xAL7iqbLHRK
lpgmdH9Rf+Nxh9ye1E2NQvt+ylwZkb8t1y0FNwD++r/dXf+LnXXVlr8bLFQwY1aoU+fLxbBp5Nzc
pMlsIMFQgQGdWUNoggZklbOi2g9Sr/Yz6XIcL1JdwMVB15emz4lA2ZuW7MzQFwZ+f9nSfa9tJazM
yuh3Yzn6WUvdpaIQ8rv11xlWegLpRzfhAJ62rCJXLMX2Oe6H7mj3u+N05wxhl21MvCmDc1X2ylX2
Bu530rDnoPyyyiuIDrfZ2Mwj1vy3BY1LB4djo3GZ2UsA7nlGz/Z/HpJpIwZh2YCg6EOow3Z71Cax
4SiGZ2cbvUhJXVJmU33XvX1xk/a741DE4Jp3An+gRCO+4nHd4w8uJUmtAMlSDHDLuwgP4Y/c4IMw
XHV4DFgF3ey+3X8hEOxV2eIBrEPjEeALLs2UV1zRevYAWi8OIrwKgYqfwlwSvLOPufURRtmmF+0F
A9tfsxBzDCZOOngUnCMShh7W54/qOQDYWjeF0+q6Tbow9V86DqdELgqy6rUyGvxxD9PykjDHnQxe
mJi/zxgwKI4q+yWWZKk7bVUzyEzVuP/URdjVx1aOmm18I7ohAsRXLj82XN1t0fPJnll+F18i8cll
coxjjjyr+BrbZw6W1K3TCJk3KK2Frs+fJUCLtP2XnUiy+FmjxeqnVZPf8i12NbWtxelO/Gz2okkN
3FSnqx1rNVkvxLmlmYb7UUKr34veag7XjVfXJCBTln5lyG/o/M+6SW90HFZ/r6j0TxOa9slptAnU
BwR/LWrEhTzztbCu96BuczixcUvNIUH2TWEpx2aFsThbPMaPUGFShkkAH8eQ4ZNMRW39Fl7BTGiT
vCswSyWCedBi5VUgCgMwlovNRrI6AjXa3vDFwifXycbqBjfzXXJrkPc0+ZUpPXd/zv15suwbQnyy
mMD4TNASpHClsakZB52d7MvNzYfijBPXQZwRPuXMhbgwpr+dwbWKt+OoCXBV0iqDKG7dGbIV6nlI
Zc3J50PFwvwM0ToMMI8JX4uePM9eBnzOydFWQbEi4GxTF70F0gyG7yyQSI9YvJfFTfH9hMaCB/qZ
Z0FtZ+A5MSGm4SRRBqgpelE9SmvRy+vs7KS6ApbczOnbxtDUNMPdFyPKHrycMrugOct2mAyj560w
Rwm+MhpWQitSSJ0iQD1Hmkv+ZWqeUzQHEACb5sThEr+IsxojMFCKXiTQIkwFdqUG2tTvvIjlriQa
ZldbKHbKD6JNF6PmTmtKIvooEYQqL1unxpYT0lfUf89hjprQmgzjX9RaSA1P8fUqmdR+VRNx4uFH
r9Pn/5bsaH4PmjNiUwOKC+wcl8BNLxAV2LaByHwRFW2XIBE7M2SGQoxwEc0cKDozdNG+HZJzq+fp
wcrLWc1r1AkuLgWFebHKKur3do4W9JnJoND41Fd2UtKh/bzoqJDfF/g7mAbSvbv5a4+GnTZXX2i+
3njbYE9CImOHDzVEE0AEgT7GhJUERIEojjwSwcF8taYbx8O/zKc96xjOGi+2bW/tx1DYAIFYdjjG
AHurtMESyjIKdFFoU4lh0GVHC5FAmXyAcB7tQgzAdbNpnLXepiobLMrBNVtFyv2QAlSOwsBvajUj
i3qcfKpSmFr0F+1VwpvlNNOHTfbiR7pLXHyAlXpsbFmVuAkr8rOrR//BaGkDg4vOF1SNxy9VeqzS
O00KolQvFePUqqxeD0wOJXr0OCyHPc/xvtXx322qFwIbyVF3+FgGpnzvv2RqilS3l6j0jz1bHjDb
ltks6VwdLeCuI5HfQEmJKGrePmtcWfUjgF51mW3SrEc8pD/W6FmH1y9nL3n5zorurOC/7U3OYaVq
YLWPIXiDvwU9iUXQeKzsLMIcPmnv0VlFVg1ndswrmqisYpWWHU9fMrWpQRX8Nf1m8D3tpyyBlxJ/
N7lQ6fHZu5K+v1llLFqIp41L1UBQDt8IJRlODNzHKFLfA6T8QLlg0ws+AEn7A9LrjlQKo1tjvDyp
+3B5jl3zHDilkakuozytNXptN/630XthhHruEiVBi3cWCLkO85V8ifBRx/AM+Ato5DP0+TeD8XTw
UVfm65XLbME+QzUkhvUubXhzCDx07yAG62SwcqcanwS7em2LV9Y2BFNUqQZyOjc2O+iuXvBrG8vT
SUTUIaWgMUiS86sFwtdCAfNSBw6PlPI4bq07RWF/D53+SUR2cAduxgy1uUxje61L35TAO8Kojssf
UWgTIOe26SxQwur6Ebu5mXVHsShmiqdweNvk2M2iixZP97SElXHHF28fFahrlQHLd51QDpMFIdPL
oSxI96uvHdA9ofYKXZYyhN8vrTjpDoW1EiQcf3/VUrc1zmuEpP3NQxn7ID6Q0j+CgIODQgHYFzi2
WcCK93waOf+uN9H7jXxLovcg/79AWgGy2JigNDsIUMTsWAHj2Bz+UtTsuSA0WD3XCEXXMqQlHLXH
FPm+Qcq0+TOCl2vnRzkXvAZd0VN0D6E8MgTr7YVfMAAdE/03QKFKbVj8YF664cLp7ggMjk2ygzUh
rrPUQEhxDRyQWTkCXaySZHsFz59BP31MLzodoq6xV+2w0DmLTJlb3Zv4dKgHZVmyBhVMvc+J6SMC
Xx0diiW/H07l8PQRJidO5W4DXVAY4xowSHuxctXoA6pnvgUblmGWnnW7ZSPitYDphWDoipWFjODP
qR9rswkuM/I1154RmX1kN5oVKHaM+fMKJFjV+e/NHGQX16nRhU8CGFfT4QtZbPhFHFIeKbslh7jP
PEDqXOpRwTOTrByFPZZZ7pFRG36SXMUl4uqxNpH/gIAPKXBkCGggStapqHDO9dHfKIaKkyBAUdNR
LD3imMNMH8xjJwt51xXAg0owC+e9ctUReiVbhEgvjea95ELsH14kQgRNqF7v+nOqoRiO3h5HPa2/
ycUD0Vr734ZST2uVJtiFvrYJ5T05Nwevy08qT3OVcQVfwDGQCrTKV9yUvVL90jZtbdLguW2G2Al3
41Nzy/rmBMU/7PSSXY9PAKY3wMeKH2oenvDPHlFKL3ljKYlh9CYWXncL8ejFapCt+KN+VYacn+HQ
gvtRH6Lf9Ft9bYnrHCLpdmxN+DvgokM4E2nOqjwPXZaw6LrEwTIWVCD2j2TxdngNHoR4OmlwOyiL
QR0gyLWxjNn4Afq8JehNKJ8yJ1NVtQQ0rj1HZ5AN8yYim6UO35PGw5Sxn05WTxspOmMplCjziqE1
Lv0xWJfjZ1l7/Dl4bGdV+9+t6oOsRFT9OoRqQWFFT8p46SBjPeEBB87IKU5PQdAFeTX9h2z3C47B
vqXHZfhS0DoPGPsMsvKApNNjWZEyOMXrBpsUbueMn5qNaGQOcsk4qskhpBOGPrR//VmC2puQqSb8
dLz8qBbEzJL7ty+M4di58kaSUiqSpJwF+bseqmTMWEZCC4WBI9aB/RaXhvJzEEJYjBVoarRMfbfh
DgtE9lhuOi4119lraKjIUXvC1Dt2jSjxOhSFZizOiAGstpvZ/GH9+VGrWoOLzakn6ka7PS6yaVCR
TAm65KXYgy88f04LQTcaC7no3H1g3/0Hb5S0GojrniKarsLHaW5j5ZQDVHzNP6rkJYpNMoDy9kgY
ta/w0riWqbxhRbuiLIHeN/aCWO0BOUU57GyBQiBs3nrGQdyxVrKUPRuRjtAP+P2xRisMnQ23/zg2
q7nDeSgsIbfjDdo79Otxouzov224SMkwWyF+RawsMy+FaSQMAapPArZZRYC1Adcsy2LUpgt2jisb
tECV+tN79yc5ADMgY5yBbbAgChNuzJaZle6xhStbbglD3lW6jOdo+fKfSLpRDJeoL6kBGDDLRdWY
OWzMBtV2RRWqE7oUGxlHvYS5Jw8nYSAyfselW4MpI+YZhcubrFLO8R68pwctCj6RTX+FyOnluz2p
u9tKkcyZ1Hs8sgE/MZ6rmg+OeVniMoUNhUDrm0fF+2TUtFSwb8NLksixztbHIUyqlpnrNqEFBAlq
aGQ3sCmqPHuCZb4wCTu9kXxLE4LHzM16bbm0ioCF66/yfsSx6F62yQGZ9fZSu54FGjHP3FkIn4Ui
aXuUgK5XVaBxsVcgLH6Jubxyf/MIkW8CpOuMAyzr3Kge8v26RyrKV+MIuLt+Rc1MlCtlgprBOqZE
zs9JcpifabwXi4P2dZDJfa/7BDaq0TthP4rs3MB4ohdl26dB0w3lQLG6rNOsmABRPGhV4E+MHmsi
gqiAuBzDskezMzgtgIJ9qBi4iqbSSVRR6Fl81UdSLp+U5SpswhbXPDKn3JrKPsrTdcQce7kDxf0R
bxLRS/ga8KSRaHbHDWvhf5MPlypJRKTROzczu+DD/NwUIVm8GJXVuVBokZAd+EGUyR0Zw1qT7sZW
Th8NyPhjsY+t8asYdbZe4VYTf7BBkD5HmaurPJKx+5zPe6GbFnHFVisdxc+bGvFQYhDaoEuyCotG
RM3ANw8niP0xxFJqRdliF1oCJvvfVOTu9XBuOnUdXwdy488145TPw2w5wvCJfitzlvxqWrfrqsGT
dcW0RkniPMiIoHgreUswMewmyL46NO/AkJnYrb0AuugEZgyo7uJqTnA2WS4qblh1OEDJOlrr3/E9
WvIk0USp7i+bdqbgS5emN/OjaL4D9o5RqZGL9LNo6tvPLCqCqqsR4NplqhnpIHqQMH24Uv8fv3Pt
pfDIxrEKtGGUuRN7xYggv3eJSH94HcizYiW0xiGeYX3i3yOvq+kKDWZDcQ8drbMmQ7GFkHG3EsUi
7xxTWEMFQYM3O+CS4m0Rui/n5uW+VoZ9xZJq4SMCAyu2Rxo/COAM73hA5ZIZ/PCMopUidap9Y8YV
Ym6rz5uf1SMFZjBhn8mBVDNPsbGp38O2/110mAcFJ/Nl7AsXE3OgoNUuAFDdka6GJ9VYtQhKFdQD
O1loMOwIXlnDoXT8gA+MPeQW6/soncm5f4WxmcpRZj0BfphqFc4tsaGtQlgRBRam77MxUwQnooBm
laLp3gLT8SPKewpF6fdFLSNLhSFyjxedWVneshzojIMm560YyWTaVUx4zCIlFq2PR7icFZRYxrJL
D8oIZvGKmNWYyZ9REkFToffxyqDV0KE/ZjKiC/AEf2oSUH+EX0tSwMgog8Muu4YLi51E0gt/Jpp1
loV5G9ZdBemcFyRPWTbq23RprqPMgzecxcho8+zJujBfVOj8aht4G9xAbbsYPvaaAqid+sPpdtVL
KoppgFebaucAE5AHaEhYRfj03tlN/EJFl7EwrZobFZiXpLpO430UZDTq4PVY9hePhPNKV4cYXiZU
8hw9jqKU5kaKe2TQ3hVocZU5/+J2pv3oge1aPMwl+vIDiPb05GT5ZB7qLYW0UP+Aq4xYTz34RNgG
m3swfAW49diFPrfCbR/xgt423PNFSTIX68NtBFnGYfAwoow8bNVppBJgzFw0V5daI0Zriadf5sHX
S9Ky3FP6jxTdAP+IWOZEF2C/NkUXpqtPGMEqjAHGpIA2F3IevXb5UxI+tRp++ij3NGMrIU1KFQ+G
q+IPHBokWlfskGqFsLg2OBdxqanZ6Yp+SQEKXGj5ux9YVvrRWdApVt3HqnTCOsftRYi1BoDRiGAJ
2QloDkGlfuK+AXQFV9YnRkCLzsrchbP4I3jkegT0OPA9CC88Yq6rGN2EAydFhxDWHSj2fzGQOOwB
C0eJqgaOhrSYWVGM9WswJinLTLkseKztbPe0mWleDxwjuZUSNVLldVVJPB9CRXmRJk3JXeSFq+YM
nSSxx6eysMofH6Ml7/r7wPWsPBw1Upreu2y8N75QdgIi83D8nxyJIxOTprlHdS0PbDlV+OelU/Sg
BmhVr+W6jisMM/9g2K0rRf3Sf6IGNX5UXTaq4uWS7aUdLfIegfjyOKA/2MjYW5iiEfj5+9mNIM9C
nGd0cl226Cx9pxwDMkhyIlslt2N8JyLA3mstmVqda0QWkH+/xjHGjI5MeIzKyIUedlGyKXSPP9lG
zlOSvH/nLH1Sy1cEdXpBo8JzWVWtGA5WeEiDPR30+n6wtmJkqQ3y/TbspWy5oHKjXREVkXs7UYni
y3XS/vvqGR8GCXYwX9ydsf9wFBzSLx1MG5Nm/oEqbD0lQt8LF+xkH0nwV8I/8ypo/j/jP0XYTqrL
BRvy7IR8Xu+jjoMVPNncgqyQg6uEFTlhRZV4Ml86FGY8bbzMRbikKlJv44jafXzugBsQ0a/fdeo3
DLAiw9Abz7XQTY4VTd4mnGRrKUhk+9cz4kk9Pp/J9z9ee5+GZ0Vfog0EL09kcNNQrGvzOgwlSVHd
hWWjep2ETHL7/9JxN3fiNcUgmN/YXiN43jcR7UO8yZxklTl8yeRzBBHwGSwOu8nlKjJytRUoNPsU
amPlT2k+mxzI+SwlX9esS4qCMoTi89j5q/COVioGx3WRFgDo+NtfpZbYPoWslzfq7BTs3E0B+rdl
3+c5pIvWxcKC6zZcJ6iDMOidaRwe500b7znlPNSb+pHlhQis2kCioiEiNZ6Ll6ly/g7LfCOe0XvK
QQC1zkAXfU8z2nj5493zRqmSrmXmCJ3p6GgpB5clN4j14jqglszYW8FqvDT5zdlUjvryQ0D49QkJ
OJAWnTVzpMEQGHzrmbTv2N5d+BkDvi0VFSJ2WMNyduNIimTkI+Cpid4USE85JHU43FL+tJZ9w6Sg
I49pkOH9kwM3pZOL2/+aOw5mmE6+6Io2d9PE3KokkusL0eW27Vca5xvBpaEmixx2kciC2qTjWgzz
GMjxP3jYiOQvEyGf/kqyCMpwUc9nNCSz6Jdxb+9KWSO2EqWM6aaO6w3PryGBvnPBBAFfdiMWhHX5
7moonTxRePiIkYY4gG0e3UJqd957dyXdPoknJresLOV1rpFH60xIylG0aNdb536gg2mLq1huyVY9
EV8b2kkj53nBHno3mUqLvbb90Hw8N6GUM9/nxtGxkS9Eex06vhxePOL9JszbFFZVH21oTP3hJdyJ
/TMFPyhMteueig0ksnzcoVUZIitEAXHlTo5L5/OWtdb8us8/NJSjYObZ79A3MmefsTuwttcakpFl
R4I3YU2aeSp7iaKDQqQKApkyAsxOLeulwl3BCALdaZtdNP8n3+czjtIVyUk8MEHu+ERck2JTD4if
91MBN8NJXVvQFb4vbwUJft6df6HKQw+wyVVk+KyYcbtHfz+hkDDslYosdkDodEH730lt4gZi/xZN
oI/qqNGC/0uONNC8Twgd+qKR7O163DY9GCLnBGC8A27YPoRVgjJtazrEgqIaO12ylvYJFkbw3tcT
OVOz8GNrRYTA+5O/jmbERrV98i6SGWOIt3BcUevmn0xUCQ9WwxCfOXAwGoy1e+8CBRupmIlKdRwL
dd+9yXJAutJ6gwdIHBl90OgP6IlSWzV5qQAzMNZC0e1mEF0ek97yguwvKyGLqrtHyeEJeRteEhbL
phxTUYIorSZeXE7rcCr4NiHV2Xm8B2tf+IK3jYbcBmUmpuZCshXxBUXF7YkdWu/IFScmfPxPbRxP
BUrYjLFNFkU1fypLTRSqovZvZ84sRn2ifgjUB6jFw/6wuLWhwuFig444nSeMi2lkN1dvplV1CgrZ
6N+wMhkVg4Ce93BPZuNmHBWc+4mSt+gY/kJJYw/yEFnIMyvYm4wH/6Isk64Dhh+iJz3D2sRTUruu
IdZKV6beE+zg4Bqq35h3VFB0VOufX27ytfXM9pxo734w6B8dCT1w3W2fABDdfZWHsPoDP4ymU6te
PrwlzhD7WEvmuodinTSGRoXNOU2ziiWqLqr0AkmqXNPUepLhg8C1yPJE1CEHu1t4lJCnyo1ahy1Z
251kd29FKQc89YGtMKHrYeLPlZH5GDWm0GgQSbNI4PaTLY8XoxvQztfnyANIk0fXE8rQ81yKQJFb
8QGxgcIcInCuvf2Eh+bgZI8LaqbjiT9NDsymaJ0ex/8OeosBk3VsnBby/IAVl0Hc8iCFq+6/wYtX
3vnvOfZ/XzEOZCGtsKDS8Fv6UTdENxN5arBiG7YktuNJqat7DKnLDSopxINuDoXwsuNzZkkvB6UD
RDadr6Cl/dZMaEevyKNP1zbZzAXf1AhzSUB3Fjdwybo7v+zGL5kmNz95kaPaHrIjDetAo+1khuHE
Tqn7Gi1yygS3wwj4NludehdL+8VM0ty8smyWXog2bro4LqiTzOJDMhdTayCT12DQTtMKJpxi9wM/
Zwc2Z7UlG477A9/NPk9Fqpz8F9P49CL+hkRSL865deyGyL4RjqMmGOvwi26Tz0cM9qScCxw/R94V
qNLmCtGx/UwKQRIErpxRCMaffonExYwXIDie7vDLKzfQkCxVFWWx8YoK91qITThY2Fa6RcHlwYgU
g+Rxrl3P0onwqvD5dNA1HAz9L32h5R951U20VKyupyHjFEYDJ4EaeUInLnw3/19T1MExmt58BZ78
PnqjVbbF0aNSlxpdUtbTwTI2fohXpAeEHr6eqrLapz3yTCh1XT2l2cuAZS0AR0gDBrU7kbm1+nDx
FCJG0flnd17zY0SAzTJral0Bisj4RW9Hkr0e4mb/Y6M7d9A1vZ6xZq2g2Lns50Gn3LViUrzikxeP
d/Dtu4iWmDzXe/5bPQXkZZM2mWEoalsAOpKx7Z5ny/zhvZ6NA+POEOSvDV6O1o9EP+LKWjQ4AikO
WOXbl1cr/+AsTr7nqHkpj8N7ECvVSOCrAYPIHbGD6HWEoTJbQQJPhtVSg/JlFcFH/+HLTLG1oGS5
LX8FOAPYwYJAyrXyiw+vwZFiyxdAL/gKI+9QtF+i+bMDsfWE3LGAbI2/r8gM5D7KTnGuK9MXRFt5
rvbNNAA7f8+/K9LHxmFHqxg/9Vw04+l1egxOJJ11O4/W9ahJuYHwPYyg2gsZg1uUKsy78JkQHncA
PcKSQYyyh4w5OqpxCZnLOKlDn+2pI4ZPvLUIsQ27dZUf6L7MZ2zZI30kTpVfu8MOMSIywRIVHDcz
yDGTLM/foonQ3jSzSi/CdsHyoctzApBAYAA3vrjWOUReMksd6wFNXWQDcLl4Rz6A/SNHsDV38WUX
qlGr/1Cicgio9y8A0XJOl0yjqjAujC/htAXvp85EgpQAQUiM4+2VmOowZVUXX2ukn6VEPoKd9wIG
XstZw7/JUfEtPEYu3xESV+OfwYdycy18Eo+5G3AqN5fR+6lVvbjrLF3ZbEw82Zjy1lwYavH0K+9d
ow/YHCoy+lq+aU/Z2K7YUqgMvekNor8R5PQAoR56Wk7DhIjevUiBqMGUjomP1jkNJOgTT4ju4coo
upJZvBPTN6bzU9wMv9IVj2SSajzdmOuqgeAwnayTmPAb+WRSkcuOWdPizF3Yvtd1nZ2i3D/FZBHP
Lz+lsXtz9sHVtgWhVsyDpf/wQXlT/jkxILZPQGSul9gkiiZBjba+8KeJuLXqDMyAXwdcbfs5K5AA
eIFwYYvet7cjhR4bsbwto6REK+nJmPT/r/CyFpNk1VLmjjyl/Wtd2HQpMFTAoq1mVVGN9vK0cGjG
r1JQcZGGbkVQXdmHQMuJviwtL6AmkesodN7O/puxyD6mH10rJMu7fNOoz2pobLjk1vUdq2g7/iUp
m4gJBHHc2MvlGgtw/aWGJmvlI4OKgIvf2M+mkBC75lE4aFrUMTJqZO0v7xCJhUhbNk9+VUXcPr4+
44c0cS+RB/cFegd8zuKWNkHZ6eqF7b8UIHCnId0RTdzJ4j7PxF0OJEo4Txz1cCc6Zjk+eV+8nFA4
Xkj/G0ALzO5othafHMIsVn774Uh+NLOaMAwWglOmKSZ2a+4mAdpQkR7ZLivwAc4i8uWNpMlJcOss
l0ryO34SHjd4rSaEXNpCaqdYgX3avrwhSZC4/vBHK6iBfRUxePL8qkZ1WRtyE+uFhHK1BbtDzBkS
ylWfGw9sQTyxdVwaLia61uWgvL6mBdEKkUGzEAuTJncr2lsJ+K8qdFOrlLvZmXKRRr7FXJgn2w58
MFaZzCaNY+tpJAwF4VwSsIRl4pkI3WCRjTJwwNudN/vxuYwnT/JYr8Q3j8xRX/FoR01nyqPk8XSx
N1yRqzAYfEPcI86UTlM9KrbgD+IzsyJL2ahEFcSLj6kCN9bncW6P8QVYDz60eUwtII5OZnlHLZO7
G8X+7C3dtatVk1pEb1DsBcI9gSzozF9aRpXTQn5E1YofekMh2L+ZyEAakqe98ihePu4JRf9AvunT
yKFxU2pmr+yOukZjhn+x2Fq50KCXjNPUN52Z1RHJ2rdLvFSEbc8IZMksVKnkFwfPg78EHVN+bHCc
GPMpQChfalCRVhwRO+NBWIs+oARLJIGrU3ilTni1pvexovXRfjcM5a1BDuI68ei7eUx0oQTvPwNc
lSGpjuvlgxBqzraJ3pYoH9A6cYUv/1QrhwO/7bZKngi1jSOsEGa6y02Wec+XGhKHYs2zljyYfd42
u+vAufw0fKPwI5ZCd8fLaXd2dpvV9jpD6FYae6SrELrDBURsvqUXRzr67mx4mnSV2ZFTLIiU6jpJ
lfB1OyLpuPKnMmQ/IRU/9rmVfkPQEMwTh93WCzZpj8H8lvN8EfoAeLXW3myiBpwNGRxM+wYmkSfU
sTeyBhzpuQpWNhPO77q44FNWobp5DhQU8N/0jhRkQOMFqPfag4zvBLCkvDIJCnSblp3kgRj5Bp5n
pBm4lNUiNRLh6uxkfh1QJ/y0muXiIbHoSQHcmR/TND0rwBwITMqoLpl/peY/w+uybayClW9GzbkQ
XUB+/yWdY/FMhOjoJAlSHxaBtW2eUCDPHjyzo/Jj2qKiu5brkdBexlMn03ttPhtIXxOP5vKYfOia
leuEI49SUNPy9OxnxIExP49y5Z8U+RYeMrs0xl3gJS1lfsKYSAvn8UntMNW4CRgEZJqPEJ1Z+TZR
am1fv5TmMgDwdR7sMta0eEfcb9FOSHtyYbIEf6D65RX8f0fPPcY55Ek4qpLNqCRX6EIsT5Kmk5qy
pIBU2AMX+LaDFcAmih8R4A40JOQl9avXPJ0CSoa9Kt9OZusOSIW6X22TgOdjX8/yzR7zjUrkARdE
g6EORgjXWhNSdPh3LyxxMVPniSHpUekjYkkKY+Kr7aB6kP7oKV+dnnOGJmK3iM8icgci/38XCmUt
O617gbcQGW077FYQjcaMphr43HbkGSdh3lvI1nsxAlAa2zbhPi07sUTwPI5uwKaZsjcjEpNc2STy
X+pIIBK+/Vjw18uwe5JJKEH1eUFWyoEUuKnCkmnejr4PeTkf8U+Zfb1GSwdxpeGbd5XUil99haNB
GQ5k3DbSqFxi6O1wkFubHYZPOBnVrzsJYML2YGP4QRhU7EbbGcbdBVwa6uz67NKSPwNJ5mXFw4wL
CthbmG1kPK6tgVJtqOEzVKKIRGK1fThCxNC7M2QHLK4CJIgIjzxwNxq1KQgbvkh/6hJBJ3R5f/jT
Urluj6FkrZGc5CoJuEoNKF7aVUphhaYtS6DRWq3ePFElCbXoVsxm0E4xP/MEeapLu8QmMucZle9W
FI7wp6UijdGMKsGTjtDxrtop4IOkWGyxiRw6QeNMtdjnqfaYmGr6RPe9jN7ljAQo3JpqWS2LwwhW
G1puCFk3BK8JId10EDiUnI0K6AX3MkK98/2Dr12qa24WVB1f2J72dGyISpVJ7f4H3TdiCbgVgDqf
ALUIV+3m1jcjtbDPEXpC6VWjTOXsg/fTqAH+rMI2lZCmzy2b8t0SWPNm3ptC7ZMAUyYkUwSIlAHT
APaqPbCZM88nA/ZmwiL6cKqsP9Y5t7DyyzWEks7Q3Ib04461KIwAFiySoOjR5tvdAzga7sts1gW1
xDlR3WkyAY4imz7l9z3LtDKNAukLaTc0/s0s2nAO5zWSUYurhvxzVRN6XNw2LbRK19X+rAm7g2Qg
GYukPB4AmHZkpnixRiwhYi+arkQxWxgnRTEEz+5cY4aFkc/6xXj0Js8FSigfLN3uMIPi3pjqrkiB
rye9vWSV4itIdKsz21gc5lVRx4+kpHV2yFBHMBLfXX81XQx/ORLPaEndZmlvn7SbbRwXJpUpsl1m
Zz/S6QSqQ5D7EqAijkmcCFtkm7MNhB+PMyindUXPXkk7VYHhICvRbnM8Bx6enaLkqly8/On4M5PE
AzfrZf+VB0JWhtI5LEzwdaKYvRmvhtYOKF4KU/fVuwRzfQ69hOjXcYCVtAoiySyfTcxwGMZwz5lz
eyyKP078bOxBSifvL62pIFbudnpj6VEgi1m7p/iDkSxzf8nJ9tGeBWyDzNIkfOHQqU7paHoVaejg
aM4HfXgryEMBeO0LZvpcvkCH4DjFDJpEbVAat4+4ChJ9uQkikWWkAKd0bvyOAKdQqA6JZkDbbxeR
iIAn5+nOc4B96tuvR3YqRqD3gOHoza2GXFfr8aixf1G75LCFZZk1XzYAvqDARVFaxvsa6aT+kTXW
IDki1TkMnSGXb8KeSQrBsBuWTWafRc9+0GuBSFpMZUlg3uw8heFje48kU+K3Rhr97vkMvPJdk6rH
2wdmXc+NtF3OIkwAaUAFdEyzReBKJhhk7URzxZtecuRTQlex0kgF3btYKM3DsCIr8l/Rvp5DeY4C
etwm/q1xUViN8dysB8n5aj20nlbRT2vgZ0js+7uYG76c68z42UaBjOyYoocRT7PYXPv5/pAQvwdL
VfVsl/nS/PIMyc7rubUT9FBsnc1kDQbNLHXBdQh+p4g5GAjOb33lG1ouzLR38ZSg+MsvDjpWxxXK
QNS88NLCuHuJ+MopJr8fD3yhKjNHPIIfAYvzEXoywRdIxQSYh15CHSSpFlfsZVWDVtZrkqST/CzU
XacGVtWRIiY3ECTRGWv24VIhZXAT2lNyoI8Uyuqtkar/IM2Y0iwncQsQmEd7uoi07gNgrV54sbqg
34BXibbsgP3FSGjHbgpfA6HVkZIgT55YvbRGXJq4niKoSouEx8WUnWGL+APDopUMQnf7guOrMtg8
uN5aLRZk19w3LWG6QTFWYnFAnyFsBTeIJDY6zZTto93wyXvnBqQbfvYKv3LIaafVfFK0obzuwcSB
XTz1xW0hxPiwt2l3/dK6vkA21LrB/h3g48oJxEg77DitXg7GsLEoVh+7Xl6Ve57/OePfMcW7GGMd
CIoxiX4ebccr7XAkhAOIbasosOFGXsFV8klgHvvl+qhUeFloGUEWcCSOPBXCsIq+EEciDpcxBvAC
Xvh7RvOg6dWO4utIJWjWI/B6BjXFyzIm6K3j6/fWYZ1c18F81tsruhPBRm9+SVg4ToQSOvwtBv6W
fxBpqhjE7ExsYlAkNXk8oo4SzJLzmirggv1kk8m4EtqLfjUYB15+Si5WWycRnfpgbm3QSOoOL90t
ISbEriDk/l0Pq2OdKgb5ckY6w8hyYTw6aFa2+mwsYuS+pEgtbecuqdBe7cM3KYdRh2FDaeqCVd5w
46CEsYLaoebHQPtICQCiJdJOfTKSeYinTY5V19hAo3QrvJviekrqgg98pCi3OH4TsXOwAy0vxJI5
XyGbqESUZ/kq/EAIVdpPcio0PjIOgxUKW2BlUiOoRsdLabiFi4uYr0/8m2P5n/QRWmz+aDuUdVzF
r14B0RWWZ6oVA+9p+wjG+Exm9w/ExVcv28QBV8wHam5ON9uAg5faAH+R7csA2E56ryjJfrkIFwxo
b5pfdysq4koG9XMaLiLJa0SApNeM9xEFQdyHFkzWGCOE7uYXMVL9VQ0Ebqc36xxS8SY+gKYqxyyl
fadhYX1llNahq5/AVel9lPqOdTOZkoPGt/qoD7xIV2SjUW4CshjICyXEytaWC5sP3HFqzenM5sHN
csPEWGkicFWbPdJtAnFzKY7Dx2RDnflcvrUzYkg0HIa4ln0qIcr+WkuojjtncDMfrjXbXCrPVOd3
4tW0V4vJCxI/mKM7QPDK6nvrH1jmHT4XVz1pQN9lahZxhyfU74TeXCZN+48eqjYL7CaqtEDwXfTg
0/sTX/Gk/b67UEB3XD6h28GCy0QpYXH82hpjBAilyqHS1zC6TDY1bvYVyiVDGtjNR9aXvHf6W5kY
1yJDh4UBouiCJ40T3ImdPwNJv4oc74PBBknDCnjRK0adUfNgwQw7gXQQ7WJzRto0aJMtC6nvL3hO
4jW2+B4SWfYxA4ykD0h0a6DChaf+7514xTRs48luEI23RCjIHluAz71hxFeLtkLROjv5cjgWYcJ3
d3XKsv2pYl8sgB7vrvjutEbc0zK+7sEntuFvYxN5n4z48e/Li99uTHu/vFd5sQcMwYDebhVXEY7j
ZOIE2oprRDVpANZdslumcM3oeB5B0KEjp3+9uSyrgXAC99CdnYxxGITGv9k+f1xotoUmGGVUddnm
oHllLM976fjwRCRAhTQid5d2Xdk7qw8YxQ5LIkSVLTZbJfoIYQr2zqbw6YsEfK1m/akB0NEZyjlY
Kr9+aJ0aQIi3T10/PSR47qyncHknTvJmKxoryALAKUET4HY7zo1sTWmB8HJz7A/B2cp4SMFlrX6K
82yvufFRpe60bhNJjTWtDjlPhVBiH3ypYYGZmUrGqKqaBeZwL3Tb3n0QTzzp5neqtKprL9g6vpD9
Frs5QteYhi+wpuYv0OY59F9wz1y6Qv5/M6mzZ+cLCbIuDXHAAOcOZWjXN03N75kyNOrf2PeOerKT
rPkZiLNNYbOHpcbn+XQylrGp4pCCHoEjeVfZev6LiYLDitTlBL1pmw6nZBHPFJ05z7HSg3UHKbid
v779VmG9HfhIUaQ+QiLPdVvvphSqXWik16hFpQX2KGeVTcrlxz5jcqinsSjJfoaNZ8bO8GnX8Mch
PpmeKiMQpHGlhq8IHJO/X0ZNhAVGZsPeS29DNFuKtg2/SH+6676EdGU+KIFwGOqpxGHPI8ex79tP
yi+HeTQIGhtJBZL7k6KLMZPc3BD6t/mL8QoeOfppKJTF/xNdM8DQAcPBFi1Sfwy/FHNIdXa+7+o1
xfzrwv4DzO/QKuA7N2xentXiZs8bjwo+VztedDbx8XtEIh+hpGWcFf6dpzJ/aPxu1It5+9QaV1HT
FVv6lFCw9Ez+2/7bKAbXFstJNVfimvBbf7Uo3pwZmzsLQXygDUtJ2DRisHucU8j9JfqMhtGFPpRF
ji0t1clz992o1bAfqeWqVwPpGSTuk2+KxkKQi3Y6mcjho1XnbfNxZ0rlz1r+Dl8743fX91TKr3kD
3+zBObOGTJh9whQIEksFAZM+blWUFDO9SCHJQpDUMWpU3eIm5P/f7qnx4cuAUXbb37PqKriIWJU9
4e93hO72ilH7xb9dN0V5spmFnKeBr0Wdn7EFHXnzrF+XDdz7wNjANZxrz9hrYW3wmEuadJ+fU1zX
L3s0cWIqOgHJ5CcnkKaqIqiWFFqUXABss/Sk7e8zWwfu/S20b7LvIpTexza30UpsxG6s5M1btsPk
LXqsaR4leTpB9njY1BfQ8pV2PBmGHjbovnrXHJeD1npZ/FCOFoPznnpF8zafpmMDdZUSeESGPowT
xEY0Q54ZfVvbW3yAB+NV9q39gt8KUKmDg/RKniSYKeyUt8yNdPN+zJQQhR6qLN76PjCqQIkNoL6x
RDCLAl5sB5xyTTxVOcQC/Mm5PIEoXbe2imbx99EG4ASEjC1yZDGpQia2jwexnltjLiRESPEHY9MY
d8ahucCjLN8b47mro7pG+7NNTw00kOQRhCyyE+lfHWQG1BLRMNcBi9xigCNu5kktA7lYq95HXIXe
JA8eYjuG4AD3P3IMxzIlfKTLWlBvAmSCnqpGwaAQe1b1PTuic+dSaiaRzAEdijdJRZQqHDG5F+Bk
G5FbEY04gHQ1+4K3JwXT0Khq+B5tmfB/tR5ud9tWPQNttzoIrHrMGgWQsIOLrH7NbYYDC/RPgRhO
pcuqVb/rqVKeIS/UCYPB4C4heUS2WHhBOpxBvXOHHSWyPgz8YYSj/OPKD6buPqMpifpXPzlkH5ZO
pfL6fqWWVbhrPTvGkfS8j2WEcf7UI/mZZtcCwJPxRzfZrao1Jw0Xv5RQX9b6mqBtfih4N6U2X9AP
wT+kXkjUoxXGv0Gqcx86puThpQOA3r93uyZ5aZwg87TD4o43P0FhBILvjUj4HEsLf38D5Tnm+7SM
+5KecpXRpuDwLN+1FuL7OZMEwYYaamVrRmP3w6ZJATFs9Gw7e25Nn0jKURxczvNpNl6epRy88BAI
L6UBYiM9Edf74JOlLvlWIeYdnnf+JsTmb3XqtlNId2zE3a5VmY+gkelGNQOYw8Q/Yi2OOw/nNY81
657iFmdAKuRWoQWtEkGmkxvJ9lVSNfQdHfUEtIwAvkXY/UnfBKHcLRchkF1DLVN03Eh8CmqABKWi
xK+6ULeb2YzwYPJWj04O20RmUl7Kxm9wq8HXtGBFe9GadLNdJeKGbGLaj5m6F5fl8Oq6AXJwiGpQ
qBZEhSvb2WAA2EubM7+9ZTFMELAU/VPoYazYMrmzYsq8H67vaZH8ZNdTGxmJBcEwHumkbMiPidOV
iilcHovZ9XxoM3PkOnyCUY2vax8LmF722TizSaMSzD7JZrFDtsKKEwbxnoYE1flrmsKOo5EDlSj/
CfbztpdD7X7DJ3leX15pLNclKDeZ8JbNE3sT+SlxehZMRdPKA2DMy+lg8dViAb3DKgBUimqjkUnk
hhAoXKh49PMFp2bxa1w+TH3ijDvIg3ViFdzcpKZZqmkfeLypjqg2z3kRYSz60C02NDaU873G184t
uMu7BIjdbgo+GOybu6v1XLySVSIUxPjpzqHASdp/YOvk2JVZMFfWgAtwa6LXCKXiVPc7i/L+6KNV
ws1t5XiBt9EsCVPcuzz4rmue/3aymLpLZVjCj0GZC8Ize9CDbkAnbKc3FHSyx4qHzL6vNw5I0ghE
MZsaqpTN+RLOeE0f5NRWTh5Y0EwpOVkM45pe10ot7GwbGyNmUXDr6yJAio3Eh3fTgUqd1v0EmSbU
kNy18bbdFqswCgVmwM7vuAt/AWSRZuvBb/aOOaXpxvw9/fftlFDFyDZyX266aCI9CtD7YXt1FJ9R
YLdGjVnsj9ZI7zvBY8Y1YM1hfETifOcLa8JLjJZ3hhsfcDSF5j5kmgt94rNWmQTK2pCoXt+JwoAb
Jwc+fCvHLjdYcUcgKysg8U7lp4Juu5O64NF4nQe6ccOSWI66rUMbd46vQwp0xH/+J6fm8zAI23gA
xRCyN68RIW0Vd18sckdLN3Y88yhn7YHEexfimoFr4VVC2HDTyCF+mGPNA3xAEemyO2FaLogs1xo+
XxeyKQnsK2FDdwBwnzhgs9JM3JDlEPmvklhDfET0199vILmC7HLrzvBMU4O0Gh8I1Ul2STmSqMaY
aVh5Ni9L7yqTog0NQex7mbncylu/XZitRx7loRnuC/1RrIJG6gGaSv/X/zEWOnb6lkOT3Fdv00We
PGmKCiUNPUXTvxkYHR4Gesva6Tn6Vxn3PRb7aBB20RfA7GvN7j+awwfIxupRhpDDSyIVXcF2+A7X
Bq1rjnmyrtCuIZlffq6ik6Sp98HDaTkKh8wQsOHDeeXhQW5jkziB0pVOo0AY1R5FX2kgQZ8EomEx
zP7tPeH8aVNfmGc/b44HBjrZPppMMa9i0AzaZ7AO/0dRfZY+tJ6Xd/AACML2EuB1HtVdczjIwiEf
B5Y7TJHLDQhR6gPSPkZR1wx56Vv1JD+7GrThN8y6IBwolyZsNDRjXJQ5OTwilt0gScHfcaeTjc2y
Fi7BLzI+Rv5VO/4EzKEQBwq3SLlrVGCMiqhs7xBCy4oIPCaVTfHy50GBR/gDlarE57Ri8dmR13sk
CGPjhFAAytG86cQNNfJ0gxiq1m5aNxz9YK2Hy5+vD4HuQOEr5r4YrNqQF3ZBoJMB6FA6szYsYNGH
EB/ciCBiHYTxFwz9WwTs2k+a+Uifxd0jK8IgECuyFMyEj+zmIAJAT0OdFzaHqATeFHDWJO1F5ICe
G75etdWq8fPUsQXnyigJsw5iOfYyHL0I1ljm6ReFvE/W98jQQBKKMYIJT/rJpDaZRNpnwFypW/AJ
ISLl6snmCOTOn1rtKsyj43mZuyJzUBQpLejbgQVHxn8tyiO/Nx4GBfoHtlFr1pcAHcoZKvfixrxf
eAlcNPx4wAPhOCUI3IsLOVWsXtkbjlneSw8aUgXVusZP/6Q+3Y0ZpPPu1uzwssPUrFh4rX6SKlO+
/HdcOSofeFyrutZz+phBAPrP01NzlooFaWoyEC65kMi9zOP5p5thPkHsNvVclGIDruuFMcy0kvR4
py0eSDX2ijHL+vqXrwGCi57UmpqTkfw7zoshr/1yj7uBM5a4t4cMJnCXX5P2JVrGmPQsjH62F3ps
R3Jp/toHyHIBUU1lmtwqZiEOfeqxmg6Cm9LCgXMFi2uc3F/VPcbG4LRz//Z2ZPtRZ2cJzEMb5BPf
nmfOoDbgEpEGHGiyCFEUwcWbnNXqpeCLtlsaa45vqbJqDOsOu0wivGEv9FHTVeSfNH2biE2NG/yl
acwfbeYEAgPuODQ79j9tbapFDTLpFR73lrcu29M1Xw8QYHsFFrAttUxKLpZpe6pt7pgdhXhIxDaD
igkB+SDL7KAraM2gkt7uJ/fWjzy11RhPoK4djo0CrnYteBAQdDUBEVENvqeFaINxf5zarQ9Jq7ra
RTw5XT83gQZHA8PxCrAsMSSriQ2qe942rpOtMVIjbbdEbe2gZWKWroTdTs2C0yPMtrGIwmeIa1Oh
h+j3X87Cij/pdKyL2O5SBEchmb5ijSOfdOydi//LI3BjGcTyYvExrFHICN0mzV9wDHywsed0K67o
31+bUd54czbZ4Ub2DghjklKwZissT3ZhjRDm9Fa279NizKn5AmCVXYdhf4CDR4V86FNGwrkTrVvC
cDlA4rIOr9NFGIzw98XOTjMjBvvdny59XCyTkNpf9gVj8NQ4swhFUUwvNWUpUfDiWjzZGBt6YpWr
BP5KFCH0KxIINMqEj5pFIJnGcFxLWqDun+70AGjrxSKX9v4tlbWLg79AaGdDOAn9KqKoUMq9HSHd
un3Uo6aUNH6IMac79FunVFklFocopTY3aTSnXiqFlVTyvmZE6Cil95eAhTYemwDJvyzcm3a0Yufp
fb8YP0dBTp/0KfGAmsVKT7fA+F1PqJ3ZDIOkxykN4+gSFzXBQ3VkItKcnIHD8naC9v70s0M6BQJN
L/sALhwm/Gez+ZZdzJMGG7t/7HJ6YNfcLqnoXKwAK9utJ8G3H2cs7AaaExse1pLOjtOIL+BUfpO6
+t2kZIF96f4fBcSI9RYD0G+6sVEKhPfh1aAyyLZq4fB+5YaEvaKmEmBj5fjoWWACak6T3t07LDjA
n7vtWpDfBqyBs0CopcqzKoqUE+uDGBepfLZyiCu9KtXZnJbzBwtXjvwH0iU2H2SkPnH96yQ1hUub
d8GdMij1/QHMDd78wkq0EjMZqR+uIYvLm7KUCV+pXJP4T7So3+9EIIK+D1mG/xqPPUG9stu7lt+u
fGqUK/A6h5kRn3x+U6xes8pCC546C26OBI0ze2V7HtKacdwZPNIPvAIKw6PamyAjDm8I0jO8oBvM
VdPTdLEHyDDBCmsX9V/QqLbkZaqCkpe6LrHf+Abb1R30yX6HoeCzrUvK5m5pN5v2r+wS6r6ioqXy
bVBRm+EP2BMTipbm6OhKXa9/ZvJD3mrisVK1AUJkAamo6yWc+z4XB5mGn7oCEXkHKAbwWeoWcwp7
4OakYgDCFRXtpY3h4s7uv57Mw34Vdb9wSRLqGwMyYnGhE1Wf94ej0CG9p1eqk74e+3tjxIgN9erh
22F9SEjvtHb41xIpoFXDI970PT2yIScALxLcSTIvo2mEdHJo3RF/Ft5dsJP0FGfPmCpm4nyDHbhD
sA7Jz89cWp6dNts1vET/AoF2XZAQYDkFYx7HBNxL7r4sf/qRUxsmzPNc0s5A92KhPE/uWk4JIJHq
5lfM64eDbtDUoOKTpg3bB+tRpOXeCyxigcD1mOqc1gHhj6AkKOrwOmWFtzZ8TRUN5CoRV+p1uM8U
Or5+mc0ycEUmIX3wHDNoOD8om/33ELF+Ikb+a+wk+yoewF8HNxxzwCnt07Z8vM8l+rz41YhpAKJk
PsjrdfVkbfFGqmMy5BiWRxHIm3jaQd+z5N7tu1oXulK9eK191czuv9bx9pKcGvZZqBiZOs3UMkgU
qLBkOWPgzVsJaheo43THox4WWbKCrGSwiw5pZHnXjY456CJOX0J4cVBKHx2aB0KBWcaA9RkZFxPT
kfuzzwukbnIpAwH2buFx7LlyTMK5OnxAZyKeJLq0mbDxXJbxLopb/eH0YFr8MjgmQeCU61BxXplT
fJQkPofKikZUA6XYDCorGQxgayZcefc3gG1KXfuc0qFK00WZKI4qp6F6iGQo7HULIRL86RhUz7V5
2G5LvackICGP5itQWthXS01WDUmHefn+ut4Fka4ca+r5klqJ3HnnIdGd/4eZsBf3ZK8a+CCzGDpZ
rqX3GJ2XI/F3IMlJGFQzZwwPuM3KkqGpqu9k5BqI9uqJIEThUhMgEwMV60OtFqcB1uBDg3HgCDft
+AKuX070wyl7NkCibMMCUMVuABt3TDFryJSwiGl76bZBYEgxkzzAO+vHZCwFEAwH/SkcpbbNPR4R
xifBb83SmLRYSZ47wR2k7GvoHkCb6AXo4zfjjgoV6yMQCPjsOJncIEduseuz4DQPt+RAv2TbjVVu
Hwn/9UYA39YotBUzGJwXTXy/8Wy+pyZ5ZrAzT5SbIJ+oyNpc9bkgsJQsVxDt2nclQ57zFENFJmhO
jTY98jivAAV9actvK2seUX2KGFDhqLYInwVLRMz3vKC58xuPcIiiyNicM7SFJvIvYt0AbgGe83M+
ocpDD2uHhqR+virYPd3uAWB8THzhfyGZ4TacL1NMCXYlBIF9YZyhetHBXnNjgfF8QXDVA146eR8o
QA/6FwqZBFpk5iSRUMTpaJd2Z/iC2na5kC1IZxOioxKwzudDik+tlUTHV+vhQOie6VO7My9y7Qqb
pOy8M4RGcpzZup4GZ2kKJG88DnUwhpbtEfjzPX8wAOmA14/T56RQnRx5g2rZjPAzGY8jpjL3gv3B
Gk+EABsFtx42TZNJhZZn7qkeLGdIBqNtiqORasOh625HPYIXyqqEn1hLRDTjtixklx9bWTpwpjvP
KiDIpL9uPbKoSUp/Egi2kyxIV5C5/zL8d40VbuVrdWOofWp/ROEu2+9QxeeEXCAtinh5HBMIRh7T
IOGvbU/Fm//ml/rYKrcf2WB4eLh9/cGpLlOdGzj9a6zAgy9Ff73IF6+/5hC0GlhcgobICzoZDoGa
xH623rEaezUB5iORLTncLpEV4W0MOF3PZllfeylIwh8YVfFqQMReq7PDE21skFAcdSX1SYkE9uQJ
1asYx8qkZi/EZKAV+5qA9qj2z+besxSQrRd4MUnNKj3FQhTfD1dF9ZR9yHXFyaUGiFUSjtB9zenj
wg2LUXBxI02o7xCgJI8MwVc/4PpjsUbdRJgZwyIX5TzrKRMZTyR7hBUEOpuk405e3y9hoto1OQGp
Lv3MEqaStJIxjpcU+B2w5HB1/Zi+DmcHgRDRgCxQXcTHGQDiNjc41V8QJhztB/Oxao3fD/K1X2HE
E8Bkj+8GNg3BVFmG2mzwECarLQ8OqFVafJUZ1OTAEPgDbRtZWSIVg6FCwydcIcurbLy2KvBwtzjO
ign4aSaFrNxhbaSx5A95PaI3DL3dkLyswWpI7UwpEuaeHB4puFuaEY+vkSexxefDwWjYH71vcGwH
zRoR3ickc4nIAYesQX10pQ7qXRVg6oIvLAT7gHl4W0Cr40lj1uil/yJTxzfQeux5irxuVc0TWHmL
Ou2FFlGASF6eYJJFaqT3xvhqBKcnPpHpIP7vC3QTxDk+9ZjNtEBggqgchUm7GptM50WO0BgVrnZo
2hOqfRwb7E+2NiueKIL/lLGzGvuQOM6t+2EKDFmPiac/LCXa0fV8wmsFNbOiFUB2xBJ5fSP1kw8M
FVLBdZOXx0w3toJdD59g+VBte8fkH2e3sYDPgT4FelnTW3/CxNRrhDnlQ6XGJ0AFqE1RBI1N/nmT
rXq2GVto9n6fBkzNOp0nWcfRgpaRGDtRLeIplJUKArwQhXhvtL7b3r9ylstRmq9j0ngeMvdAnzKm
HYGhtS/fvU6LytWjesWnhe0lqqtAeiXmcgC6dRPSdU1KRvY5ly1vrqgHtsTomet31y441z53TIZL
fRSZyE0oCBDyed4G/4Y0lJLP+pWOAdj51EPD5TyUyLILny2c5p6pOU9muHhfgZ3o4xy46gbyOUIg
pKtK2LLk8mBRAt9nMRysy00BIlJ3m5lpIIvrl+puuBkXigSGtzV1XcI12I6PuN+rgxrSxTp3786N
qdeIQ02ggNTBUKiOyl3ziPhvIizfZZlv7Scnj51af/hnX1kBQpW9quQbddZn0FnY730GPVKlq0C0
JO4g/6hKeYBbfRATbMLERWm6wyLxhbBwHPSaSPPlFessrVpzYFg2g9ZhAZNnhkoO4h4T6E8CFt6k
uwXgEULJPB1PJciNxMqMcW5ocBlt8VEnkC3TQbegHoaQQ1KRPsJOu3zYHrHwxZ5A2cmECdbqSvFU
vCwHMVG+5horrYD2L8/V8hBrmOir5HYTvi68LblmrbiacjOFh9LyC/4NFK4AjgMsstT19N5n7u1b
8k5d9zP1zxL4NXeP7O/EeYYRD243VCQhhrpl6qII1s6UW2iB5IODmBqYACNlocT1kU1c8NYlZd8p
CbwvgX8BTPaahVvEusLg2joaLyCp169VNdPhpzk2IEkj07Zd/98yk0yvNYSn1jbPm4pl8dJDn6/c
Ic+zH+Hpp6ldNAD0/bygJp4fWPo2D2XkJYMGTdIj7zmv1yN0L/prsVUQU7ASKMJwg+iAUcs/3kwe
GS6MU3KC1om478Tzqwd0FS6mw9BxCfZCP/1tP9fiS8Cz3xzAdJa9gJzXATNRi2n8SzpYJlQadYQH
RvXMZmpjtcFn/IO5Fj/nzn/o3QFOdSgjCNU+uNh1poxpJUtT/MYbqljTKyNWSvX1PmUnQLvP6P5I
eVAd76UQgmaqwY+WhLVzPQzty55+KT1oRMP+vgjLB6mYoH7r+5Kt+CCDPRmmRBSvd/KzOxoII3UM
V6OYDPt/sV9y6+eQzTeh1hxcu9cQCNA+wQvdK2HwVBnL25Eu12hvCZ4gT4UN9Tj0BqCekLszQWQ8
PwRSNmEpkU3hwm0Hm/1TzMUoAjCf8kMg4p29cwBn4LJ8EH1gBik5RFn9Uwvm2814XI9mwjxaQB38
Wzv7zF4B1Fd/IlMYPjSCi7g0m8LUZsSN0/oCAWIU5T0tSDyAf81s2hHauBF9NMM+tRj6SWDM84vO
5XiTeoPc2AJ6wrHFD22DUc4h4KBG9kFa6s7rlQR8HDC+/X+GP6Z32srEbwuKRAh962ySHtSYMD6e
rOdhdn6bAgA9QEJeVfDo6pu0axkEcqYxvu/LU9RP7P/A4bfrDzDTumUa9tRHoFyhZw77wE3bPMJj
OOfAiSfuT4wpw9C8r1o9b3KBlj0carZwQAzHrnd806OI8pxnMKsaZxeKgPk1E4IzHrJ9D+U1evtU
ylOUnT6gAznLsu6C0B8HkwMbAnznmcIZOlQRphKv1jLfej31FZGktxEV+CT9pzrbcw8+FTKME51C
TI2lWmmm3VRsLzyMFeIRb/tFbHUEwQmEkMf6ghSe1+2+jS36I4FvnGPLB6G8gp5J4cvJ7iMGV1ti
BNkiwjZNlm0gcS0H04K+KFhJSHyE0MbIIJtNW/jq0FpJK87A+k9xVcF9X+FwJtAzST5aM3OMG649
SZoHN4E8SOfDe/l/fCmyj9i8ABuvJdlcdYY3gGUxiiPPGeHqilPxdAwVDKz8rZ25ZlN7/ABZ+o1k
HraqTdONgG3WdH8jJ0BIk1qgA82nZMg3GMWy3c6fb7YU1bPTAjWigtg5cIu4NQ1ZZbVHLsN3GgDN
e/puB+9YDhbjH5rIqXDOMSYRacJYImtAtQzfwKm0CFkUVTO82phO9CjpdfT/mtdXh7r5ZpgPxsbu
fmr6qAFKoO+ZLT+LPpaq19y/b7KRT2B5Z67dfNh4MXL8d2nPxbP/bRT02xiLTtBZ52xVZANR9C6w
d6LZEZX81bSBwtBGzikg54PizAudT/rIen8d0XBMpCbTTzNZS4TACcQ4m21gyJXcSY8ij0iwLs/F
SYDx/FRhRiR/w7YCtGbMky9ts6opKfcCjHf5/XSwRKuWTKadoJ1HsLZx1e4vOppU33iURffEeuce
rHXQVBAXfE/xwwqSYGtg94zgqXK4KaKthMh4sDOtWu7U7IFE0mNUXJLUskCdma4DhykMviMP5SEm
SOjPxiTXTqVotMu/pIGXWmZboE3WtQZ00NB4SXOyOsFtTW3ROQhAIX7R85eHId3qTgozXR6V/lHW
0BHoq5vCXs5gSzO52UwN9aJw1GjbE4RdUQzRXRWoUbLr/Y04wTDan/g6L7vmbWRArx6IZL/AYFjz
LaK4X3Lt1F+zj2EY6gVW4ZQAz+WxaBxoZ6Epyrh4Fde8N7YOzi48rNSUgSeNakKOrufKuAClFrmG
FtQyD4D03MGDQhU9sXp8znrhRDLBrcj1u8Gsz+Bj2vjAdVfSs6mncNf6vHIzwCRZ+llhSUKE/173
nHMeRN7Nk8PyODJze+t9nU3F/yJdyM1m/IPFuzfNq0P96VoaXWvvT9zIodqa8PqC01KzfSm7KQk/
bbKf0JwwEeTcqv71zG14jeO71tntw7l7C4nzdJHc8w3t8RulAg36k/qzhfoxPIREV9cdYeFDNAs+
hlArk762Gz9S/p7ernMfwdTJ3NYDS6fqa8Pq83OrMsxQXzHUNs4+s8k9D/ozUj2urziujfFa0gWv
ixoP7eGq2oT4f+uVzN5KNbTDZfKZ+9AiwtcMU0jhd9GxioBpe5RDAzgx7EXvssmIAbyZdl/wxCBd
7BCKAgVxJSvgyKlZaRq2SmcPZGhifZ85lLr2ldlzn8XwnLePrj9Qre8hrFwlEbdf4kwbay7hPDlO
9WkeCOIJgBpRyFrwYABU6mPMszYCcWbrF5ltSzbC7+eIrnXZrXlrk17H4WeZXIUYxQmr5B4eR82t
5xbR5JQgIP8RtBi9hxgT/A4GAq50vM+lnkcLUiit2bsLcSPQ1uhQdEqYcCi4Q0sJSz+u54VhKrED
csaGtvoqHyAyF/V7eMj+BmE7LWDV3I1Lz/gJq9rFSn9osrvRCgMs0lf0fTDT4eQ7uixYoM3Om9jZ
7DFGqWW7TXFhyVbzxxbw6EEx/TwIg+dJ1SR4w9Dv5F8Li8LvR7GnrEsFeP265rEDsrkt5OwHmcJ1
PNwvJc/hHuPuLjTUmF20ZvWa7Jo6iLDzHgTssnMTbCmwSt7k/yBIqk85I2w+tILmcfe88Doj0h9p
meH9E2+a0CNQoEKzLc/lnSrxuWlvvk5UiBeljgIB7V1KO/ytnLBnSEQHtrt+8oTonmGvzsUaQoPm
l65zERmBCMVjHs1KKY9MR5Rs6d8wPz6FfIYSZjDF9xWSjQDXEaRkrRRnAIKR4qXc4InqzV+Z5Nh8
QklaECP7t+tn6G9I1zE1mXNUhXk3xxr4wv75cauZ264s7XZ+8lGyvHdyUJTLVSU50c3oyMtb2dCr
mzLbPbwA1aabOCGelYY6C5gWvCWxZN3u3/YXaqFM+kpm1ksFq2nYN0xfB6fk/qWSE52+g2zEX95q
t9FP5xrTHmuiloI6egxJfkOJ5I5qe/XB7/Tf561l9rPQpcoQPcpQCoZnoYZqFkdH7BG4uPhwGXad
Yx1djQMndFoIjlSzXDHQxdpYrVv6/QYDWfUH3Br41KigjvLmazVhz7uNOBV+YTzfMWeyhbXRDPsK
/zNctxaeH/5uijmdxEU71EzP2Pr2NX90YL26tZX7O8V+ky2G0Je4YJ2HU10ev6vSGIJvoRhBjAeU
nHJTr24yU/1j5784u/Ox9HrQ5NhcZyDEWLM0o5lVqW5DQlEzyislTBxfySDWGAHwEhS8QpEKRqF8
ZMkJ03i2uUEPKfORGn7gRUjUIbhYBHEO8hEEFtWXKOcI155hjKjYgV7xsh+IdZ+WUGL59t0TiWNt
Igcor6YNrbFEJ+Up30sW5oiGO4ZMfgjpJj6qbhRYBOHJXTr0AhHsl+9S8AUWktVFk1Os98uTJF3d
E+iYWeOJLDmc8aZb7sjWA6u7mnZhZ4s8Vdzz929NbxWRZhoN9HqVhN0Q/vmMZKjrQIk2l60FIdiq
P8ykdNlJ3HTZUpU8/2TdN+DplXi0K1h3U/d7Ls8F581fcIgugd2pYfhWjLSNMpAA+AE0D7t+RO3S
BU0W9jj+um7F4vUJQ2099IxfuhGZaHitql4WtgfV611Gl4hNb0GVHormdQkk2MqpykONIoq3MSWT
IL3qLmKUJt4Rabb4VFkWIyfR2/sidNIcfOLtTlRwWAZJ7TxP6F4VTzlfHv32kcfBX7G3Iw0JTdM9
SwSRv/CB2rDi95VUKWMdZ/532VcZKgkofKk7m68NT46yYj3NbJ0z4k5aoEG7DMynd5hoZKlPAfGu
3iVrWyv57lQ/oarEfrhBOBDNu+oPIGAdUOWAOvpIj7NCMFQUrV9nJ/Ak8U5dwXjYQn+2NLoB1pBz
XJ6C1IDyl+1OggR6rM/8Fv7T6WYw6URHi4PZ8EDm25uemOaZjRcVUw148wzZNGumAi8I2vsIEuSb
2c8ZlEt5r+nRL2f6hYYTFUbtMNB6ti9+6ICRblstGqL32tppRCHxfOkpR7fpubfK1qVBav7OH9kH
5EGsFqGW5J8LIQp4tHG30G5Fw5JpclnuC7aC3ghwdjbvkWmkSU183tgosICEd08iOO3C69cZ63eY
Q4vPlee69cWlZVsMHghCn6lt8fJlLyBp9gGqoBvDC5lIqJ7JNdyRV2P71hxdlNHC36AO6QvSdXof
pHuzc1ULCfOLF+nXCMFgG8YZl7ElWnGT7qdraIyKrTIYQ1/CpFHts0d1iOTU8RWyA/0bjfuK1sJQ
CeNlhniXUormiToQmX7FYNTpUyvgami9Jm+GzuIOFOFUL3bwbWmWeY0+wxQTYP8KvqO31QJt3GPd
MbEYFIMzR0sAVLLAawyajlfmICvhQpqN7fv+5I1rxNOpvrTlJVXDPXEvN8R/yhigrQmcDiEcw6oN
6hw8rqUrREal/cvHIO/tpQin0lD9sz1hreawa9x6IGjuiwR8Y+GWTB4VnCrQA3BLod1+CB69Xh1Z
gDidCOor/b8sj943Xkjxgj2wjcqxlYFcoxyItU0tNqkjEv4ylHDINjDgIazAfy2sDdqmP/BZVygi
MqwrmDj3n3DWfbJjv/csjsoYN8c/GK4o+vO2gX8pW1KDPWS5bS1Iv9qkMSND5edFpgwWCbK43Opd
ps6xjkr7cZn9axwZ/nLfmA40iXjJ/lmTbQHBQcPIh7g8BsYzyzVHRRJ5KRps4K6dJ8X6vBAmHMbs
jX54tZM7WGZ+jKrXBw9gJBOHNrMR9FzehAxLtdH9Q6FlV5/my/IRVCmERpJKC1CXlz0Dq+4rdod9
f9p4f3r8uNl8NAXJy2Pkobeqo31VtnRu6GFRe0F16VLn+5TAwFKuxciyUaEk3fqIcea7tyRs3IWj
migUrGQagn4i3OIzsjOiNoxkfAWuPCCg66xhEYZoCxS106ZLxkjzO6K0yeB1Fvvl9vy6s8UEtxex
EWbI4505ZJAw3TX6EsGpT1eOO4jfsImzgndoxfUkPU9TohY1cSVeQjniH3YUvFTPj3Q/skmBfu2Y
AAAFe0Pe3eET/xCbECj2IQ+Rnah0lOCyd9GV9A0wtf9amZ/omY5gnNV+zT0gvuLK8lNh4EK4cFUz
Gaq3auDJpD+iz70jsL+vQ+Kmoul1APKMbcJQwDLXlKkjIGX/VzxYUi+Og3p/ArsPZUuIn5uj0gWM
398ieItaBDX3w0wbMc9LGXIoglMGK/Kehp5qchoh80Q9C5MP+h+Pwo7qoShaccEV6cCWsZSZyAfz
FpMQ1MSw8/3yJGTfygQcFUIVa+R87P9KOS0UltZdNWQjMTsx4PgLSwG23lN41s2sLjKcwP5NnxtS
Ps8g6IdOBC1ZaUz/3IAbQup2FDW5XHJ1ZkVpLBiGOAZvEtaDLeXgzv+0JOt0JgTN/2a9pygSrxQp
PLwqHkmEldO7dOXekswt3nG0Ix+u8vJeuahLw/D0yZQVOpzNWVnDuMwoTk2AmG24CkqZD9TP+QtC
+xrg6lrqTGBF+LQ0hUQN1ySVCdNv2OlZWF3EjgG6+f0Ln5lh9D0cbtPfN3oNHpWL97VbePYsquT8
Na7aj4oNg+ggm+dMp8ELj/W8Dq1G0fzgneVuxOxExpGcshEU1IMSBgZsQY4vRYpbZ/IukjzuBFEG
nhzW3Q+j0nardNiBNrXkky41OWnfvmJ8jrJPX/Abb4vaKdevZAvLAEJlGGUoaiZX2hhTcqT1xFZz
uX5BZIwIXitV3Eh9oUIqkMoCMBIrolp8gYGx599aYKJ1xkp5DHyZqhWU6LpZLZZjgzGZUTqvVnQ3
XF+peMkV6XjhrwmTYSzKt8bg2gYBFP+lj7TE2UAPBLCxS7q15DTG3nHQhnw7NhzYQubNliMdcbg8
p9Ay9IQoEganTbet7HZqmfAM9/r/AriWD8pRMKAjq3dR7KCdt5ToFE5AquNQUEhBUIymLkgiAuOk
EtUTkQAZ8k+88FzPcw/JlVZWCqfggol6pCqQrqtFcGrEAiKu+8jwBGhfhwAGlLsw1K831EMB1b4m
RP9ND5ail+ogQypvlaoFbzr3hL4wiQ2z1aZ7dj/2TDkBbfk2UQNAcXDz5FGvRzf7al9Q0KFaxSAV
2V8Zha4Mc6q/qRNyRZLOLf0tdPyCmy250ONFAfU3AUlNSJten2qnzQDF0nK8YJ0IgQbMiaDI+/K2
lT+wvmiUh/V0Iq7tbyvI321UbsFsKL0C7U0XWgAY/3vTe2NpWwKRGaidz8HlXSf8y4oxOdbrucVi
+3tBHqUfFUiUT/IOMY+3xu4nLLsP39RjiSArxucXTw+5XNQbQXClTZPi3WSIG1Qni9Zk+EiqCUQg
UUcWbem0uphrQNgWXEoWZ9RAVdRBAsaaWwTRU4dGY/zzZtjAX/PARkL0qpngBh92H/G+tQkC+Njm
g0tYh4wLhGejy7U1zyvriOZN2PVeDu/XxrV7bOhq1u+x+pCEOEjnxXF8rG5m6h5tUcS4j6nnq2Aq
VxSWwjNFd5m8rLMeUEDmgtc2g7ms43RY0JiDzd2c9bIARKio1wrs9n+A2f4BKxk/dqrKvZwRfyTB
6EhK0TP3K7z9sGVxDixVk/7yNtjcFA9CR8hAM/ViIc4Dm0dwDDknIJBAu4BtlCVW8juv005vRmVU
nidW9C9PM9W1DC48wH1CC9U++RsdjBnC0Veo/WcbHaFQLZaj8c0ByAXFsP5coAX7zcwC7NpnpI90
3tmu/9LVsKosltqKwDN02+ZwNfXuBZpUOe6+7z7ZKKWUIJZjuaKT29DGApSLter9amkZBXNti6gS
UL9g7A1nlUmGXZrVnO2LLJPjaDbwzD2Yirt5Zl1wJZFx8nck2DKRenXsDeflsQLxZmajhJpgQEcX
Ok/mkvOkkHgkIABL1ioV8TyT+BR5GlbAVRvNdKcye3lGYDJIr6lWwLmUw+PTkkoKu4e4NLiMtNU+
HSvhM75P17q4orW0vxwLRavELnMsDyjaB58dJhhT/CogMkD3C7YyucK1ADl4rNf0qDTqj0J55jn6
HOAMNbX55MA4UHkqaNhgrDyC04LAVg7N3Hlx6KPbo8ujc3+knqKEraunWwa16dvk8tQsloTqh6tD
uWynw9vRrMbOMGQwHx91qpyfuZjj173rw4dMj1rtlt+z13s99RTwfU3AHpIDyvbGV0PKI9jy11um
i19ETg4rMpiNS04HPfWG/kJ8Jx7WP84TpgKils4UNUs0EBsewUpi8x5IwirjFpKyi8CmcVgbaxL7
/q7qQh4w1vPZ+Om2Ai/uHnxzB6gLS6nhGoAe6wqld10ZuVymCRAXo30sct1ZZl7mD4Yngp9BdK8M
MnsAPtMJ30RvKZTOnoy/MZRjae7DCSOIBeNzc+dp+tY6Y2P6k1+U2ZsK9XU62EzrxqEqRktPMJmB
WKO5s0j2I/f4Up8MzZ5ZBT3I/1RqtEXmGPeVsfu8MCLwMm9TSNANyGAco7BrcBhcNRZFyy7euIm0
kfL57JKHzPB5j8ANRH8ZJKRM9O/a/Je2+MyueWgwzQo5QM8TnvVTEJyZzeR5JgEL4ZMkuNBoICQO
h9r15G2r0047B/21hYov0+o3Q57GBidZoXwPK8ASKmnwrXuEA0+KZe0W1xeJzi8krkOg4L0fDGeg
svzoVf1Xk8G/oxS4sSbDl/mT5hubsU176wOKAbMdE9lf/KK8ZnF+h6LWWVwAgqLLLkAZBgT66TXb
uNcuv5Kt9OQ+uZaI6sCgp/OB2Haz1+pWXH+07INV2lwtnw5h31Bu/etGHM0ojTv48Y4O4Bt4TW4J
ZSdkJmrYwovO1x1tfLMnHEL7EY7ntJ+0W6dWrQnz1CWEnZ8dO7UPBcZGbZMsBlVHkE57OafmDTK4
OREwHIGXcfVfZE3JcUi/oks+4Z+RP9o4/cvRcOll/dm0vWuh+tAVFyRnLMBO8GLQoEGteohz3xRP
GyJd4Vt5JwP2g8SPNDN0aOHM2DwQjQBvyOT/ZStEqjU0xEChJjObj7aazBIiCK8IHQuTf9do4g36
nshZV8UJw+Yr7iwtdWPh3HLTxdSpIIz7RrJm3RGzpik68MdVutf7WvRhRjH1PZTa0NHgQc6TMBCG
JfPw4N4XhDwnQqpQt52UmwfKkrgx+qVjeLFUxOJ8Lk8mFz4HF9C9ZO7hBsRiLGdmB7mi58wIy8Em
CPlEiEuh3wT6WezNukXfLQUxQlgFoSFRWWLWIzUU6TgKccGtnwXjfdkj4UDvkzds5gKLFIRXRMvQ
7kEKy3ryEAfSWu3RDWegV1cX8QmE9gFmETfdiMWx38U461i+U7yIY7f4Y12fcKapTXD941BWbj0c
7sisjSF+ShcBhfQnzFaZTkfQLztthAtm/2xPMDuTgPkNkWevbqYbzpptp8CQTRslKI9dvkzEAfTa
hIHBezDeNuDeWbVjwRNeFDpXPG90Y5FHYms5/y8AniNaerhyTdeCjyq6dtcYdJ6WNPKE5z3d6q3x
0XyOYtqJcKER9D9f2x+mLh2t+IRXPnKFP/mccoAWsGD2eAfNux7cXsu6cgYiOlQIVdnmkNVoK2V7
G84NxmnSam//M1hyBtzrH3jWDIjkfLe42nnyVDs96iVOhPqzFAewjxFa2LCRWq8ydYwdZetfc04H
YnYZcwTxXwnBXpln6DSvITU9yfL9sRIAysC4Ps520OHntyaoRHPDg2pbZPmW4EZti++bLbugrBHW
QWfKTALqyMAlEV4fofBGOHcqCHzGZ6z6IuG9+WKM3I2tojuwQTTpmf3jVYY8ut3atvb4oXGlRwqS
/TC1ECnU2XdK50N+tHy1v2y2VETbxGpPtF7sOZexIDB/jKf8ZWmcMl0VRHP2kN9y95gDwUMk0nvP
eVUYwYZDj5Whc1bCR/cYpYvtYpdB/unPUI3i9hZISVRQAuC9/pcaf9Cp4n9atZ5XdY9I1fV+3EGB
C6bRipQ8pp+UdRaSANDExQ2QLnLAAMiyVaiTLmz41PeSiuJoyCSpQZLOy+KTzpeWYAb/w7vHDz+0
NwpcG3cz11EodsCGJvGwVPuta6k/9dOni2UBmW2ft/GcnDRrVJKY7SazYw1eBR0ONKwUNz0dpf4L
5ZEbz9E+FC360BBGjFLutUWq8Ey12itcSf27AWt4YUPxVDyvUQuNYau81uO3uODYKUlr1o0yuWIq
2l0RS+isGfUofTADXjAYy3zM2kZKDPIXdpHRGr+/IWOC+9uFAYTME7uf9n8CbTwYctAsBQDR3Ar6
2Ev2D6wEVaAphG7KrY0wnm46Xy/gjAo7RVVZg9RLk84XSw2DhwMhfilb0CRr5SvFvGB6dNqwk/JL
0XjJzEO4Mf3McmNR9ykpgRUw/0k2aM4B7Uax+4SiOR+4z+hqjscLsUwnfB/l5N9k6zCNxtrUR8Jp
nVf7xQSMGPQU2vlWdIHOSm8IPZvIkXLLy2fqwjjXumxca7Wgffz6UVwkvGu1cJI5gceiqYXCdQnY
e2LsKyzpFj8bKEMRNQSmc22rpNwWGgt1+TOfBAExOe0TM8Mnj/DG2mL3W2FGS/tsKGITd84tv080
QAIvpSL6gv5KJh6VDB5Wf2zkeIMgJm92/Peqd9DHKNTcDtmG/nj0cbS/5rxreO5l3C1n83xgAJo0
Dw5/8AW25FD2+4sCkpofTiLx5ZxnWSdhF0qN8Bi694o9Em5SgzFZnPUDajFkEpJiq/+WQYnDZfAK
m+GGk49wb7fKxMMJCkp9x7s3Pr+xYMidDnWi9P6tCEUf0bi8ho4pXQVyHF9CqY8Lh9LkkfQmlZfo
DOZUDJMOSanvAGrL8i1gPsdzf3E6XFMpcQDFNqpkAycs1x87SlhXaw7s8oOa68p10/66VG8qfFdj
jnwhFzynX2hYzOQUAytvm8zwRQyi5UfQZ4b69c+m8PtWe41AWIG8jIA/HMEYFRQCYy8T6bV7NjnE
NLxzift2PMfE88kEMgbc448sI548+BHSyyJ7A6mhqpdRxW+07CEiLWUVzGMQLQzLvgNhjAxgW249
9uzLXI/6Xy+KcU5+BGoRqGLAJjF7WEirhYhoA1LJMna/RZDrPgoqKEiuLu4Z1DppAtBn06miNED9
JtomDQirLJPwcn0Qk8mg6D03gWQBYHfJRHuNUfeMLEL+fcd5GLf3TlN0WUDhKyzqmHlGxLiTih9H
jKD1Z0efDFpWen3QcxjE6y3E1IFG+4pCKI7iTCo5SnVNqKDuMb3bO6p8eyHSlEkAztsLRxJW3Cnm
zgKx38Y+95mZ+AcNBrH2aM3H6xE0GQyY0JmY5Yyp3O+XqYsAZZWv60TLHscmEnGlMd9rCOYc8dqr
3V1dR9c7/EQ1uQmOZaw45ObHUO/MD5Ojis2XRA1VjzPbI2P2+Vgj+APuUeS2gnn6Uungl9rQw+9R
9Eaj8pS0NfIEw3UQPg9T9t6okMlMjrMF1LbllO+KGeIkeRcoa5y87+pWbm/M9HAb8OxGLg2UqPuI
3661nKPNovE9lyZ/qHPnuIqF+VIk4TiH6XYNFNRenNakf9KL7/yUR1TPcjQhJaKlNnWFMyIs46Wr
Eyl+w7B+RvF7vtokODSZiNaaie5MHceMelnd+8hqPfY+DS+Gj9WbLfOB60pdm1Vvy7aKtM8LOoPa
yS9PXqPSO+fvf8poeLbgL5jfgxLkdq+TesdWTqZFha8UhL6eNAIMj0mOdgRoMgA3j/MK+8Ev8T+B
/wQG6EpuKwK5c6I1EJLsJW8iSbUqIQeL9jZtiPN+F8MDQ05cSZLyhkqtXQvu+Fdc1dKViCVOVMjY
slFCfG3z39YLcLA08/eULzJ3+Ph/P3I76sXB06qOhDFRTK6j5aHx57q79fMnpPwg8UD1cnCO+wJE
GwQtMBgMNNqVBdh0pZAoQt7GA8cDtllygrTgxptjtfX5xx5p9OF4jTucwu3E+8+rMA8hqS9SdsK5
iVuayz7aZHytjYgX/SsSNNcpzKLo6cJD4+x/SuvZihk3GtTlEcxs3LP0V1TLgXHFUzJuSla5TsUS
V441s2u1i7voVT5wOd6bMqJuGolBHl+b82YY+lqA7d6e8m9aXJ8bjUYvQK+Vj/cLgIgrEiExi8gk
SDJkIGVYRUvapo2ZJiqbEQ6qfi8SDyNrGFGxrSWbN6UiaPXy3pSeOh5s7x2NQxvxY9L2XX8KVGRu
gB7vr5RekwFy4HEBry3s8kDkbccvTMAuCru47Sdw+CcWJTxOounxkmkf3z5JZCgYfyBxhf19XZSR
8iw9lsIh3kcnbrk8vNbE58/DIUdm9CYncyCHosgD7ABAFigYt3M6+g7FVZrMfglTnvTBic8WonTt
saW+T1wz1Zk9QLfIi2F7xY/utefQiFA8T+BmgywuLQq5a02CWydXEo/rI5pzeLd6kaUPsh0N129M
C2BgU2RWzYPKGqAuL3FVSDBhgJQIKjg74WuoIK50kDNMJP0qMvbbmBklP2SqgDK8NP1NHGmVyUuw
JeSPQ8FwFjy1qB9DBjqQu/0g5c03TVflhn0m3RPhagAdu3FzQePvgJ1GLz8nSh2P8E/qDDFB/rPK
Nm4DA0qJzsBbvK6SpAatNRmq/oDftVEoYmSLbR0oUCzPKGB5SNgZBimHpttT+RtxJrtSZzdu83ld
Gp0xuUHJ8OySvDfQf7x1rFIdCqjHAbo1mKvxnm2BkrIkkhoe0Igtao3+cNfsY15851Qu+PZVIXAx
GlZm62SyC6PBiCC4WI2SeVCcs2suBp1qJJBqVBUSfLycB4cv2BjEkL7UrMKEDmakKeaPaAkk3Tvr
in3QlJL/xMVD7UVkpuftfkVDDALY0hVI7AxCOzJpBkeBby1iKMT3oVl5sTHicMySX1Sl4o6UyzV4
CXvdrPZCu0q6TVoQR/eOr7aCnIhcbMRdfIzXs2/pYsgxxzbL/9+5WhTSP2NJZmt6Tmk1kb8+Go2W
IcQ1c42dvEHyR1SpFG2Ljbyu3awXA4cTTOBnLB1CNtl8S5m9d2+LhTloGmQuGi78O+FbmwzACBm3
8X2N/YHlLNP3i9HolyMfwhiJsabfNWLFaKK1Uu8tv8XZ5aTgw8eEu3tPxHNxPNOg3Rzvdg84I7uE
ob8M+XwQXkVkTMsoBo//B5gaGvhSkLjv/1fKtvZWcK4hJ4uXXNMZDPVtmXgkskYl3opK2ispt6cN
uZmuxfmyabjuJFAHOEkG/lX3zO2FBfl2ETCxNUVxdqwQoNOZ/58Ffx2e7aXMalFAF5fuEBLepFBX
FsHdQ0ZHuX2g2u/feYNqAOnzaq2kxogdE2U0VZP2c0/OfKeC9XEE2DcHikOShT89LLRG4IUSFXuQ
Fm4GqbtGoGTg7RRSZtRxXyAhk0MAzg6hwabpZBmmEo41MNK8QMiU4WDKuVIpycpIfeAeWrJJckH8
lz6ya+hUzv1J70cQ43YPaE3+DB3xetdkpCwZ9U/JHC6kuoHPm7o01hjGe6MG/u/9vCAG1cNlH3IK
v59j7RQ/eE7+hVR3eMq7jJloykwJJahQVyB3wBcxu0IFX2SS1iBMaqaIh9UVKIOXjpT/aeToK6fN
gK7Tt5BwcNMJIyusp5dL45YiK5Bkk8YhrIEx11tlC/Z2I4tE1Z8A+vd3lHl/mdM87bK6jWpsFwM4
/DI+CFb+R3F2l4SblJAlFJsCCtJMsmQCdL4bCF36DO4OHP5N56ofFlB4UJ8lGpS7dV9BPwEZqASi
sDyUpqMLHqTlY4qpRBtml4wD3X51TOEuGLAopms/s0DLAK7btQ2sEmuYfBgOn73sopz5l6uENHGO
LETD2NlhZn2tvVCmrNN71D6mgSLQrgRG8uuYoTIYPZ/YNgPhTZ16zUIs/G6U0m+wpS4R2aWF6bXD
MEETsb7kw6Tg8mnBaN7voIhRuEO1IsdYxWOjXTcL6UPcsWICv7cQ3vWHeUA5FgQvCX5lxKLSz5gf
Mt5rf2+qS5lU358jJ54+DIbxejqSxAiCVXRvhNcDWufznj5UeXrcK3bwX4Hg1DLkpjz+LQKZtTyO
ls3uhYIH6YxuD1vxud11A3JwwcqXj6kio+XhGOhCtAmKY8HVj9Optkk5Nk9igFPeiJzYr/i1vRIf
vOV7XVLcF+Xusplgrx1q276PjwjwFbFmArmeDAXT0UHN/oxRM3bQAe8Ulv0TUg6HZIkFpFcbcL3t
V/GNRovu5/zVBLXeVaSAtgQ7eTYP6s/ZrTaF6l7XPAXVjle4tcJt+bxqh+dYPgR4GaaFypGR9gWa
6Y28FH3v7IemJkz9OTLDoMOXON2aSY69K/yBcmDjTuYBF6yZh7jayjBpXrXLItwuzhdEOjNsOneF
uEBxw+CTaH8hC0tJCuEbvIHWqkfB1BIOMkrvz5Z7l6Ph+9MCiX+uyCRmjUq/FOHoFrStPpN/aKFp
fNJAo32MI+cSFnxDb+eQIJP4izZl+lBOwM/yE2ukY5Wh7u3P0jXf4KhO4e9cfxE1FnQ0UGP2ikUg
DXQ41ccot82xu8WYz+sXZjMMB7FhifoN/bySk39a889Jm3B8ETWmqOTwfBMU1osIKFXwXACng0UK
w1PLmPfnfCmveAPdoPhlSfs5eu8LCiXhQpwYaGYakEP0MTkGSPBE0Qu9ePkd6JIOmeAh7wxVLZs/
0nZK4xXfpINB5GjVDyuXHplqBZMKtHnIy7QSw9w0NWqMF3vpiD6CtOY9F2XepawmZST1XY5k1EAR
vuUOGPWhGpPzmS6ZxXXE75x2yL1ZcZKQkAsoB0ve7uTcKCsfWJjCg5vdy5s2lZyqTxZWQZu1CSYf
XIZlK9z8KxcqapcDdwpqgjJljyAZOcNK8Muet0VioJbp7ZViFdxIHR40NW6purBlAF1Wuue9sMc8
5glfcXzDIdEzgeua140FFXy3m3N797GwiYRN7lL3Q6DqdKatI14cNa3p8R7Ktr6bxFBpHjc7easa
nQdOF1SmDO+g5uHWne3FZHOmh/qH1r7QJUBes8ZGMP9LrpT759iKa7Io6RQesqrAufm5fa7ypWUi
lcxr3wi4UXrdwO8UIuJDqmDrmNkeiZpyn1ifZEKOGBXIjb15ZS6MjexuJX7AwsOWdhA0mF5IDz5F
Vnc/W8tTveCwE3Gl93GXmYOlrQRlaIrkLDdxTL0SN9QfPSLoOt0yhnIj/lAmF4cwV1xoEODxmDwM
67rXnskROgGuczpPMC23ZGoeT0+nWOYJH3kEI1gHmLV0iQNv0uDbUyQKewc72Lux9XT8NVwR3bn1
WIbRG62N0w9Q/4xM8TjZsgwXu0+ukMNtS+i82dvfOeXA6EW9Ku+BeRJSNk6AUwm1B4+D4kZaq0US
rS6wBUVyb8vaKRpv3rouSyzebjNHjDkSzL5nPpt4i0Ykd+nqjZmpx+UR6szVFCAyS06XFe7WCD2H
LVfw49I0rHKkNbvY7dPMZGDV/O55OAH01wKPKtqqEcKKuiH8vO02b4pmwGxkxl7wH0U0/iPjOv+I
D9VGyXjG0/A5YKmFcR/Ra1Q2Bj8BnNx+CyMhu8wJYvh1Wf3lGSWutKzNPDZ2Iwp0WGZqSoz8dKKb
uNgjqW2bW14R0PDLT1ZR8dHaFFj8gmxgTXkM4NZgENZgD5/bUo/lzrMQRmATcQ113nAW1xpQ+QK8
98DIVb7u6RIZXurzfrpIkDHITeVvSPbrdft+7zmqY/v+9+u/YkiPwujaZZNEBVOTlnq9UpFIBmXt
FuI7xaoeuxdxljmCwjEeiFPW3SLLUwwYoWGiP/tmoxuFtAWGpllFgkL85fx8LqZ/4urWc+3hqXll
6Z/q4ii/JEL8+F61m2/r/AkfWLfNUJGJC7LC6js6mrpLDHPg1ccHM9pN0sBjIMTA08UXEeGwcu7M
ZtgVl263cyPkF0kV5oQ2xpJzW1O3tDszlPfwtsm7YKnaac8yCwYJlajiOMf4wCLfTH6ihSBKW9a7
pSfrkshi8pe70PsMIkYJaUeP7MWC4SfhSUMXjMLJbsTeaECyHNOAkO9uitiyC4/x5lxQgLoAolMN
PeRtRcXsw9QR6ITIa/JPIvGvOPSErmbTInLH6vc9QsEa0raYkCq+olF8ks19ZZUU2zommOsqIXfM
47s1J+utXQA9mC70BK6RE6j+3cPdlOYEFOoNIrCcI0pouw0fp0DV91czqyM4y6v3lli5abpzj3m/
0tqRo8iniu8utUYrbJs+1+B2IV/wXbCk1H1zU2Z/O7NgQjPPlyF0N9bKBWrFKRYZBcNiLzxtkkuh
PgBIJIXsWc24DF0J6nDJCDB7qldLg/rnebAkhIfRhDQ50uovdEDIZzob7sYaXXd8pzLGJECzgN7X
9TarcZO2yEQLTp/tvD9JLvXqYGlACQ9yMh8M0cWA5t0uIywf7lFg2wzstee2CuveMUiKuj1qRZAW
/NGhyFmSxkFzNEHP4nTYcth98w3kdMADsTXQ0eDPpxvY23b4SFM+XA8+2EXUYHaQ+eSj1LKS0AoH
FxXSBOAzjl6Kp11IeOExB/ydBSjznpHEJNBdo4JD9MtezijESJ1i9+Jx1YljW3fZMvTjIMABVs97
bDcngvvBns4vdtbHA3MGF9IUUMbHPA6x5pCbrOCtoshnvLItjvj6UvcUpbIfM432xawzJRoBMm2H
udpqYiIsOiy5TZS3ZMMk7ZYbL8Z0A8kT1WnB4ur6tvnWkdqlD5l0kWHx8+olBal75EPn6UOQNdWa
9ISfZBJ0d/6CPY/0T8PQE6mBsUc22Aj7qoIaHQ0q/28VSZpRCWTC3YNeIUdRxKZi6e+5jMB2YoAt
1HntzykrNoLBQDy8LMPk3NjHbCiybA1saYGnvv0DcMZAQDGDUAgGQ7+1o+3k/tKjxNLJGcnIflM6
Ba+BBrMi3vRrPZoEkg62bUJEBK+M+mtlNDtGiu1toTtOIsAmW92ZAXNMx9gTuX2xkTM7ra377IYt
UW5r8h856HzVUnFaF8B/jbhay4c13/myOJ/uelY8nFnvCmAvq4OSN0L6DJuFAnwDJ3U2n7T44M84
l2ewkfCSUOHo0IlHmsziZYRTG7B8xmavhmWpehJvyfCOOMULncsPnY5vlo5NNV0YhByh9+ySNEwC
G4yEvZAuGByybin3jSx1+rPn43i9chkcNOMqduPNpGB/pITRT6fUy7sFCG8Mx5X6hL7aQVW4uDyb
ca9v7lsXGTb/owsY8rztImqmVqoA8Y++imkGbJkyxympFyEvl5qRPuqWHDgOKVUVQUdL9mn2wa29
R9s0VK0iYjLDTU7D+gS7hhnZ2QO0377NGGNWWfrKTT9ZS/bQELP9cb7lZqAYdfTeV8953QQ2ZhQI
fE4q41qzWjX6ROde0ZgTZP2Zb+YV8BD/1sriYGrnfuV0GVbhLClQU9/J5cxPG4lqQePvSmf8MG85
fxvymc+CeG3AGU9coeR6Ftm5qY14QJTlg3gFKM05FnntogtjGiEdxrX+z5IUpKRdsNWYIR1rUXdh
rgUBiOKjLgvU9SZdc0pKtOX9VzU86TwMZarjGbdgHvYQWLn23T0H9eoaX+p0bz+HS8lqFKchJsJG
bQ0AktuHh+73XKGuOm4zeok02W7OInff7KBpuZNlddXNv6xw9f37Y0Q2t+fsaEuOgMqutX+lwVff
VAAEmqCQbUPph9cAOgmJ0j6n4l+4wWWCDEI5nA8TQonQSfkmgUAn7498pCIxmZS+msiULwYmtfP/
C2JZ+XlnGUnZ9aLCZqR8vT5v8TyT5T0Q4KRM2ZAHgKDfqlh6mxDid1HNrAH+SBzpW7Q3KQzs3BxE
hxHBBgjOywFHo3NCucu8yQ7Jcxfc8T32g+HH9411CPnBay9qgWAtoSyM5IyAgDKqtyvgLPjF459n
jperwY9jbT5CAFWqlMHAj4P0Qlp5ERUbHF+iMK/EKl+Q1emL2jyY/OzMCZhjzJb1hMJoz7sI+HTX
nJqp5tCItDmq1JX+2o1jU1fGLydgjZqVSoNfDXwJHjk5Hdg5JHPMS38lRRLhM2ELhcS7OwllxhPq
zzRTOc+rKNqkU+BI0NdRcB2eb3j6ndguh8dGqMugzkfCvnF96emdqR84gX9QP1YUkz5unzXhmH8w
Ob2KqtstUbissk1CGjF2aG3TS9AAPQhKxRJMlA0keXm00SjubE2vauri6gDDGE1GTIRfMab2C4Qa
7v6PkLy//7x4hcCBqLoftyrHgyhL18IIdZttsTwGK1b2lLht5QVcAFqvOa9w2oxzNySyb3ufryDp
8BEaTL2dAXxH08lYeKcwmD/A6cm4TrWMCeKnaN02XzkovPukdN53DhlX9GsB/x9T36pYP+TJP0Bd
gqPAbl9XDzKY7bGy80ekOTSmLFQLchTTGF6hWHW1gj3vBB0SffLR0qW0QmAfh/ehzkkc0FsfJWQx
HinZBmIwiQmy4iXVN9isKBHVl6b4mUiEcd9GE9bjPB3XVhnqmTYMofw0dlPLDQVhE1F6W6xbJDlb
ALrbPSsiB0RmO3DxGu6HDPd8rZYw+XCh08yGf2Nf4C2gD4xxD+vjZolYFk4wRXxPghUyRVgvWKWN
cdl6qQiGaAT0+9bzg5Ag08Qy/31P/goV93Pp8W8cEDXXm72/3PgL/eS54mIz874p/y9gFiJ1u4lp
F+0sTbhKLxGMcPTlJOiruRZti3sQpRVE35+8K/nRGfBhyBW7UKENf2HyKQIG3qiP/TO4MuCQMddx
idaKYiugxX3DZzwaIIQbzynLKM/YkU9fOd0fAzulb3p9gjkcy8E/Z6p78Bmn5cV9pY8rYkXMQddg
UaJw+DQ6Vs9BL6tQM7XX/OgxBh32iCZdV7EEqCbKZxNWpXXoVI+2hu+F4K9e0yg5G76V8IDTE9YK
fWDik6XkMan4OL6XlDhP68A1CPbTdQYxd94EOw+CejHpBqSD+vmt+3HpUlnEh+IZPnrKzpsf4VE7
TVZeagHQ6cVfvQUaV3sZ+BDxcsDmfGm7dxjCYMSCbiVUGut4VVVKT67dXPg5QULd4vFmQh714GCY
MQrgeFJmOwDLFq5iK0Sfu1j6SO/ckRshYpEhkPKGtoLppNQttNWGVlEGo4YQbe5KYS4218dOWQgO
/YcIDkt9mg+EgzWYUOAONOpBKPqvh0GZxWgPgi4dBtv7pM5qP+lKx7KB5ey8/Y24kplNc1niPSpb
PurXXOx2xIyoclpLR4LJBIBIpIsCWI/oxD9D5jRdGMra4WsLG603gc27oY90rF7QfplpWsRe1xqg
jJEtRrGBqPNlCnz+XMqzuq2h5iyWYt5f8t5MtmIE0QhGJCV0kRHPw2exaPG/UCtmrUu/Nb9UAww+
mnG02j6yn7Uf7eV8qSbR4c5OQppKgdwgr6++VlKNSW8eh2A21fVV4b4Xd2I5iGuzoZ8dJX8IQGOZ
njSvL7A393X+i9GZL66pOFeL6mBNqsD6XwNA4yHukoTfMI0XsJuxo4dfY/xd+R0QiHLMS/QXC9SZ
KblahoMWL/WG44IlQJTEE5LLYYpgNxbB0xWtmi1YTmLbEUl7DNEH2ctqnXIxBnvbGx4PWLvxLdDo
c/hGTb/xSv3yGgrXfp2Z2NVnk1kHl4tAeBKkvt86IRVwurQEe+Ll2fBK1p/W/Adp1PQZovHSieNA
BHBu2Orrd6EGCbvcfujw7kYAxfzHmJQ++7LBy5zS1nlEw8vYA4bfG+vQRxmEzZvanxmv6UYUi2Au
CtcKfMXG+pGfgs1ybmfEeD8Q1iS5m5kJcQKCSvWc/qOlejKNbilRci/1mkOi9FaWZa4n7KNVzD1p
iDLqM7h9uCCko0TRxiGQl5DLv6siL8dz+PlS0UHYj45EGVP5SqDlosrpMoBvO0yiQvi1/ZlX2ugN
cFfWRXhAdaj2afZsdNJZKgDpJg7JPJDALweHnK/xJQKWrcd0ApreO/DmcILrVRn2dPg/la4Q2ZN1
2WhYA4+/Zb28hNtI1qRE0b+mUK9GuKJJBecq8vL2hc35wi2eto6hD3sgkL7icEolmNy0BJHrwjff
ge0TEP2qbZh4b2Aznd9nVFdI2nWxiOcr+o/DeXTIzmo533dn8dBD3SQ+aFYAuB63oyZOM4vqXqRd
Emg2aZJq6JDrBb9DfHtq7PzMBwohbLn8PwQ82UKNu2mLvlaJlHlSAM0Kjnu4MlCMDqkjWg7JSrIE
LUiyPhK8usaKj7INQzaGeKFn0qS6ygq7gcDENq3HqchjeDyvX+on1F9S46yM0PAKJ87n0qy0pyNh
EsDa4KztYr3nOQg5j7TvjvGNrHltyGjv6XgpdAfvbzUtWJeN4773ADhHFvv39lIL2EbD/V8KQmja
rsmWhwi+3KDIDEalGkYGYqlaHceLBmtWbKBo6HHAObdHSjvkqZZVkBWd0/skYerYFeFDfWUrJ6UY
kK6yiZ6ZEksM1kJduxd87QcpJ3PKCLuF8No+PXZgzg5RZw701hA5+14Ls+K/gJH/JCM2c3hUcDiN
fHN+vBP+oCiCDqSmOObkDffmRIz42DMaL/iA7eWpaLo2ZLlHofOFpH+Aes//Hxa0aniDbW2WPhj/
w7UnW+3G8f7gjzYSDN6fV0ae3eEXx3DUvtfub/BLrAlBbEKWCORqgBnaU12fAHfGzGcC6zWQWKTs
oCrA0jsCxPegBJxOyWSDzWYYiRr8R9+XQt5sbhPpuWHe/RZO0hRhTTcpwJ56jKHsoISdp2sGCqip
+7JNP1rV322azbjIAemCWVEpOyOpJGhq6oF14JPzy7T+2H++p1hy7C2lQF2NBZIchwgUYjIu6AmK
00x2yIzswbpoEHIkSMlNH7eWkynUR5gP7ZV1xC4+R/mF/IL63VBd0Hs9fL/86x01kS/4hsIf1agj
8RA5DN4M/2mu4IQ/O5avEz9thrGQ1bSShob+y+Rw0alledVtIGX/EV8+b1g6DuO6kMM/u65LwYaO
lARFmMAx2/LlMEjb2ZFgtA68T3xIpnI0McKG5B0qM2S0bs/elefnzfYf7dkVp49/b4mC0mW5yBe4
U+P0o6wnTS087tYAYHWFTHuUijbBfwQrMdu/uLxvTJeRr0PtHJtidIeC33e4wT8Ard7AhksflsWL
byk//zOzVnbvKnRwgKU3N1gYS9Rk4m9YIxf2nM49X5hh30DFVVMplhhZndat38MQpaW9dD+oSpUE
rs9/ddeLBO05YtJ8vJqvLySasqEKB2b3LkJBIiRV+nCVS9uOdvROCxqXzwDyeDnBnH+EemPi7vmT
iKq3Wlo6o+fppJnLI3gHBN13pExaHyCKxM9j1L/+hUOCDOvn5eKYd62yyJS8aQ+VkEPXPBAvlmQF
XLKUeUqxPQBLYIqjQqJOuqS1KXuOkztCLRNUlHsNdcwJb6iQV+hcjHIICjKPM7oJ36M3W0rZUu0r
hm1ADuDYpPZOJOY3D2ngAVr0hZqH7gn6xTUtYXZo9L04v/nWcOIgXLHIA8zr58tPBUsK0gwGKu5z
JazIFsyQ9hTRBifDdOVzl/Z0aBeSrVZTW7iiZVuUllhka6nUWQegY32CllIQIAbl6FWi28CfMD5R
RXH8aPhFrxyA4ZohsNuFfITKx8N5eY1yPiRFJOZgu6B8TH/BIhXkf4daxIP+3PCXVFelXjuHI8g7
MVqXGp3ZqXeaCcrDJ7wxb5slBi64Ny5QDfu/497QS5Ftgp1nHCF1+wlTTW4Fb6q1EtfdGRBVj3NP
DSo9Qql9e1fh4PvMlEffTwdq6wL6yRSViMmaIec3MOGUUsFSr6MMHTnR4Pz4Q0U3iyTd0B2aW8AF
cFc7k9PCh5lqBZNASj4GMxiQ75HUSK584bc7LLYViV1awUOB7iOg4jreqXpKxKohMKsXqLxIq+dq
EGW6AldG5IrEMOjISjcFoKYIqiyW+ZS/8+87IZFhx8Ey+88bVC7kGQGdWsbZGYG5YTDH6Mgnv1Z4
MUtopNMwbgDnkXmCY6tIJHl+HSa/cnCXbGJNGnT3Tr+7bETOA1LMBO/R3FuVD6R5KoQctLKXjVlI
NzS3nZUmatSoTd5ax7es8mHmT7YJgn/rvwIKpuq1nLxVusv/W7RluUI4OKvpGs9m2lFvcOGjy3Tz
DulfkLFTadE4lywJuqjhf1rII6wYnIh4YPtWJVpDxmdxUna+7JQ3YAjGhrR3h9UCM4qbiqXjYoRI
uv0r6xJeoScSSp9hKY3J84VKRCB4B6gfLfWU54cqGlOsLEq27duvKAv4/OSxmfCMsIt8Ohv6dFUZ
a+UAPuAuaREChbjVg6ZlHQJreiHIj4GwCdsT9cPBK77O638XN6Ol0+3tBtgx97Qo4EF2d/QDhnWj
cX8kA5I0tIx49iBO6VOL9FM4rSuBfGuS2sKIIOOh3RFrMZEClecVsjKr8vm1nycAF/Eu7OHkGiss
SRqDOuz1o1Wbt0/j8seiukV4skcrfbJNRiEPARsQhawDVQ3K6w12rWxPmOgUBl+xYXUhj6MJIF26
1oZI6m6bpMRdEUHyjnUZrgZpuMBe7x63JJoM51J8GYFsZhqqwEl/kCU4t4Ysu2qJLozhx4stmxaw
OpNNO4taV2Ym35pACHY14AKzQ0qOBNJA/oGGVWvoFnmsYOuypwSOyvuz266DKACQVPHgQruBXHzn
CrRi5DVVWCC73HokbF+VbhvVQBZqcP+NOM4eQQEEnhSpiO2DyEeZ5gVdKoIh2ZT/3bddY7mQ7Ypo
5xnh65MLB6XGmtn2hxpYtsyV1DkOtit8SDcIQOOMz5UFM7hNqc+XEFdvovADLciTXhZIDucinYge
tKPB0X83bxFmPg/Cfj0+c/UOAKa3ll84GBBC7gpsOh0k+rbMhjAEaIFJ2TlVna9XJkhCI3htnpF3
sb9XbiB0pH0DXpM3xzat84z18ijB6PapEyhCEcsxNUOPNtej7ec8NwS57LEmYnnyRwKmuxgZangk
uc84bu4MENOapI0IT3Q3nVCwFcPxW7tmpMO7vwHLwYzUAh9BOnZZVXeW76b0nAFtPIMJU+2w+MiL
RvKTBw5ZGMbejvWXZ2Q3hrop0MqHtSFqh0JiHAlI1vUNV3GeNVUm9dSvGzoK6WtqKdhGK+CmRIZS
E6eqjHaV34aLO4+aFaFaHHhxyaNzHz7nx3Gqdcb9TZDcK4VAU+y5uS5wn/lhVZDZpJ3CNYZE1n5s
jrk9nmZROcsqfFJRutvQ4wkukxIdijHsAaTpZSoMjbk64cKCamqPjZWlvNRzs2NvFcShYhl8vvnB
gDdd6NDRfFozsK4VAY5bIUmBHSI5aS5g00UAiVkzAh7eO67OB/sGP2H6Mi4D2/UZBYEmBwcW6da6
8R9bkpXz8YhkNSSiCrvroStR+8zBGotu8Ys5RgPNwejUXomGZL1cqYvPcVCsOY5W+goNtVtlPxMe
GRfIGUZZfNA+l86n4xVP244toVPp2i1N6fhRU+UktVH/R7EEP9cRaVApQE+VctZnkdQvYdovMArq
DQvxOA5G7y372qn0kUkRNx5ll6Pd0zT+99OrlbG4/bQ1ELZY8u7F5edYmAK8l/HqB+tilgc1nGVF
NdXGcu+Z4ZJ4AOF00fGuZ/EIIyLfsCnLRK8EA07wPvyEHIlu2oaPw9RRsKNM0TncbB6KeWhi1VIx
iU50XVXDHpMsROO7IPHUNQUVtad+XDmrG1nmmyzG01sGh5+QTG1j7zku7IyAawmrbvjVpRCguXPI
UaaK9E09KfN/o7J8nYAneznzc22yddGR38VQw6TKUtf3kSPvhP9AP3+yZhlcgDdG7lNAEka7bnH6
kyyFPftGsXmFye1Cxj4ZHP+jlrVqjC8hy5eKz9fI8217F+OXN6kszX2x0b3zFVE1e1t3F4NC4CEy
83KEA3MOL6CY5YWbJ/p5AJfdtPKNFEOpNalG8vUr/0xh2I3yW2J+fQI1IjcEiBkpPYVjJHRh74qJ
/i2Dq0TdGmwlRcCA6a+MrWjRbwB4oOMrAu4j7dxd5v6SgR+f+AEv16tfi/jV9qVF/A9bm0X5HhYc
UYIOMYY0Vla2vI1LuxCbmgUpRkj87Yo2pmSkUICduz3A2lwekxEHxyu8kzbc1fjJ9tigJChF2Hcr
rsb9wA2k19KHZsJwqiId4EcGePAj4LnZjTc9U5UQUDL95GaYuWs5QUmjFfZqMKzMywqo4Oe80H9y
GzvPXY02KF+AhLvPjj1FzJquBnG6AGCOnCK0Xvd5c5RUlYvM60utNgfwxgADx5of3i/u/VVq9+YB
IroPLd5DeGsqLr9s3oIv3uOwW5PXAf19cOzntZ5fFgWl9QsG0OzdxZZ+d1cmAm4k0kAzYDdAHQzC
b5L5c/zz0H6MzG57nS7J7G3lPRTZKJRI9aMyvh+MEVy6rpdHlu/btsESO0CPBG32ikPdPtc6Zxwh
fEi6eB/r819O9MJ2Dm/FwycORZSBr9wTP+uN+m93UGR6NfviOw3HWW4C7jNLBy8c1rH52bn314j6
mXzA7hdkn96EEC2n+JWzQQ5nBBJ5arW3DApjXa1zW68ZmEUtW0CLSPkkRjR4/MO9szDRDDvcRGZ6
euAY9ZgRpR6C4qb2rPLn5GBl0m3ZUJFHspyPn/g4GYW4d+cMpf+j/5hXjnzRnWQ6MiYgXzmHrvff
0hKOw7DC5fg8Mxen5A3wfsuoxUzTpgJva/3Bf0JOjWlKbQgqc0hUOUloZcuSZQiPJfTReUKtfR4h
ClPUXkjCGoSrrf/oRrH8ZQh/fE/guvGFVJmyoLyb6kL1lu15d2OMXtN/D3qDnCL48WcC112Gf25J
ef3+YRZXGimcwWTGA3SLyXdSx7wQebqaehyhWiJOVqereUzUcfhGwrdPrrkOrI5RHewOgU2eUKen
Yxc1A/HYz5Rz0HDXb8MWAj0Seabz2x/Z7FEpYt3M9TARHBcPD5sKcBbHiADlKAwnMZ2cxIvdiGE6
SkdZ9nrdcFCJRqUoTDRJZgGxkqBwVBtobIPZJKzWbkMf7uGm6vR9EZuAkMNEJtZYnM+LyHCzWp6G
BLHb34sR42MQum4QS7L2QSptCnlnszWFpJl3B5VTfgA5mm7yUzvIc2mY6aCBtKGKTYNwhpFELZJQ
IDVuemxy9WziVfo6vmwdRcDurmenIYU4l8Jq6wJnHIZVEoJskj3M5eu6FuBmj+8V7P9MjkU1A8Xp
b2of75qE/c/jj21xjxzt99p5MzNOv1s3Yy/R1psi10fCv7hBBBB3IOq/SE8lZqdEV+Xjm3VqJ6p6
WPwYtj/8y3rpSO+/0KwSgjIvoeQsNSouWmhXFG6di0YPaEOURKItnM35gSXwDp78X6hsRuIrmAuY
nce9unmm0aBIbMIhaUiCL/GXAaY4LpDmZ6Ea4tgVmqNNbICUoVInqC9nxoWLwHl7MhgOfHj6W6mF
D6+0+S3Y3+LvLkHYLXJqaboGmSW0oSafXyBxDtqw0ZFe3BovEo//b/BIojrMDSefdFAQDyV1LR8b
SKvcoQYmgRSL2eZF4j9jiidrtSjkai7bgYTYUR/Hp77MrgnONdTfXABFRysezxRUEv1o6/+2N7jg
wy65mJnPJFpDj9a10UuONxYQr9aNaiT5ZQXl40qBsLTIQPk96fL8R8WakqYeqyvLp5rlbxQF+8xE
Q+uYZYarkbD1nFg6ld+uOyO+ugNcMMXyv5/6B8QOzesSrUJGErxRpw5KinEiQWHhvEs7h+1mHhrF
WSoH9IHPOhwn+9RuPFlMmZKwwVm0fbUgwsYO6plUYm4NpIK0zELrEcJ3nSdsona3SbyiJ2XFp0qq
G/w/RuF34V9OtuoA75FaJiQhZs6DIc567+NWaB30sLxAQfe4ndk7pdTXm/X2ZRlqzeCiNv6MnsNm
Sjm2ZunSr0BKvzpq5LPjTQgOeJTE3TEdu7uBwBe+wW+Tv/TTNhpqnoI9SoHdGzrzVW81zRshtN7f
pcCITgv1XA7i2DZcDl5rEk5gMwyyr7TdIqhKF7YFPh1GUdOHvJ8xImQay0WpN3ps4DsJ+HPYfNYQ
eSi3areaTAKpQS5gjQR6/eYat+OCQPWPhGlel+3LVnyLXijrsAY+iSlGhojPjUGOjzmsznuyutOv
lclufCJ3C8Hb9wSCy2NlY5iYzFy9Pk7hAwhN1XQnawfilRe/RS1HbIgoJTRjpEQJ71sGlcgFJhXF
YTSWuWCdvbOqHyLG4hOiuZbPexmVMX02BcfQFHXO5lAlI59u6amIU/277kodWzkv48q275gAG2Kj
zQvtcollGU31ssU7SPmKw2CA9WYmziQiEynQiQVdJAFjmecWNfuI8I4mAs+d3t9eJdpF8hEjh/Bv
PuDIjSr8Ca84NlMv6ZchPPkeLDdnJbef9Ziu4Mp2qeccwNjqHJKUxLf7SqKCgvR3V7ZC78wpwCw8
kgvLwAuiZagQ5MbXbSWGLHkssYDXOPHYqruwCsnxLQC7SSHywR6UBiQIHyevy2wU6aI+S/VpIF+9
lYbJgOOhDTen5xXznsZEj72ZduFRyfv5r9b1YyewY+aWfadnq/P9D6pO+gT7Ld+as40fQ0R5LCWv
8Fr3g6f3C1aqrUg73U8vB5u633Vrc4hJqnBbQ5lhxbDQGFa3cThTV+NmCKl8S1Z3Z4kwNaX+tOSS
/HwFVk30LPn2hI+kMT307Zd2qClHrjZIce82m+71LAtUZBLkFpT6LjYJ9Zm3V96RQ8AkxS6rz0ho
PMNgO7ZHkRdgefug1YDcIsAAVDIkaNZJOK5xM+9iruudQK/1XARWM/nVjYV65oK3MphBh99F9JPN
+WrtigKr019tiXL0a3cSegW7IU5M6guqjImL5Wyk7pkNGdHCZQOg7oha2VNSCyd0PtCJSgYEakoq
P4ej8qNdwWMoh8Qa+4l0RRbG+DEmScMCWNbSBlF/n/L0W97L7b48KyHstOZTYNuwO7NYdx8AtbKH
X7PL8FBeIvKUzjmX3cogs2EhbjZstsDpbY+23iUyXIdiEI4JZwxbIdpNjIu1YaxYyVfoBlAljTVi
lkXri0pumdk/t8bBVIe8ZGPxiQNuPWRHzDV1h14lwVsSF2rzM78Y5NW3XZuCVTbwU/mmByEAs2bs
lcj8s8aEzKvkzZ2139Zzg/kGo0SdGFmpzPJj+vkO9u+2zveg3Yo19uweVsnraHwnSvN+S5oStZL4
7W/CGLyqIKAeAJC2GtIUpyF+qaSzq0c9jIduCB6MYONdb0Wv/XGkQK3bObK28JUxMcqgR25n0RTa
LppwztVbFs7bC2najrzMcLSK+flpZ2blZ9xlAuVr73GVs6MAmea73p5EyE+yXcQgCZdxoNS1xHk5
TImcWNJVGVGJlspWBuZbbTUQ+mwgBAGuuO1vtD3XxgIxMGoJaj6jCBieSPVYL2lK+sAz5EITL+dB
TKKLxPuCnOEiQEsXqUekhqalmq+sWFPdUXI5NOc5j2FzLfRclbhC4OWRXQ44Rtt9E+hiD60MI1Po
OJjP+30zG8CIHjVD0viibb0BO45YIo76vNvf5OG1cVXwUeJIXZTM3tqijlQsVhu/3zlPGVFSDCKC
5lm6mak1K6C47UX9txp/QfCuaKoBHixgFBX/ewBm2bgil1SpCz5SxDM7bb0BJw1I3pIBaceZILNJ
vzP5jYky9VJ065YUMdC2pAdGN7hHNd0wMJikVBYSWW/iQ5QiUVuGF5XxEL93o2w625gPx99W8aKa
rM9lVYIutd4UWSzexE9PDfOsLOEBmYglAbzYDFrRaGlNQ+IHIHdMuQcgZJRSBjWIe7uJza/x2ZKB
Fr9VWIKI/C+42IrfEoqttravbAMZ7cmk2ebTYgmdq1bbKI9y6RptXv0r5GuLRS0A5ZKg6CRGytEP
Uz2BjxTPle+EUA6Y8dM1pdfcGMU4aHmJXyblBlL8I3pgOM1qK1oRBRZysA0to5A7MRsbenWcSTQq
NFOGu7j0F8xjJW3veHUwD5XmgWwUJ8VsjgPxeET+Bn9b9IgZDZTiJwFlgZz9vzv9QCaxtgxm+M0I
h0C02+c+jhdINO3lzeHf3T7+wGesguIznlaQYI/coNkPHGfNfdXl4IILpZV7Wy/bgfcGyLoUy9S2
GZWxDgUqmdEaW7Cz1UcwFwx0nBe+KfzcmmV6tvB16ehgVxa/TnyjG8JJ2WPZBqCKwZr1k12Vlu50
295SyE7RAGWAYU+tiU1GUKDnXNCBaVDGkgM0SHKYoSTM2pAhg5mgx72GxOjv5ql1N+5m9e341c5D
Nckcb/Vru1HR1EDyq3wYpP4VtIZIohnulDbkGz/z9p7kaJ6uIjy4FP5M8UWc/GgnkmsXRqfU8dw7
/ThdEGo7c6M8UWHdPUagirzic5TZHzDb71jNn40j2wDyXzperOmU+FZz69PUue01zz7qHiPHw8Zu
4u500+21UGzb2fHgBzTKRR1I2sbxcWokRX8ZCanYTe8Azrl36buTwLfGHx2Vg/Fz9gHtajBIm1Gw
NlHVzRj9iTR/CoMb5C4roLoaqN0iVQeWk3rwTYJRos6tnzvUO4CA00/vJTWo1a9s02kA07/aEKKB
+krCjWJMlaafAw8m5uwrFIC8feL7+ldGaMCRR4KZwHAPvYHY/vbwmJXPYJSh8LzCDueX60UtQyQV
2KePhu1EzogIFXTflK/DKjZrijx2fRapN5m6Q5mOT3AyPsiRFSdga7XYtVbWN2asWFl60Vqx5qW/
XMeo7sD134TXQTdHFZLhz6v/j1NK2uy37PRkgXbhSEZef4f4mzPKqvt8yTQ0VIFtdPqwQgIbgz+o
dH8+ZuR+wF4cFy63F+FXElPPD8XPzW603Ui67idQacxx0ffzpIk/u0BDgKtlUKWqzqt7VAUPVLEn
hZ8YJfGCb13LGS2Ps1UBiZcrWaWHjGjR2/NYitaV8HN8XJIz8HTlqOOLjWIbyTeaRIs85e0e1Py7
r+TmgCnoUjMf0RoTfoiTfPbPilYZ6Kzcrg6F4OcenLMqwSI6yF1f3I3mpVNWqhXZ1S0Z+nM8v/kL
7GC65Jn+WOtJND3tx5oj/4RVvUR+fRrB5A8xuUK8UByWdRuf9Mc2cAv/G28+ucZbcrIpAV5M0824
v/ncZdnL7v6PuVv+5fL/x1K3OFf+BXR0e5ywKLmiX7/o/HsoPzIDZM/kcBgF7v0T+dCp3DxTx8kL
S+SXWHzTFxHJ8zXmRLQbEJL+hIqEO0NrsTQtE+F+SKNmyaNXpBNnVmgEyYi4aRATKnVLfuR6mnIw
6D1Veo/dNCVQkHVBKVtz/37B6p/iVqc8uoTgFFj0flQOgP6oFSPEv2Gd4epDX+Aj9oiZTSvqwfzG
VEykPZdI4GV69FaU9ie5mGt3ppwt/RUWBnRHhDwZOM8FKAh9XTQ45Q8vdxlZIIn5C3Vsh9ZtXYsL
cxiZdXRuLYfj+3IX83WuXM72U+h9ZZmb2IVxYCB1ZioersfqMvb3bpYCMjEjuURtbcRwJH4zTC34
u5IOFIsyE9d5PTjlWFWXXkmm4tIO2YAr8QZmAui9ubLXUYwp87tUMl6agIMedH2n09ZLDuVlN+OQ
XMgR4AI+K8X2ukBwJbQWSnoFwfr8Ujchl42nn9YukANskkVHPjrd+ze1yKxS3Bjo0ratl4ysoTHr
shpq11DDfe6hxJgwUsnH0NEarpGFFh27xuVWo0tFhflVnwf/3xJwL35J9AtOH+g1hUmxiWS3TtX1
VpB9uuhfph2rGWewIaI3QSCHBTVmYOeekvM0yqBH+L/ifXo2T3ObqhzdB483OTkmHliLxlgauKcy
8YiwjMfbtU+DOVVJhI63orxJjiyaPH0PWn342tWr8ZCb5FIirIsJdO6P1ecnUmOahgLmBF8oIvft
rWWQAdHlcXbdP1iIobk0qe2kRtcP1xiFw8mi/TPQz0ZW1K/OQrrTSuH7B1x9MULFh8RM/SFDD4x/
RAMEabKX9/ba34B4wiwbVlaLvQZyywQ4/epx43YxekEOOGs/kxhK67ACxHzE4V2v22nCWjHM9zut
4uoLWX5OhYZcU/dvHblljspi2CKfRNi5NqjodiWwrgcFyK+k1WY+aDM83aRayUU4JP4SR1hYRdDD
wYiMR5d4+5fkEfQt5gknsLi8eZ+1mhcoIpvUIaXyOCj/pg6P1Lq1e4OLIAMxP6UIaA9SBAZD9XVg
mtdefSWKoMq4PUwAzwXrPSgeGVefTNopMy6JjAdMmbb0wgC++t0RQGCr72Ztlq8DHRW9Ej1SlBbQ
XBMyDOonukdlcPpCZB8oY1HzJNgxjk4JvXK2JaU+FJ0DVQScxgOi9ljTzgRieCvCZ5GN01C3wZZp
178NFcVBzFxv5fG1l1CGpxhx3p1sp+/cVB7F6JHew4tiSFNYXorbOA0EMvd2oE69gTFnWiUdOJqJ
Vf5k4SQ+SqHoT1nM0doT0CXtBKzm/U/8HaMQpTMvmp8CWUJkJtXtk92I021nCfgsRfFTbqILPuth
7/uERPgEAwywHyfYoMTAybLtVhFRKZNavdUwm49Wi/3avy8sQNm4+53mpQDhlMKCASQ0Jodp9tG8
V6z+hzFG+rW3M2Ctj694XWoHzBBYc0ZQFl4xvu3YbIpwH1N5H1dpn6RwBuM+zgc0XhH/V2mYqXU9
YhsxYUsxZFu+gbUqXfvD21LOHbKWVM2MzJ0UeIgokw+WmdyYHaajJGvhRrAP1hPM9RprzTvOLJuK
+UM1gkmuKXtgbXqQ/7mBX8O2airppkrYf9dQ2hjZMWpbXgKx7EZsmM+FdvNLEDYIuFjEkh2HodGn
DrL2Q/uNsUXBBDTHWZukW6Ic5+W4KFjf2xEI9SdGcRuban4iOMJ/fcjFM+llnu6wyytIPhZTJt1H
9QCZztr93xqbVyGNPjyhdMjb5Qe1M+2BWgCvJHbFn2QYEMl/dMf3Pz9mJebYH6+k7PNsB2Y8V+h5
KuFGeYDf+/Ina/VBDXPqOVA3nyrG+Dc3s4kWlMOnFSG11n3LmKZUnMF5bz4m4Lo3zrnWl2DfwFDu
3dO7uXqaQXA7gF96G+Yg9rTvAkiCpE1fANdjvTZZ/nc62slBesUvo41w5WO9v4r+tPL+9gpOd0XF
GQjQYNoKXwSnKmuovHPP8U22lGKqTix7aQwKvTa6KMmepr+IL05YiCMHcWYDiEOmcPCJ95mPYhxn
ibYKf8iher3W1c3h5QaVLjfyemX5edh0+V90L+YkdYE8gxoIaUKghhK5sR6w8Uo7C6Fn0GrUzJxH
KflOS0tCnd/93/1RQehNW5aesfv/nGsswC7iG71PIiRuQR3TSMVNx0f9tKojymR6fGqZTwt/aIYU
j6UrTnW3CCCwvBUSin2uUS4RuOfBXsZFZxW1kPj01C7G6IbrHuWhE5+Vsx5o27+4PVzuHqUqSyRz
PYO3HztzWsEv5ek6hJt2zplWMSiDFbBIr2BwckDM+6ZiLO6yIU3YrE1AKPNM4eB6nsJ2ADcktIMc
jE0J9tO9Zfl3Gy99iWwIJrhd37xWY5qEjJ5A8yFAPGhoW9i+rblr2uCxRsoVxVgUrajSuIFSjB3A
UiAsG9JgS2pqTa5e2g3M65AuNOO7vWlaMgRdP5NgXy4muZZV8BAMbpGcMYdnmiwQ7/KDLps77/Hy
ff9IEiHgjI6eK7X+30SHi9PMtmHRqjUvub+rgbbkC4Yp/vvC3jRAhJdYV2jgnfXTOmBXzQSwc3bd
hgOZKWNn/mZ29+GaqtlGXLmgld5k8NYt4Dbsqet4ZU4QvYfSJTc9ZmDUkF1NRTkKXc6pZadn58Ne
UyJH0rO/cMpcJI2Fy+MU3F2Fprmo3xEq5yHd1os03wTrcd4UgUK4arvfUltquKl4Fa51MjdsJ2Px
udXQJhtzlTntGFDDEEmAG8bkclFadd8XGFLmE6sbwKRJ3c0LkyCwcUR5cOmEFgP/M19sU1y4Apb6
h3+LIBpZgyysRtmPPSPAVlvV1B2wxLko6+8BFNngdq3DGYbGiBhGB1uUbYjFiu3/EYywM4JCaN46
+us7b0tnQ7+YUdO4ooB2vjrivKUJkYC029u+itCwWzrecKXaVHsxc08IQhuV+RoujVBiLn+sacCK
2tfqWn4LGhv+LYJnA76ZEVianLGyd5AuSbE87hIO3pBp0MeWUPtucRuDF3/Q+RcKEcjTKmAdyLrg
qoeT/0/ZnVtlmI4pky5aBBPvAzUab5wxf77vWnMa07QEyBfsASZ0F/Dx9yhS/srQhzMPU7jsl9wN
n/tqCdR6vh/ICTPaEUfiIZm6h9A1qJqDex/ShVyZv/KVNcSWXsVson1CHy4yufC4FvvfFXJQtpzu
4POlk14tDH3CGbeeCjK8mS8wDzyq4ZuzCUy65jfN8RGMObwX9j/ZW27DsLdOuwHKm6jwF7VumnUz
Q5mpt6jxdM2nK8qOd1m1fLkpHpgYg7QryQy3cRcNjW1ndfBm84bdO25UMyvbcW05uddu0KFwch1/
+rXFR8vrMF4JQPmn7Jg8/nvtkUMkEU24GAFg03h3ZYE74L1EaIqy8EMvAmW5X2K+kxjkRVID7mA7
Xbm3J1W7VNMaj7BDjJs+m8Zf4e1gfsFl33w/o/OGb/anZw5aRCG0Flfae4TzF2Bjmjx5C/hlCFlS
mjd2yo2CIAgJR6qKEXz8tn/axL7WVOji39lOc2OgGpRiC7S57kI/RlG+JLR4hbWppBqIg6zyROlk
7S6Hko62zNT/mMZ41Ld48bXmYOFdRIUp4c7a1evsPiiWREYKWIh8XL3oNCQ+QICXl3//8jxi4Shv
9v6R1HPxndau3zGQqH+uUBHjsoGuH97bnZ/k+GxDnqdPlcFAdoWknAVOcpAqKDjBelgIVBPJFFZe
ZH0Sv+dK2GIZmX4NAq5MjnhDjfGilIPm870evHarxexGVuHswQdFJPHbk8DcJKuemkEf6jqRa1x0
qTxh7AtnI7bO+42xY+q4Ktijg/siNUMpuqpIZkoHUZPOpNIXFj4VhHjpnIsmX9TRcR+Wt2SexbCa
XQ28wPd2xswS4R3k9YVRjJR57EEVX1cAViKpRN2uH6WJItS+8Jkl1Mmmqnn9SgCRxiKLXPzWdlzD
EjFGaYuLr94E+TJibDXFTfLWNGU55VUUQvereuol7ZQkvC+trSzg/w6Tx2/TH4/BULv139474qnn
V3fFQnMReuZ1uxvpmZ0/bLWAAi2XH1TzsS/mUG9ns0waqM9K2Fg89w/HpFFZPeu/AQ+QAYLvPrzT
OCcc7Omb1hqsVnPtRSi4boMvQnRr/uEZZHq/g5Subwv0etVYnUG3B7aanV7sf5b5y+mey6iopUy/
ngaTVCvXxwH3Mizj2tai9R1ExAybDCZ3cuLBzcno0DqTRRlPPXQFs8mT1/CX4/92VmX7wfSUVRJe
f8ddKrVndC7nLKJf+DUl7hTOFvSL1DCq3VRJ1L/PoKsD1aJ1QUfLTb+WTCbwL7uuNn+fsmeRqgBT
t/IH8KGsu1PVmCSVsgxLBdeO5iERYEz0xy/85zV91eA/CySzThQZ88EB2FzKlmegG95rdPhB1GpF
bb6Mp63BFeguW32z4w/7794mxEK67qOk6zmcYJSCIbeAIA3zyrhyYQvSZEmK7Y5WHFvwQUo8UshT
x++T0u2m8JGQGuLZHo9UA9tT9nJpjWgysSzrnTZlxVlej5ciOSpL5SxTGhVdivB+m1BsLFiAhK8z
FLxh0TKfridr3eccGL2JIXg8opYAfJfr5FQWIxluvB/O1CLtp76LI5I1YgSCEU/SGdbJYzWpCYjK
OD64XylzmXh4Am4NoVA6qetxTkWZ4ccJPQMYDYvEapDXyhDiB5EO+XDHU0C8/wQeTRrj4Ar+cD/G
fWV/tn+NscBusgQcGbR4vQyQkEmE82v23HjS4c2pfdGXVZuSfsp5FO8AvB2CY7kCP5av/RXbFdzx
SH4vX2pcAhoJZ/mHCIYfFf8eoyJ/Ty4Fir0YGScEMg7HcTJtxI7Snbc9u0YjUJ/qj72/yE0T+3K3
yvKjl2T/TlBvXnglkuxVw72fNNbwYwnAduMbPVU1ywgCS6aBF2MkNKRgqArjhnCqRTlDjOhyewcA
pMP4KMNlg/anFk0tSXbbp+GEJGQ6PQaxzymqZIGSowprNvLB9zsrv6C3FCr/WS9Gthi33WPMEHxt
rjYnr8KVJzMdMfN6rmg0nU1pEqDahI+gF7vWyermBeKJhmGsYqGAGze84NCa6lfRG8yFLH7EquYh
vyatsNBWqd7R5WK8XcbTG3Kmggtp6udJVr4FtSghGvOdHWigftjoeZcPnaZAOiHg9bCSd1mbzgt9
Re19Yay7rvzdZZT5r8Uthtg2s4QO9PQ5dKcaFKpwdqoTIS4hs+7eCSInJ7cyhJiiWDZdNsA+IIJR
v2zzDfAtSv1xsGDlBTIM0Jw6DW7YOT9IvzJi0f2H5zfoWWFshwMBbTUFRUwFzy5HtJX7tdEeVPpZ
9nnfwnS0OTB8Z3QpdDLVhR7RWv7Trfp8i0rzQDwiq46ZvvO4dAmVF6MPX8ee3uotdOQE0kybg2Kt
xzfD8cXhmTuCzwUjgWbgJUIm6osXAcabQ5jqPIbKx4Itnlq96VukCiilaidI61iF+e2+cZ2lQLrH
KeFQ0bvcu9MXw3Y/adLan+TdU8YhbvQ4ki9bC65U3Q0a201lxAyCkw32xbUEGx1Z+eTOCRBrZebC
cwI5paTwnjRCb1cJQ5uo5uo7hqtCokSNDTabZOtY1HxlUb5gkMCDgMRPAUBSEYw1gfwbAMLexJHo
O5Mwt1rj9STKwSpbTTcTlevqjykRpocALjywk0zHJU5hHH7L996ZvmDjfC5W3cBRmuXe7/o1XLUB
wIJEUACecE4WxOxPtkaNlonyUnHRDj4CED2VEtNr9Pq4WFH6cj5nqUKR7zAx0hSN8uq182Z/G9RN
6nzUAOIQb+BHTkhEyUmOAMltKzW5p5ny27mHgELzeWiOekOXkts7vY3gIMV+Lf1BE4KcrJIj1qU7
7F/YTtQ8ZnNUDhYZUj8/iuUA9PLdMClObSxCngUq7uljxPJkQdtCmVtotXsotfTWft+PuspBhXyu
w6veTT14IU+tvqd/ticPvlweio6ktQxsaOzNtfpiIOO0BXEacdcSQVJkab4apyyjlPf95cKYOJXm
v8+EU+onzOj/X5TeECHYPk1hZPVkcZnCPYYyhASSDU+RApC0Xkj+ULSBXS17lDva1mP8JTwTLNvW
himrdQQ0jpSCecjUvptH0fw9frtCnwPeDhwUImx/UTbMCMGL7V/aguxFk0cXPIKCFJS+Ms3mSr4A
JPrervacPBQSFnoIBPe63Sr3SW6XIFKQlMknD28QGFrjQ5b4vbZmulwNGWbDDgXJvggNAry1L3qP
+wmErv55n6fafAsdjQ3/HAfrqPXh77EAO6e/+WJDAgv8E3GJUrjcgByYOnTlG52x/97XlxHz+4ud
bMw4XFYAw18H6F46pQea0sMMFjvuABCWDXxb7ez6v7rJ0AMYcqX7AHsmSzRPwgDc1PbfzdfGiML1
xT7mYXDHJGQYCCLKAm7E4tJoLU2NBRQVCy9FwpbNsh8TzCHLD8jegjZkwT0u7pWEGZJFoJUVORXw
uskJUfOgfvvREzZryua7ndqPkZ5YR17LU46OhBVA5ntC3wRUMlscsiw67S9T5CyH5+OaPkdT8WvN
5/i3WUDP9Oat2l2YyaAWDD3nclKHGZyMkqwdCwCqP+2pNJpd6Al/QUzLJXvU9n0A/IyC9a5ypWbV
3QYogS0QENe4OzqlJNRKAToyHu9eaOllXDvV0+tGEd9OPbIL0bxBu3C7NzBzx3pxFKVxa70pWIoR
gOunIc0MSOaQGgd5dRNi6dDj3tO/Gubprn8fjN2IUlXhKfVb8rnNY/pO4z4V60lMy/65LGyJR2k3
NXwiVFDF9pPP5oagafb4QonBkHKGfT4xPYCfwYexM0ADdvFF69qcuxDHgTP4EC4fVTLcZf1uM5yM
YjKAw5adzDeF+ehky51IUa8jnoEbnGZQqGz05LFu1tG0AQvRycPr+scw4/uDn8NfPpgtbmk6TK14
aRFrdY3fSD7kzum9Oc7zkpt5ul6ELZgF5mHGJbo6Jqs5bb6Q/QOVnI/jiBRKenIsLlOY6chhZhWH
a5WQZxD+3Z64wUrbdKaiWtuAig4ubUQneDQJ29H5wjxkWoqQtSDw0djLTss6Vrm/16A59j1zx13b
zb1fdAERx4urgxZbxUZIN4AaOffvlO4mKkhNY9YbQxgxobB/4ir6e9D7WYAo6B97Wbj2Dxbh9RzN
3aA4zxqrhjyu2FCcDL5J4cReaEpksGq1QF6CoAJlm4bou8ufwkoTYBL+RF0FHikphJwRR7pFZKEQ
qeN7/1nwgqF7Lk4utT4NM9kQouEVQKxefoykPv9ZBhKQvZBJANwtxYJdSwgmSoggQwgQjGngpC57
GQrY748cNOyEsVom9RYwNGCcawA0oAASG3Dr09agWPIha3intvHmN49N0gDY9WoJjiCS9X+p0Fso
NbAmJeHIP6Ua/X60VAT0EcwmEo+iHMQu1JxTPF9BCnUfKaGEzUE0Au0NXtbN4Fh04oAU1ta8cpgV
WsvzfbxTn/TvGS0cRjEtBEcb5MUWbn0OBfx8/maXFHIYqLAloOJ/2k880I2tmWwq9HhKrMz1CFHR
Ye3dOycQCFjWXeHKA4agGKTssmoL8t1BwUqUad28yF/tm9nG4/9J44PYDwGWC9yYt/ozW7bdbDs9
bkfExfoHxg7XoqzSEMu3qg3E6+nmg+UdA+cxdlX3yrf9W12XB4EtLRT/HIe4NvO+MRBv7dlJFZWG
IDTKZNW9ukwbR6dJ1rnZsA7o3YYQ6HtRliUeNlO/E3wLWLe6d1ke1ezCJDW+RYVCKeRWS/u2z5ge
n6WStXHpol5ngANzzQsYxIMf3t/ALeHmFNeKpH+w1UKLXN2HcS6ogpNBCN8SCbQVNo5D2qXMeN6C
Qt4DbIbsjdmBsXjNGkCkRWS/c5iVY2/mIneXyRxMLZ6VdX7WmGEQKIQ50FquMxaSZ0OnkdEd/2QT
a7DALA8rZjlbCuM5qkY9O8ksTvcvinaq0GdeKLsZf33bIcL24lgmB2KpfUeZCMw7P97EkSt1A0Nu
7aWQ1B6LJqItiQ4Bp1LuWwJjyY+4hS5OD8W53yfzaD6AsICSlZ/WOPzp4hLcSZMizm24tpT/Aqma
DpL5nSXLvaETPHntnSjidvsrVnVP2b3yNt1dPp+W/MAr7UkcWKoIVm9tEG5AiGK5zQ4+AIQ65dkD
C+cyFd0ZAXuXthonCzgqITxBp9sth8V4aUepLM5tC/2qu4B5JhbiBC/bpgA2erPASuZ+1rwnqEjA
3ypsvwNVZaQ7fVuKquktcUG+aOdqBb6WNypd2x6Vbqw+cZ9HjdEPBu0lOqbu0mgTFuuJ6i/x4E/F
SfPq1WeVA1nVi1/rh82DJDkgpKGxYm95ZeslGokzg2oBwO0/lhRcFynqnuXSsxlBxgfQ/88wsFBG
DpskveaGXpm4yEBsQl5WThkwLN6Bl+9EcgESpuegoIhyLu/Y1bFMvQrkvu722/KbjJjNH5Yvptg7
LiqDP8UPANuH1+/miMP3MbvzxSedVOqbhHTGC3luYlAbCW10PuHirYSVbn3WeddRm4TZQQY77raG
RajWY5CQb9TWPois2ZWslZVyGchqC1QyzzsPIcMfC6S2Bffi2GPgJZNEHLZYUoV5joBXscy5naw7
vWKWYi2t2Yqu+nOwD6UWYF8tJQ+Fr9+oY2VCOgYLUEniJa6Vzm2NDaGr5f8cWBS6qGOBuu202DdJ
TV8Ecn1SN2oHNS7Koi8+MSNiuQOpIlxa8Rm/hFWS7k3N61i3f2mjav51KOifZQCAYnwCo14P0MOv
FhVk36SbU1EDvCO4rgCB0SFPNngogJyiQKb68zAo0Noa6drPg3zdAijSpp6D+AML0Cf+jDhhruDR
Zj9Z/BO7HsNg9R7WY0VjD1kczZwN4d4IDItOl/zTehxbyjcDIPL09hTsJ5IOusDRcK2wvbXxNcSW
wMP+C8q0AIz6w1NwuSCNqJgyq3AxOHIP0g8aEe8yotUulOAnmCNpOEhX8N+oGfSHrkJCoTh2hrnt
VEJZ5tRrW4nAsfo3udXFEaEtoLz2SViWapj4iGpb6RgunM++cYGvT1clXZXGJk5W+OEh/SiSnP7E
feZ5MkjkLGcII1miUZXF3fGEzP8zV7eI8bap5JtrprnPR3H8BA1+W8p2PVcUL87w4PVKmRAq+7cm
dl5MTmJsWdowMIlOXVQD602FyWfLjVGIp5H6wvb5hwRTMhS/Z905aBzmB9F7HXEKZwN9lGkQTb1o
fc02dU2O2OYtAK/lGUxgE3ZL9n3oSE0S8Tm0QHfCzYPAV2WLnZ8XfYEC/56Hhe84k1uA1EzITVmh
TzBPNrTMVABtReAgX7Bs4LuNgHG/TZ9lvKVGXxRFZfw9MwUTpnOXVcArWqxw9NZqPptlbUsETh8z
dsFBLQWX7afkTysMjGah4QhlZxRbkSRfC9SJPa94ofCq1eQlS4gl2oKIGeW2p251UE4gsaAAX0Dm
0lPD1yZVYfNnVOsghyolPDYsETUpwJqboVo90DYLL0FZ3/SI5oW4TZhvs9vZjREunCDDfNjcwTOK
rCBmw6BFhPLrST/amBdSRtiPPLbv+AxeEiwXYGVmpLGysinOU374PODvnqM2nnE7jbhzNiDyhg0L
15i+yIhpbEU/TpR/RiY2XFBBpzTjsca1V4pn2pFFTv/eE/FZhOQZRfPyJGINb6sf9wHVNUyCWOo0
bSugYK3dD18S2GdNIiVeEQjcBf+6PLrFIrtQ7oB6aAFZnY/MOmXJf5hcIOGrA/LUPHAb41KbSsA0
WTFE9J2ZhThTNAyZzRHWRhHMIGKRhhI8sB3BSCyeznVaf68e3yrdWu1ZNz3XFZsMp0d8gLlnHJDn
e4cYxGaVbl4UdGPfZjAGKQlEcMYySnpRbJu9GFfX5klO5LateJOA/lEXFqzeDqqmjxGFk56D1AAK
CB104TJWJbqGl+BUmltfslWx1RQD7xN/17NEqnN0OeVMz3830IHTv770VCtkWg5a95JMkGZzBuMm
jxYumEs6ZTHhUPCnv1x8GJi6B4zA4cp17FZD4kTVi1dJ0/grNJZaVeZmjM5WnlIHaYn4iBBmMaxo
S4nyREZBaddJ+3lPmQDILEJHBRfahxIDK956mc2kF99UpPln/uXhjY+mNDQ9QaWqO3u31aG+2Vmm
KkHDKC4aOIQes1cvi7bzWQDE4u655oWLJsvn8W9QfsG0iQi5fg15T5+HDhbm1hnJ2FvpJSZdkGAW
G1EQWLt8xA58NLUqZDmVDMAMc1B183vR2EsYzmszpl7vvtiupXLeXRgZ3+eYVp292zSS4H6Jk8I2
MIo2gBOutM0nvZaOxQf5pL0oRnmyLeFWhxFL+MfYX9eLra82vEi37jPhJ9U4hfpyNgkrp54wOfjM
zv3E9Qrq4G6wUM2B9awAjqKkvArEXrOivkBE2/o07iYg1TMvYxWfreUbE5RytY3SCR5DZBxxtHg3
fOY9FaVW8beBihZUdXz1KCH5YRI2JlbHJZ0yw/t1VjP4q9S4ZdJJ0ukRMTw/PfXRQdsngAXYuaYo
CKQUUJKfBQnxe3WI/1SjowrHqEHIiPqX3vgUsHenQJROk/m+utO//EoY/711kGR1MAzLOpgBEfcD
S4gTwfmz5h7egXYb9Hj7ihXVsUM03MdEr9EOWGzahCEKThLE8X2XyXLp7LGjJFHnHd3FArx8xTTx
UbbkQluqwqFFVmqMSHYc0vhbCWGKzjitFmlaErqCLgA4PeY9oCZqll+a6I691+mYAWF+cphhE5uu
SaU6swDpjpDgcsrpfDTXKpqtKiVJLp2H2Aws+W8v1OukwV15JtOSavGPi4y9B2+dOW6trbIlsMVb
qIMFt3oR4BiBdZrZXmhXkxZRx2r28CreoGGbGn/QevRxp25SjxyFc0d+nrbAsn52QP83aqZh4ho9
9bnj6Q9mmUSISPDeLHpjfMy7vXKhxpnOTxoL9Lq/mLUoda8Ly3AfjgxZQPq/mDfnphURYcvzupRf
mfqeNt/X6sCuQHHERy6qO9d9+5rVPQqWBhfaYL99pzNQYalPC6KMF/K0uC32qSVE7MdWWJ012Q7G
31Y01qIkxYgH7eBDYlNRiTgytwRrv76j1/g5+5xcSN4d0qUqeiAKgb1PWhX+9sNnN/WTs6A03XBq
Y6ppjPBfDDxNWXwJ5iUG3cqevNGSA82sx8GJus72vD4VdD0EV1vrf3KmbMMe3FzqUcatDFjpq3TX
jmx49iOIckCRdmtEGz48+XhwBIQICaWPP47I43M5C4NZQ+E8781cHr2PEt8gANKh1oIAeGxiu+4m
gEBnRcUV0p7n4FpyCqv4A8GG/Za+S6pheX/jcbtPeLbnmSzVE5NAxdnBmtM0cAIQ/a7VeO0T5T74
o52+m2vXOk79iCEhPZOZRfJNnGbptpa/YJjC9ypzMoDmsI+xgRBm3bxsTP149QF6n6hTXzqMsH/u
hAKTW7YwUiV7BvX6//OvgYV4Tda68a32qEgXYEDSrcYNH6uBh6FNSZjkbjud1k8+bDmWu9y0DKTW
fetmk5mKCRbw9oPaazWz58gbLvwz2wVf4s4mUI8a8Yq+zKBbA1MqOGzxXfxR8PUzbY6V6QahkWit
/0HcKI+N/gdkGWxIwU2GWNwDI69btDM+YcqKrZupX1WDECtpT+3kMDPMRWe2YErP7FwtWAdkRpMj
fN8hLRlNVljFewNE80p520Gs8501DDUAaoZ5W8vWr1h9ldmfp+DlCYPvaLIv6oYPW8Efyys8hcU1
MxBKh0PmqB72DJbf6NTxbbg5GaiQat4vxhdkqM7pP1UjD/D8jQAzAhopkKnaduPgIVfm0Ipxgvnw
8YLhc9NxXwd/F6u0slO0WtWgpF8uVfgfq+oBCYkxB6WAXTvGI4J0aTdhVOBA1DHCE8B3LZEmVUPq
NlYJBPCqDCA+W1degWLYNWkQ1Ob2vUGz6WulMFvjep9xTrDzo2l1VmygLRjwbIv7S/yBd8WHS+XD
+203fg2dz+giSnRTjBhANdMM8G2T3AhvgLTacT+6mxN4GXSv4DC3ROK3CEH7z03pIZmXUxRz9eQG
qHQfO+KygZrtPQl6oTvrhdNKm3mfi++QvZfAg0pfKaEulXU+rt+1UB28SE1pv1GR3b7GQ6ILvyaf
NBkOlOCAQO9CRXHu/kNhQYGqOecb8VMsuD7g/oTfQPe/OHSTJJnhtk8NnMuImpYdD/BADq7WG4gO
9sDp4cTdI2Oz4Ra7frw3eGmKradAXTbFzEVNMvF+oqm5SEI6c+sR54VCnf2VokDD222WPNzpGY4R
9TLokrWmUpzlC/1Jx6SU2JTrAsqVNcL2G7TlfwTak/zug9p5knkpcD/YBX6cCqXl2tk7Xg6wpJ8r
hai33dqk6/s7u91hT/bRqGqvfAlwO56O1rzRcrL2a8eJVyKAM8iWfFcvMOcPWYxYv7blpBJkH+HH
p0INhMwLWhNGQ5l4CEQPc073aq1oFSHIHfy9ShWTgkx1PZLgtjpMk5wx2bS8oyg4oQMTMcybGf2W
C5SPC+GUUf+b85Hci1ZGs7PopHnEsGJNhUmcrO4XA1Vv5S5n2zz7DHCOUN/5pp4r5gjXSk5S7HOe
a02ff5OXc6HXkM3KKNTKf3nv/YqaL7Aq+EMeUK8fH1Jbi14/ASTQmQl48zq8osXZLkGKxNuNCxT+
yhkHOi7VmksmSRr7Mt4z3ZKwhYH2y5D46+6j0fiUX5iHd416XZaE8GkWLWwO7Nn9ukoK4vYa2oZ2
gXZ2lQXzbXWzci/DNMRJ310RA544/GyTLW7YtjUY+cbulbTZLSm4fTswUvs0t9avBozq17o+WwzB
OD+A7NiMMmtN2NsYetb18gjSARysFyjZlkMX+oqBiQ77YMgEsxR5OZ1r7AB7DOrdP6mLbjOUIlcF
QTR/9bMY/Sv/lgzVh4x4J+7Ay+qfoXLVaV258eQPCNtMOwG20e7f/JPzEgOn4D50kqdXQikcWIMO
hhA9Ic28eaUX90+z0jtP0rZSSidgSo0byhca3Ny6C4x/B+eRxNzmoXyElYmmnaw2QWA58KL5imAZ
QDJTYLkwzXKg+N743rq4DouoTGDTfbDo4SJEERcHlABvWwK5DMZ/+gd5ndXhk1lBPOT1wY8f18oq
TDGJuWkJx+3TDSG7TmLZmXfO3lMe96He5ZILvKdzUUWkS3dLSGy0UjVQtqDBmuRR0ZhMW9unu181
ULAU6EWFFFlLLjS3tK5CXsko7MVZBWEPj7AyWRWln0LM2O55IGLDO9EIF3bcSFSbA5ThwDwTlI1q
YsGhKzi1kzb1FWlX/NUmu0HkGdQC2uq0XwbjnUs8hCFGw6f6/RmQH3BYmjVPUZ76l55BCv8cs/to
kK7knPxmUq6WTvIEyY3SgJxbsjZ97O/37K+w5imDVVca5K0S1YFtEr5XE9yfWd6EK/VRcAk780bq
v3lmLbfyXmFSTXgsrTlWi2FlsmAmWUwFOmjg2l8wsGbdx/MJfBYYXtaP/mrO/jRhVrA1JXdGKn3I
hrVcREXVL0+wap3dCg8VirGlcUQXx6K5fNVH5J1/JzakE/GM6xUfvwMWvHn+JzE/NCrxDto524eM
dV31ukAIPC0cJzORkSwntMfTrM4cMnDhFfInI/h/SX5TlFNZ8dVOjjj5DvHVGI+/e9FexJR88sC2
kyaJ1Tsk8dUc8C29I8nfU90zMCRkvZVsUyJulH8I5v6zLPvpFq87od/EUtizqJXj6UOPvJT9GFIO
8fKNhuAiPlFvyayJBW6ep8g2jL/OmxAmER/z4ipe2sKnd1Di40JFjL2Hq66hd3NJUX+m7fDoIfbQ
Ue2OpC1a2JDS4EM7AmUbUPxeTUKHUbBdopEHPfHlYcjWKPzuZ3hsXXWwAgGE0KT9qVG25qmn8UNM
Bg3NLM4Hg6WNbxq1qhOZpiuGwE1TZXHWdkDcvxXCzjob6txvtcSBZI+vbICAk1Q4Ui6nAkmAlxkK
jXEqF/gFg5Wbu6tw/hj/fpT5+/VElEWyZJJNpGAlpAoHU4omYbjrjb12LdIbgwW4Du4/T32TuJZs
5CvzR1uKFp0z+A1dd22M3g0TzQAlfQzz/mOVi8RI3Fk2T20Jxha1lI6CrVBCUqDqktaaDSJipJ4H
lm0B2h+NgemQcjR/vYrkZrqXnM602SXaFlYyS4AvCVI8I9ImsmkzGX9LI8ul38FtNNPTjzwyJcKn
1cfV6usEvNA3se57/eyyxNzBu8MOR6/cR6EyIXbaorlaCT8k4aBSJ0MLt4Kxoz/Lci4s5rTEskf2
AazBu8j577RQ5Pi1HEJd2AA8e5v2CRKapXXDzwfYscftABbZ6Ms/1nPonClgH7/snFpIT29oOwIZ
z8wJ5nwwCJUDnzZTD5b+AG66eAgmVPIfwCwTKO+lvdYvrZRwxlJHyfXxmCHoel86qGv0GiNc3DKk
lL4DLgYpUGdK8vpWNHDjuC136diDVP9Y0WRYUmcyA2cpFG/m2AVmupsE7cs5hTMeEyfH3uT2iE3V
3qcSa/yflycVUnAld++ilYulKysdtRtIXZbY6oDcP6hWa1OHJcqaVg2mMDm4X/6Xih4QuUPYiRcq
YnI4FFoW/Mk+RkSuwttFGPisMdBZjveEpNMzH4zniVXB/snEHNO/zqZA1kTsi7bH8U5jiuNbaU1r
4Cmv+V4tJrRgpNOJLCKG/YyWAXWvQKkzuqS3o0cncTullZGOCUHEczU6ri2e+outeeYtlFO3TZFY
dCMFir/r4JXbUCrNweijdemkhpN9mJuLuEqGz/jZWUNL5mijwO0kXYf/+E6GB/KjDaMNExN2xpEj
0qWhafo2O1jHMlhYxv/eRO2eeBwgT91XS0czit277rNf5R8p4TzDXcqhaaUq9fhijjgoHAwKtLgF
+i7QbEyBSeh9Cg6OtUqK/mKnmlVX5srrs6lnsCP5fZKg13UuaFmheMIe3g2K2fm0GcghljEhoL13
rFa+/U956BPJPyN771Y+8f065x76resYO9kT6xi1txDA83dGQSAaN/XyKdsFg/IelS27gZGQxR+d
6NYwTi7zZYx2mUVhe49vDXJbvH9GQOCT7a1+TriLfTGQNAkhkQw/Lz/iDSVlmXAQXQnRHMXMjiVu
KIDuvuUXvhoCBsJZi5FjCIO8WUMnOYRM1hCPPERCPq9SceBl8mbnBCST49/AmMT1Kf+IwGE5uYVz
i6UZLjNBdRbNxPdBa9rNa0vAl+zkYpp3edOqZAOBNz71sBK2jZCbwumO7I2ZBgrVwD94/LA+NyGU
m2pfNw6gELfOSaQI8U5YlKX0uLv6u1aV49IXNdzD7a0LalWKA7ug1XNTkKqa6neZ5wnaORUXxCJi
Dk2jDHsr5t3zlenBHqYNwYdztEnIscYcp6svxHAR383Qs1gnGtcdmd4DW2Os1RU5yhRWyrngkRK9
fj9c3PNai4Y831E6Xrd5Nkr741rmYa2drUVTcFaanJt5ghM2hJm1EgivLvFizLNBZGcHaUBxSSWo
fiGmdedk+hpt8FLxnb8EJw7vNk2XBBupQ8AY+BLbX+TlPB8YmVOpV8MsVZFWs/tb3+rnwwHC3qQa
nnlFvf4+dt/UtG5cDKghIVlzQ9FCenBuCIcfYAlr+U58eKOUHVhNEoO79Iy+7jVY7mfEfZA7jxIf
zqwaAV00i93ZzOnEZM17qw8Modz9EorynwJ/mFOqY6nMETBEt9idQDe+yXqGq5ly7f9zCaFP4LQm
geaXq91icGAxpAUorhxk7MH1owL03kOz7kqwo4avyPJ9xV0dKtf76YVP9LTlTcxUrTG0AM+X0NOQ
qvIBk6pq+VoyGevnS4jTgCKFuvhS8hXbltk0iu72MRP/qvYsqvw2W9tPob36CLnN5iAS+91kS9lF
Hohg1I+/oq5i+XKEzVHDei+AC7kC+4znssD9y9As4xDn4lUg13sF7xcxNUs+w4/wf5BHSu8nF34X
9rtYtqFt5SnmT3kv5S9B1e8oYuaab4K/8c2aTgrTamfagjeW/hXm73+ZzKl8NiKgdiQcksnIC7zT
jZ+pU4HN5lX2npbGONS9p4sY0ch/Ob4ZXcNv7YRgd8ZW14K3zZ5Tv2h9xBaqFkFz3nn0RTH8XY4g
GYedsfx34H1bkniFXIrTAI0RrsXq5UYIG430k7OMp3XwFD0Xj2DlecT+yV7C6RvDGjkA5X8BCkee
W40DgOh3Jx/lCsPQDFHQigpdvNHxu5Wov/3pH54inBEv7ZLgB8AR7ExzAGXwZMgSz40BjPmYPovZ
SQXy0PncmcwZGTAOloNdl3BYyIx/UXrEg6vlxXRvZC/nKt3/O95kBe5JZ8gMbtEZYFyKRkd1aFTP
TtGh+XztMGOMrJCa9vIxJkUgyCi+i0JKc5RhJ2R/b+uttvGHG9scoVB4ksMUJAx3wEV8N9ocPm/p
EY4GBTnqPOs4aAZ8+410+shwGztL4GXzLh0eIMH+3Z1GhsRut1jq+eT4S8/53F4MaPg4YMvebTLS
1LQg83zxlWAS1RtoVYbLcJmu94b3E/jCAiPYVeI9GFFvAUqhBmYFiu3osaIPWpQ2+eE3XUWbVYI8
wnJ9GUEfjZsxdNF4dkRSqL3R+Cmi6PXbVsjs8ZnGqtN7VFZpGWgAqQj/O19YOxFqz+PuZ8Yk8c1f
aFgLJlgmP6HGREPCaOxPYVgdOdWOHCPZAuKIYsZH47s3pSgH487P1mHlBAyOW3YpL3P7Pyi5yQ8g
m9+y7MPwzrJ1pE9b1fSCk/vFakOT2JGkPFluVFgBEAkAO3EO99q+Lj+mUL88lNqPia5vyMoaDv5Q
JPyB/s8Phys4wxp4D5NIBoxtmoL2y2wfLXLdBvNtaUBW3EEPqECCUqTVDDjI2Tmyrxa12hozZkRz
SG+3seLDbMjjEGayokf78n9daCBArvwwrbn61s8/ok7o54X4AHKyfAUW797KalZewpxemUvKLPIe
pAxoyQE1FJT4kdp1ctPcV1R05S4y20kqkM80TPGz1zpGoXnJPUirSZRAzV4U82YHjSMOOm8C/x9A
7nHRm8ZRwJhEsNwW8nYBbUs8eqteNJZKWkh9S4+A7sO2HMu5TH0k0OFN92DIa9chxhJSoRQf7zoq
5B2lEA6dl0lgmV4TQFMeHMybHj7tpb+A8dSqb0AJJeeC6+WaSbOmwXMzS1vOhVj57LfLqyULwqPX
lWsd8jxlMUQwjF8AF0ZH6d1FYarbsJ3OwD8ODVHZ09O7peRi9hweIR80vm6R3jj3ECr39yiFhHSa
8vvVuJy+ZEI5HYPMBmBZDGvbG9LzEs4oLCobJLBYWCqfHxZQkmH1OlGrFqIcE5mZWjB8oNML422e
6xZKnbrbjyVRtqf1uYKn2oLIbi4q2kEOv2d55a0exoU3Sjm07y1yZQi+j3tfgAAG5It3DX+8KoVZ
bSCPCdencLuBNLf5RrkljAtvNAuYfw1FJhZcPzJVtgcdyIRClHcgBAwZ3x39pZF9WyZ5UAiCOi++
MSWz0t041fPPZrRYpKQJg+TRoHrLC/vsOGo/g0A/rdF4+D873ivX+AIH5Slobrm2Yk9c0rasJPIz
zzUFlCD0U60+OsJutK+6apQ8WEfB5SK6bHXVmlcmZPHTYkgWWed8o8kOxjilbbOlJMT3utASilaL
e4FGXmtErKR4a9Cp0vMKg2wP+9z7RGvnhTNlBQW9MacrHMd2oWy0yCJYmf3CSGQm3Tddf3iWKZzW
xpQCn3tbbU4Skm8dBR4WB8p/Lq3aZoKEsfkoR8hUcV0BMJ9sSI65JCOTKQccJwibt+27Tf+EkA50
MCY8M1e3+wgIbaf52DMSlcScOKUh4My5FAvfbzIjKjMABLXEFviJqNpu49vasWsyRXOfknVtcAff
Wh+c//+X8FfGJC5EqfvktagjF8DLfLAbtS/VfbjGE6trGK5P+85hLsyP3lANarJtazipKCW/B45g
LUroGA28eOHusnDVHM1mf+pc5+8qvGeBo3TCrijtnAH8t2zTT98PodCNhX4NOxQnXZ0xp4txk8nw
s9E4F7IVaEZ75bJ3lEEsEwHolLQKsCh8qXnigmm3BpgS2a28PJMqYDHfkhwjoNmlljEareslX5/C
JKlS3oSxi8OvsXAi9i7KxzirCZJVSFYame8xMwwYXyz8fHpShMo9sI8GX1bkENsc5sZmEkNOgn6B
1nKK+Lbjv/Z+dCWSSnKGKlttVgpHtlE4wN2d/uJCKBxDmuqGav0PAqqGmFIlq63WTCwZvc2eQjL1
Jbx3+j0BQvxiKqddJH9OVAINX0M2nYIzMoUrOWHGfGkafe037aBDsZ2oOpj12CMw197Uhu3m2QZw
zhggLsEsJrP/iNjsXaQBAO6qp8IanyQiel9kXVibZv/1qy9AjjEPe6nDZ4SPtjcNWYOm46dGhI5r
DabVZw139KN0zHl0IEw17OvMYKHJISNMjK8OonXRqRDEP9nsibFHA+1Cv1WiJjMys/GSsQ4gOOCo
ZgGRtLqlsF9FEd9rukoXnUyfdcZtbtC2OmHrOmDHf9pkiItm2hVL4tjweEpf8YnYRBweIQcGDJhU
20TpBdXU9byoY/SLca2pHzUBG3IdIk/k18yJ0cRkh3zgBB5G3INQsGNj8Ftg4OvVCmmdmrhm/SS6
u3jmDHY6W9VhgxEkIxqipKai0m3UTf+6czy/0cEZ5dEwAdfIJj2tfkM/B9WXlUwf1buIniYLQliN
e3z6O9WaeQJGbFRkyjCI3jIWANEx30lHkLdE9H9e54NsNN1JIKKGGWwrNrjHngYzMSuEUBgk0g3r
VMT2N8I2ihk9lZQIAfPVkO8MDKWIuVi1MTAvJYb9AKsiayKycta4L7otU7U1zBMxaXwPWq8/CTNZ
hWkpUlDVoVbbeNfvMn4SiPk0PitcSaytzWyKiKbIILJhN3JuxO9mgq1of8z1OJmkVJ5pPgR63VvI
gpuQNFwl0gMTCMvhNpETM8Fk9GdmB7SnYUt8bK4R67FjoAbq8Fl5GO/I33dQpKlo3wAGca/8hnNw
iI8CBco7u1rG6dYhT/nsmqYdFCAOhlHUfLy03xD9QW1N9JhsmM7xFPyarhk9Hp5EkBccDSNw6vzC
sTRmk8KPhui/OUSRldcpyjceGgVCvqZZrGKxsSBf78A8lqK69SLH6xa4WFRRWCICFdx56u4yoXie
opLNy7K/np/vit2GxzSnIiOAYZKs/Kr8EciXhyALfap3a9kVzVjuSZndAnQx9k/Y36MM+d8Q6X1q
K43/WPv51v+Lbu3HmgJ1uvf6dLmShAsbXy9xWsptWFZM1fPxGjH/DFGIThlVQJi3dvHQ22Uhw+cW
joK/LMCH/zJqfRb5bbnNCsQj1tMfwgKOrrzZUEmBF61tZQ3ykoI9igmLAKDA1T/NeNQ5CO6D1J+X
YprABznvZOHDGbkvgYzSjRmXiXMCOEz6EzsjBPSMOIc1MPzgIIwXvyRkwmImxhIsIp9qMnVRCRJq
EUhZL16IfFbllnigV0aImv4KN4eK3LdySikpqsSWjcPwLPu0wdUGfgnUHDk31FAVtiMGSn5G9heu
aO6KKXFzOeZ45FlXTtqM4bD/kD21xAYuoeK6wgkivaf2mI/PUxhyDo/hlbk5lRlAjYXHW4RDbn2M
luXty7hNJ+FRsmuoJDbxIbQSZ0v3djSnYTyUR8GOerItS9AsjpSScxFjECBiTbVzRpzC760ghhkX
YOIDFtmoY7MKn+kX09l3xg/8g8/a0C8Jqv/8aUhVnYX7EeU6KUO7AAsDDpG6XIjbZ/VPyihooWIu
k8JXs9jkP4t6bY9064rP1wOqH+3u5MMZgRJ3H3IVPsRfKxEmZFkv+CILs4OEGxD6k7nchE+M6E3w
MkM7ZPs1v2SBpxVaNEgPGOq0+M2wkMO8oOOUXl3uHgqChyw8wvSDvL0K6YGsSYnBlryFPEiFuy5Y
O+qOxV7FtdlNVEy7b1SBo6llhuyOvs+HFErsAKSS0MzZJDJpqPTh/4x+pkn1yKvLqIZqmDN/PLN4
2X/wdtPgoT3TmK7M0PqxWzNA4yv5vv+inLC0L2I4jbZaAAgZo9c3VdXAREMoqOZnJS9+xnUWNRyd
AD8A30+foiFYqzebLctOBQvxDs1ZQlGTZcI4B04FNlu04lwt+W6gCRzZLuyjpLJ/cqRCIRT+Ldbi
IF3ORduG3b90MB4bCJYhSfyCHt7G7GtxaRUF4yEPhxZnKM/73qUh10UOI9CzysYCx/3nUHFNliii
yUwNAn2x5ORvR2k9TsxpZS0470yRQgx0UBYB+fPTGnnK5PRffMTfn8XLn6tTblsned5af+uFx0Iv
G8C1ZhwX8ln1C8EdpS1hOKX5hkf2zo2DnrbYxHbeJLG91GGy+4E70BcXMoBD4cnmMEy4JeDz+cO/
Igyzs5z7NJNb95tOeNRBQ0XwTRKuqTQ6cBngZu/paPue5SIJOSXyOFt2OdZmgB4Jhs+Bf2UA1dOS
cXELkMIWiiZg/OBgHFvVGG8Ad0/uk/2eRlJgGPqZhC9cn/v7Wi7pB9jmNUg1W41KcQZaghwfDMMm
1/fyP6hmnThDKGp3Odb7UDU1vheA/divA2kClty9v9CdzyAC89GEm1iJi4hKII0pgo4qBAiz4ZWZ
NxAxB+0+qfBXRtsjPB5HollikwW34Xo+KII+/54y2ATCKQeuEHxXT/OoTuM3YDq750M3YO0s7IZE
ek6LosOtbgGFBZH5WrYBgHI2g/FRTtJ680JWeB2aawC0zun8RuE02Drvr+D4QHRw5bJLOsA58tF3
7mvyWKSBNYgxe1HvXaGOgdd27ciVWuVDrPIOMPemHwbCOx+3aG/q/Gx5DsduZ8o+tx6mLc0n4yhz
pf4Yf+7t19pkAa9p/SAFGWuwbHn6UYP4YRSy63mSbJCfgYsnx/jpMjNXD7hJ8RrUumYWlc+pAhlO
xsZ+R/qfHfE8m6ilpxM8iuDAEZARo4OdnroPEBrWFxd7Z3yysbMLpYrETEZbKecjUSdBNhqEQ9eZ
hPjI91gQ/dnVte/GIClbHugnmApsJRdCTakQ+qW3nb2bj9Y4Q/J1q7sjs3+W9E2VYx7yTCd6gK/d
V258ZDjq8W/yte+IEiM0tMP3O+v0LwocSBh5kA32cvqOfPN6UVb5A3N4WbnZcq61fkL6pDcPSjXY
NIFiont8oCN4U7iFo4y9AIJ5H2XVE5BxDdtBavzxJ5RTVVZz0DS6qQMSGSsToji6yXCBA413KO0x
bbWl63WxU/Xv2ZULa5ukfP2mbaApGGQhvofYYQ3h80g4zH6mIUlG6/7dJi87q0WWGt0jdZNSJzI0
Nx+6XYv3fwMPbDYDsrWyIERQ9tLd5i0Xs4qVAjUdOmq/bE4Eo9m9NMkvbdLISvbzOoQYvtz8kyRC
e5I9S7y2RSWLN8rKHlz4HKj/llOESD4o8McUopyTmtsaGzQLdQsN2j6zRs3NwOUEttMh13zlCUAi
hZWe207Kh7v/DlCDvcFHb35KZ0QYaQUMoCPX6g5cSK5/oCz+hncJzEMTURQJ+74HECbNw/KXdKZV
fw81Rv85AE+6JtQIh3u+IpYETbEwFRZcQTw39czyR84nFgGKXF+kzjEWNVJNMk3LCcRPnv9zj+ag
3S05zpj8aATMjpW+9yCNh5XW11V0chpQh603sqywVfotprcnKeFq6uXzLkI11QstTuH2lUnFTy39
K4MJdF1+/pOuKtxJMifFZb3TVqB+T8pdQ8NGq35dY3W9DqAq82P+CHB/po2l9R4KlI3u+UytCA6r
AYlOMr4QlkmyjaxO054N1pwV7L9mibECoQ4lLxwSO8w7WaDj9Kazk7Am4YL3f+jZiOvfzPcY0rST
WuFNgAjzzZMsPu0NiQtgWl6Ob0jg5rI219PHMl91Aev56PLlbitzyp619w1dFQK7g7WFH+vU6qw0
3DwzTI7h0bJ97f3c31ambJ6MlWIXVsHag3sXikceiygGZdEZABe2C5K2IjhilWcmLcLfXtVfncRg
0tIiZ5qPODllg0uR2AXaepxihU7v2KY2+XDpeFDvoLMHWCJ33jdq3JfU7IrAlANEiQKomwFtvYen
1IPaqfn2YPR/g5wgH3SzlsSJg7dQEKQXXplxAoeY8zKc0fDMkZE0K5ko12Clt8Xja0xvsA4egGe/
o2uL/2qoiaU7vt1bbax7zoLigJpX0hCecp4sswvDTzsCaE04Qvx6oO1TZSLIZYyiuKB0kZsZl41w
QwstrOlboO4CaVVfRaHndvTJN4uMrOOLesg2b/gXTqgLdugDslVQWatB1qc05cvS/kkCw8lXbtpl
zDsieL42UA/KNjdypeckq0xsRc1r9aww+iChFYdVKclmYE//+9PFZ2i5yw+9c9QC9bCie4zZQ5yE
+APbkZJdI/0sFSlA9wXM+Cid86odiPtB3q5qHx+Q45sdIyRshVi+0UlB0apZgUji4MoRs4KmbzqZ
qxiv9QUMpjCEj2RuLBcdKwyAG3gBPtgLZi7rlFQ9gr5Y2ZPMbPb+++++fwFyxfLP9NXE7/wwqcwK
8Wy3h+t+jD34vrWI312cjC3oDQIfUjfrCZSV2vOL+yOOOpbBpQyvnR9m70ulyDs0c+pXROQqmH6m
oJ5aW1ZwsBkTloRFKBoxV461ru6/OWRHX4YzQWsW4NcIaf7t2DoHYGJ2y+2SHr4oA2uvWoAsdWpC
z5NokaWjv6dQ0qBfcQxocb5Rz6RuD0hi6K7NdGuuK8P3trsLGrE8Z1Va8p7xkvBfSHge93cjnkYl
OY0XJMMX4kOnruMKluSTRR3cEAGTkfKz7DKmxOgaWCyY87cID0AKPNygT9ot3oAVW7SNzjlEbVXL
HyHh6qZ5DAQr4qlUS4JG/QsIsTutt2Fnkqnj84GpbpRRTWsv7FcKHEU7Zz3hzCVrK2ciNdJkR+LA
+jSEkwWgt+CwFJ7A2xY/sszJyojW0DmDWgyg1xbe4wk5XuFGJJ+yzSY4wpPhydYghK9us+k3ktsv
duyVhsI2WqdcqjxVVEzGMEavvqBCjVcJ0M2VqxE/07wfr7WK8tvC8JsngvQmMdNlYi8C8ksmriAN
b3Kj8i/C+yhr91JzASjrHuhEiBRdV4ydOczNNNDo9OTEGCMR4X0g7/5u4J3TCNZRMBlr79fLqqmg
s6pSSWVLUTklBvQ8viTtPjXrkp48h/tajcIokXakFBdfgVVXU9II27S2RZ/lTP0OdrAGKjuJTU8M
wTxeEeEHAPIrQiyWMM7j8ly2BHGUxmf4lRdMWtkJ5gLBvezc7OYKeudDAE90AKp9nksRrHtfc9Hr
r1zIJJp36rPPwCQOJrzZytBGKLEHb8E/vpLt7JxGm6eEUpIoEHsukvQgUgsq9gwn2CCZWuA18l/9
lG4zydYLVtY0NG+GnQQ6xrl7KPCTWT2nJNMjXwXfx0D6Nh5QckD3b2DBeztvPHLKHAeO1LLOrcZu
wMoqk4BuPY8vcu8bWFItfedHa3r2GDv8SJycaYpYFm9QEg0nIA2N8s/yUxi8dlXGKxLiy37GYbom
YpwYPbb+UElLHFOxfoxYHg8V6HGPTEOkmo6juvi7FDzipjfjpl3bHCOR/k1/eDfdqoCE+t7I640h
eOjX0jnMUFBSJnkOA8atHhy8TmaEG7d/zAER88wXuG+ZhEMNMXe6+QlMwv0YNgYQQzDkU1FuvDEu
c1q6fVQIU375aavvoRWQsJ/1reqaaKLV5Cs4HORGOkfdgMw/irHmZAgxxhk50wIKWUdnUby0Njxk
5SvpAWRqz2SEdgSRC5cbewEpop4PIp0r/1TIjbS6Vz7V4j0cl3QUhK6md4eqrC9voqfOladcZqHU
Fr/aocR+5UdRBBSukXwFWwY1xQj/ePAV95uDVINv5swUsQfC+D4prawRC9q/4I/JLtij/zmI3Y+5
sGjguxVLMfbtohvvdmm5Pe9W4AcIXi0ajZCUToNDUBM2msoB3dAnmfYWgKnNwhE2XxZespMOj0PT
sqdkBpIXGvZMkIgFHtJhFFIXm8hhQUleSj4zQNRIWUCYwLLWtaiKESqj5J7zhiexvSk8boCJYw22
u5DZoil/alIzmLU661jLPqKvcjB18hTSA7hlrZ0tKYKixYcVlLLVdzqifHuGRvRT7pNzExHA+21h
HYMy1/MVetDrZB3IZUZHoEdsGxI79r1ICp3jiFfFQTaRDUFjgw+2FC9c3djHUxqD53pOMDiwTO6n
L/nTALZx6WZXYepAnBvfVZqArOhMr5qrI5FwRYY9Mrwa9E6H2DebNDYh5EGy6a/C8ffBVBR5XRzX
UOnWbkgiDl4x86WHYhp0Q/F71Rm7wx+BYmYdRWV3rehTZRvga9KtJdMl7P2ZvZLQrMUfovv5zFx9
ASGQp+zVYswlz50cwSk6bgSHdjYEZV3wmrYvclQjUV3CSCeHdhhkNulDBjp79KzgS7j+q/DFS71g
sRWV9VOHt/9QXSt4rB1nqLwuqz55BPshvl6kSi6fgL8IMK8gNHEf/NV7eT5RKsx2jzChMYsE34cQ
qSNPnMa8/SJYd9lAk624CRqI7UmXAYDgFoubjxFENm5/EwCsrcRncFUqZyOKdwx/YfwCelQMcsHw
0awlUm3TWl80K9SiDlSUhH4YKuxexxnOQaWDU0CH+YuwCwGjZqh7IPR5hM0c+FbRL+4jnBwsn4Wa
Dg/YpjRfUML8dm65BNMsd4gB4T+oOZsFOhLCKDfXQeN9VYkkRLdAtqlpcCP5dOm/Cp8WnYOcKhSx
ANdAjKbutfKWmgKTz+4=
`protect end_protected
