`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
eD8hpFSXjd1TN/qwD6KGU+z2509uzOtDyaItcj8UJV6/9IqXwmzXm49sQewLHmPx+zfD6FQpyw+p
h0cjnBe4og==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
L3SB3aFsPoBeCHEa+GJTxCywCdtSUeC6UY906VBmK5CfzTgqgVyM79kYm6BdXD2tikY3hMRbv08+
R63jVwCpRcJdeLJIbr58+pkInrN5jPNeOMVT4fdRP6mG/A+kbgolgF+LCX4UlGa6A14h5xUJIQ+I
BOJCodJ7zf2U3UPN5i4=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IDpiTi+KiM/mIyaieWhkLwbuAoWvynL5XwxHTZc9uzTfzudCoilyQ4oKu2/PRnV4HtTBM1PW4epl
rd9LP+loq5H8NbcXKhoN4VzhEypgVleSbFixkcTkk7Osf7hVTnIQPy+t0WVEWaONYL5atSlOleSA
iLuTn53tMAhqoF+UIInXe7RC0RJ3+CAVLKs9w091HN93vVUPCig/wIe/MmVL56SzFtGO/87XTi/+
qJFEM7WvagMWeW2rwVCOs/gjJhh8s+7tB2d3KXQb0D4ZLH7wYYzzwMxpSMKY/l9qmmdLA/pN12/C
iPZ8yl6wlb49sIPVnHi7OqJQ2eGqj1d8h/GCTA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n2PZpcfNvKmHdedDmvoLesUJQ2ikmLTmdJZcask3j7R5PdvJhsOsZzhHEOQT+y+b0Ce84yuAo4mV
4UeOAU9ksmjuQMNYzaXBCTRBJ/9azPVm62xll1YYsfPUMZgae2g6opjWLnzr6EGMV56mIb9u4U8X
dioOTIUTaJWgJFclbBdlYBvzRfUZhUXEnrcomCpTwcrv4UMGBsBcks4xQ+VsWhI0z+YBxuv8UqTf
QS+2qmMDtaorfH1LTrd7a5VPOQUgv8WS5MYce2LEzFY0oaJsKXIx2hkLzak4Mrq2XDDE/T1TKlay
SBc7GQ9QhEM8o6S7ecjMC7LHeDgYjWYfIg4cQg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
krxjXlF5n4BmuFCvmd6vJwuZG29Bt8Nn5bI9IuWdakXt77ls/w4/DdjPmapLT+DuFzJA8V6sy1ff
03PHzhJcTL3sKmbpnRLicE1pNpQUEN6NHDi/2E/TpQisox73hVgMAHEeAX6hqX1KcbefOndlffgW
vdyTXn2uGCb4mJOm/Ae78G/J0gsKyqkTdOgDX+5yow+NUGy6giW2aNpmW9DfgDvE2F9tsjbtkma0
VNvhHKIZ+lioLu2ED3lsQ0dnEEp2ygvVvS1ddppdBZs+szrgduYOXesf1YwJWHvIPu/HsiQFg1JS
xeBAqESdHqnBdlGvxkSDTrKjmnsbw4JF2Zk9hg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mzua6Bbkphv4HsiSX3MuiRoYKwYUU/2nOENlAhZ8kCE1xmXF0EJRVzVRAWyFik36NLa5qPt/4JY+
5OOnvTAVz9IgfyiRBph7QKNgFD8o2SyGGDtkTKv8LkDm4/74EU1epI0SWiiahPioX5BRHQJ58jal
8mrVX4JcvwfOukewKWw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XiHLmnwZFcNUphRjbMDiVKrQ5P+RQz18f+vH9g6AuGZBHN1tGDOOI2rL5WdjgG6AuaNjLBJefDso
61iBX4Uz2dCM5mX2ToGKZijqAJ92uJAXNBHrP8YWyyucNadYpgTAXUHp2cyctbsuZFUR1t0UIoEH
fCY5lWwHt8wMT2a7vQG/TwGfVxQHs/AUrny7rrjnKpmRzesIpAD4wEzfZZXokHGCwm7j5H5lo4gB
VlmEIaqgi/Ys0iqQ6Ti1bze5P7OD90PsZwx121NkJMhdfC51MvaSIeBGNoz0LD+N2yNJZGNhgKuP
VKzat7Vdb0PqaMfv81PTPvMKxpMFQyzOad/byw==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 20128)
`protect data_block
EXHDKdmWe3KKmjfshDm7GGy4szG+sx8LEtajOqsZ6UKD1LBDP09PjD1QI2l4XswXm//UnA7oTX8A
vIAttB7KTfmEWUHD1h8n/hzkOHrURSiXLZXQXFQFzCmBG8gsvYlEqITBVs+C70RT7Vj5kKx/Crvt
A5HVRCwFPqLb9uCBgsPpCLQYOkbta55H9IBg3SHCgFypk/wcFTRaFj4C1ppI0ltd7Np/GVcIE0lE
lus4gqvoRY4xpYj0fh2lhjqxJ+L7gGh16mcm1Tp/OQJUY4pWo1zPkEUdzl5RKdINS42mqCLh5B1+
oRpo3O2d8ht3Vb3gKRpB09Rb3mBet0yDnf9dOx9EMXsrGHOy1wwxFi+Fmpyd4nIL6rr5mNtjUCZq
LxCKDa2LbGc16/uGZr8enlE+/5H93jtcNvimKeEgKaulXzpo0ocAw6xbfKLyy7lAwYIlLCy1bhpo
cqJsGXcauVaS0Jdxox5ErnpYiLYRcfKNc7Y2qwidWBo7GZC7dWeFZG/8XVTDbNQr44zzrdsE+300
1m6Ni/sytTgNqxwnjrwql1VUh0OOrjJ0LiQoyd7C66YfDUX7l2VpOSlf9RxoqkPa944kCfMdswGp
NCGJXv/IRc5dzidVy+y79jGCsSQNQoedps8T/N/76hZTwlstaWAbzCrflPc7HSSgrb637GlKBj6T
UOuokEs8E6VgvxaQCmn2gFNfvbdDLAVIJJgwVLy2MhTesIZ5Y8Q47/pfpUAk9rYv0o8z3ejRiQ4f
dhz2lY58lxo+62FDvOWEfiudxY+mWVaU9ut2imyU0GpvlviPKbaheT+mg7q6y2HUA9//1Xnaz1LF
ZGiMyYM95JNVE0OsKFHDqoZ4w7H55+P+HOQSnHAGcdjQzYpHVWatHNzMEgsZuLTVxwbRs2y1sQxE
mG4spFOPJoLee/VEjlK0+GLF1D+o/GK6JqCXxYicnkVcYJuJZf3lMO9eaZwjMI6K8ksBXASSgDOv
Dw8UqQltfxQTKtmyzejEae69QVjtYkntzxVfZAsdoofBEoKZTJTc/tYiQbjQK+RNKgwPanNxjlin
P9U5J7M8MBoYJF1uW64/zP+jdIVFhnLQq95le71VqTFUmWKNWXdA6p6Qg4+wU4eN0/53yNEHA8U7
YgxzVg6vufJgin6BPelEpx7mEqbVDLVMId5m5wEQkM1ODPJu3ojJ2YbAQYa0m+DktmrROQoCFyBZ
9OrRQhek0oc5WkzT5y5DZecfW1FafFvc7plVSC5k/mW1FBcd0kSml2rd0GxvS2xDRKb9f44BOyQm
mEqEHn3QHgyFsmosSPAjkkjihPv+V6DozDLwGOxknNy1HxkGZuRQszllylAFeui35DBNQim1FokX
wl4DcQOA4/FG0bcXV6sM2/I07Uu9XLhm9mo+kL9/z75K9juQ7Mau637FzIrY8qEWjmNMfcqIzUU0
4g8nCo+t2gtObNM07PwWOErE5ehrPvlbmUMSaKjWwUoSNhy8tu2ebRLhxTPs+myBUu2L4lrIjqzk
r1fB+ckBPYyYSSiyewuQl7s8wwPTndo6kcyRKJxK1Lq1y03C9pk09iZKqpE7nBRE0SAw2yepKzyy
If9WFHdB5rEZSxPQNBbr/vCkPlauklWAhvqPpIY8/G53oCUUuxWKaTMDQ+gS0MwueY/mGKQXzRef
bPfJ8R6D6MD6tiVSX+DZXaYFMv0js/3+kusien9QJbyVFVCnUx6sQw8zaTtLgDxgiprhoGasNy4/
LiFoRvuIZf6BTNj4Hu36LaVEnfLatDTbDcfNlVg4NqD1KlOXCehJ2//FpCLIrQKHO59dl3/Mqw7G
GRX5BkW5ERy7ThZ/MVG3lMqAcaMNKLYbK6GFV6ox1sjwL37SPOY52i2D1Dya8/o1rrexZaFcllAA
PUSbPCCtEEyTXGDP5iBC0HlQf2YGNlLYodlMLQRDYKrefWvo4Girmoo6zmySBd1jPvY9i8o/Pgdl
CVVmTZj5QLOAczjUjkonD5L9yzdBD+W6tPVIY6psNKlDD8/WmtuZSlw6FUiZ99g2n9ovDSdvqYNh
bw1KxRP9KnrofVUfPqhdSsq6iVLS8BntXZwOwcooIkAmw+pmsz7sLQVCsp3d6t3zSkmkapA3VepU
Fpmx7o6sn3mH7g99CFJ48mNsbkKyW7KSVnCUIqFSYfe6RkbOwm/vuYN3yF9dj9UPqUIked6hxSyh
U8xc1Jx4RzTwF4AvMEoOaD3uMxyrWAjgEFkVAopR4GPhodtnd7O40WGyS5G24+RSukGqnt32WwQ1
Xp1cBHAmUCzm4hd/k9vSeuoIyNvS2ljPsfj834nebBHExn9cZ2Xu/n29NA+oJOdQQaHphqwV458h
7L/ye6ErT04F+Njvjv6WW1exEbSwabPrRyNq4+GVKS+Rkt0MD9LquyQupKRIM0c7eYirBYsMGHec
ztzyL3i6yhptshshIkU/vTfS+tX3FO9z7VGm+etWnae0T6TLY00YHgHutiMHu4cbIS37XeBmBcLH
FNTTMdwm6+oUIdm4A8IRRl9COahEAq3xkaBR/HOXWIQdMAYN0HexaqQcqwkmULkC/jasGzkdQbgm
cu36XuVJv5rHGPiMFhn3toZloQivUBBYVCdZGAbCdBi2oMxzKMt8bR7AeupcGlcCm34x6Mz//HvX
OPcrLEEMNZXI64LrHDzeCr+Acwv4gwi+mQwIKJefsKL1ggmGsfKOkCetjk6y+2uw7ca9Kc6QJwPS
5hxsYEqt97T5MLSTZzdelILQfNzRBsO0+d6o6nXtJDgA3BudL8OigXiNSRw0BCIdQRu8Vi5smEii
NYgkbWhUbLbxvxXtNSR3LjfErxHXM1AZ3DcT+S0QAEi+QPHj9YK587Mnk0pqOZwdLhhfOnaYLrxB
DwuXlhrGznAl/llduJRgTjDAkphLr0lxjyoHP4zDE0wBM3P8F+m+Gi4AOfDKd99teo4A1zLdP8/I
rOHRdN/DA1KOz+C/+hzVfQwFlY3TvPM16FpXRqhwdT5Mq55nHiJ5lZNeJk2BW1UxPkYBe0ZcJ/7p
TiW2gYku+nnOVxtSNVLYjqgyH6Zhgy2sAqYz7+VruSnQCID/obBShFMNQGOb9TmrmQIHB7NxxCuC
aSdx31cb+tW4V22XpQExfH98/zQXJakCWzOe2cUrIksEm3lpcYi8I68EAIsTQ+6o2aJXwRcfWCAJ
b4+9EGsYnaBApftYsq2AAMjRhea8kFLKdh1YsjiVAC06pkW6ypYtrGKQwz44oPSfAVU/IkcpMt0f
vprP0yueYjhuotNIl3PX9E9hXGsF+RiPiOMAdD+e2RltBlJm60fFiMAerTHInfYt1j2YQaD/Y9OK
jZn6wSWMY6MdJb6x9qncCmuPFi3SWI7q1F47ljMn2TE3Jj7LCbA3Sr8PYWSPFx9Z9vuXMU6tAx5Z
z7dTNjmEek3WO5jJRGnugYPaal0aMYo9varSx0P2xd0FftDe03Jr5Yfub2QChGzk85gI03vTebTL
XPsO5RtXhJKVNMqqqKYDszon72VYI/aIFXVW9LW//jgMetqI2EqO8z9C8RsCY1299vtBBE1TrK5z
m8t5BAdqr9rcuT0JZbbGU8xHN/5pMsnsSjUS7gp12JTUTiPulpd1npvFAAQ+LErKE9xJ25vtoCkO
4quRJGztxlKg5M1gUGsvt1HKu2q7VYTcYh8yXHmB+/wqVJfsnxUk28lkrR/Mo1k3l0S2M+H4cPHS
Xgrj32U+ftmqb4nPK0czwxWp4ARkHWwlro3QXkGxGzxQg1F3amCAnhBCeBrAzKi/7JPkMGdhjqu3
bJ1zHcpVQDeIG/U3TXrFS8+1/zzKDyhJnjz6x2goLw8W4RTCmZcmksGQem9ZEhuDNueIQuQrU3RQ
h7WNzwUgg2Kay9Q64M3zErZC78NMAtXaNbtlL3LWyYuCohikNI4SSxvcODjYTTVPZFTFDKhwLZE5
8RCVLoMqQHZP1Y2/vyRGnxhZVwxOphwrNpFNq41nGbpxFbe4Mae/2/UBxFthlYsl3yiPL4peORT8
U4DaDvdQj3XvaKT3pLXgUT9JCNpCZ1zv1V6RnBfSzz5YAcGrv5Mv9rlnWrY+OxQTJe7zlvzXaNGO
Tj/uMQJ+a8EtijpBXMAxL+B1xoLPp+eJld7z3uYoFAoWwJxQfUcwEOBAYimIwYStideMtdCfnjOI
TgenYlazWmT96BIOPeRfVF5thBDNmiZO3ly/CACFNbbm2JLkg9KQqrKC1E5i426b4wzOheCpJ/tR
c2bQqGsreIvOahrj5xel4nGtnkkzip0zasnaiNakija1U2fZEO8FwsbW+h5Ip+TweJTl8+czfXqA
oLLwqcTjJ8+UIgLN19HEb0tnA7JDPS9uyJ4llx6xohTko1RfQahjsBtg1GfRDLYLxhHL13JvRoly
DE67fOnLMbpETOApSPr8TjgsaXX9epH5ZCaLwoko5+Umuvdf3gdMYUHlaGtFbhzJREn7/TM0km/B
oEKP3G78LPAD+Is+tI5sgxLCAVCEphkB5HnKwv+EpyORy88LoMlrt/z/zS5+0YT0PCGoOIUlRT2I
mviPYgZ9QqGqVSNc0XZzyAilIxzOcd0vM5QJNNpuhm2mw+pTETwJM2FNcaqCUi4amv9g80XLGAWE
T2kGezR0U0uwW4z75MZ9M2Xin8mQSvEtQaM9Dm3dg/OWO0eVV6Kyv8XnDUxgytrfiHAYMloPe4/y
bEd61G1qR1SVAT7ErDEs4zIkplSma9aMhiV43UxECgSXr9pv1fyjeOzlmAdp+mrK5w6I4TNSYe98
VYyVzy9IjIlYj67olq9CJy5OCeousTxWQvT3QFE4cSEarFMWctHh/Uij/2QhDZq6s40yCwdeLa9L
V4hXOPMuesfrM63ujY9oKDJV50YTjaH1MeewJrwxyu1Itfsvv0pCT/ClhhtqkiyBzY6xZiiyUDgR
VMwULMfCKixO0uYISy3TJIdg86SlkrJUn661csXs22HcMY1t6xrSikpp58dOPkAzl9WLCFwp8Tdj
SrUJox9ixH4zcOGcKrTi4rK6nv99vzgf0eiI3xIjFwDAjMjuOo5st2p17b8fcBl+inguIOiViaJc
3MiZaJeNV4nH3VHRLEIW7VEtaSMFKQISveut6MWFc/bROdsEs99uqDQ75Kz3AHqqocqI311i27bF
4jHjIrYj6HgF2ik7lDDX43rPR1MWY5JMaXtoY6X384G7Ydfrk7MyHf6Tf4BvETBdDVq2ZvqiJjS5
SrJF8REsqlHr24ocIYAetSCKHtg/PQaZHjBlJYgeeIJkmtrt1yKSlZ7PvysP90MKlsRlDH3w2b0H
TPayWa5DdNNI5dFwzIRnik4MiQ5aRGiCHmtaRLAMzFfT2Gul48GT42uwnVFxBTrdB/qOXhlvhiT3
C3W8Ahl2rY+1RjFIihIZwuyXuNu4rL6pF6T+9Fx1SWO9O43n+0h9XCXg8Y8UfEqcDQsKRjHqEs3S
kOnN8jPiadxyVxiwJ/6sheYzppyi9OrO+q2jmp72rsHt8X5ESY6pEoKeEOyfx8+N8b7HmbZb5WWW
JYbRhUqdOyRsn2tUcYa4wND7qVMtpROZeRmHaSW+OvpdNsWbnAPaJdjdeEqf6Iy1mdOrw1WhfbJ5
YgtDH74U+vBc5NHohkP2/PBI4NkgdeoR0Ktg876wLYDW+7f5pCKyy7wfK4mXiiaPqh0YZgF+moYi
yyPhe17hqtjeiyj+k0aTU9jGvZeaJoIYgbMY4woDtfEwH0JzyGPHRoj3Zi5B8lLoO7K+ds7fwmq8
jrZUkXi8QHRDmsL4uoj+zIUQ8+WT/NvdByGcxMtIUTqq6WI0dOP/aBawnPbfNt7GtSH1I2lqXGWX
w9FErMBvdgW89cNJzvVLIYCorWuPDXGucRQbRbbtICnQcqPAflWjjcRsgly0qrkqu/1aXMQSsBrp
BP82N5p6/K/0SqLBIW6HEptZmusm++PJY0Bf3Xk7J27MP3ACAGA/Hv5tsAWAoNkUyleNpRgvFODS
7W6OWuVu5hJpqJJYDgoSpDtBSzPcmQw1G1M0b+96vKQhFLAsMSzLumOAxuSFy6n1DZFy6FQblRa3
AjHehEATlRJSO/v8t/5JxAyqJhyxd8cEBuDJJrTy8NBBo8IBbcdeob9o4X5W7NgSh8jk08jZbmRe
0xPKCtrHDWn4u4XX9pJ4M1fifpHNaeZId/zCk7gBVrdclDrrUKNP1WJ94zRhDkhwPzYRZzmTPqzT
avzWccteLx/wTRiR7cqeWR7BU01n9fW/xoXexkn0bamBMNI9ODdrvMSjffy573dz0Gm+hRDaxT1A
VKmv3hdZLfRDemGBv8LgFVrujgyYLCylA3MsXsPwjmX3i0tjf9b2BxXNGwFBJdpInLStoSCu2k4c
T315CRXRKf9vemV5gTBUVRA/sKNC4zjdvg5sztLwYwcPvCd48ENFvVK3anHwLApcv408GTMrGx3s
5vjCVfuuVGPT0RJmUE4QtkhGRxHrntq9XMDmXTBwHeXg4WKkiIBRsrHIg7OPfNHMaAtkQIAROEGm
hwuhrHHB1KQqh0DysQkwuqDcMxgiCeloy5SpXh6TzFuwVdrSG6yegt1kIvQLT0awzfsvToy57i3O
d+wEjK8RpypQTbSFEOiWQswji74ep9+YDzd71DXaEnu8/oK0CeM3wRfzJcxE3KdhcWgDhkmPRCNf
j6yJxusoYeVuF9/Uzuh71xnFX/JM8ZX1neqfO7Vavsnf/B8kmJAIVfHeLYa9zC5kkElyV6pKEMJK
KfWfeTAFXverLb86tn0U57CN2VDJhW9vZ1c8cvSp8PwN6BlTryQX1xXFOhGF+E7QOPDBN74ZXD9g
mGvbd0qBk5oB3sDc7AEbHzLOEpaNL6O6inuLmXH2Zk6iASJtssUYG3USV+j5VHY/weq9f8PP3K54
6I457GwpJS20F7iut/Lr6p9nDPoCsmFfzS0mjWg5gh2tb91JsPZrkGQXSqwR0q2W+tcb2p/7cDOc
XVz1HQflqbzmrGW6KW3lnM9mbaRSIP8ITsXb/8foy6RRGNSYEeNJDQVBqGLIhO/2leqcbOtxRBv6
eRGqCdAoEpVbIiG21/D4H4cK/9xQco3jaiqxlawrL+0qS+6VcZANKNh/BNYtOzfEkWg4PIWHGjYx
S/kdHeS9NPuiXcx1OqFERGP5oRxPKBVq8oeV4gly0Ve9WP0dFu3LDUgmgsnD9TDfxvOkyvIX4aPa
jjjEX2AQiUQL4GypnWRzuCqMuym+6eTUz6xlz3+1rxEZEL7x1kcp6l5N26ox1tAAmze1/v8bDZNd
JLxVS2aQW03ppVMcL2S5nNOL3tLNgw+Nh1OpgVpluCOcOBUv3WVzgjDfh4f/M9szHD++uYq7PyMq
PMrRNXTicGwbDuODRAT68W1ioTHSrmL0/1xwfcbUnayFCWluL/7awBikLGWStPlwD0tqC9n33Ipm
d3a8UA7uDu3pumwgApQ1krf6Kkn0ZncT4szsDIAKowAJQtMvIxrMLrMCLcR+OBypVmNt2oHkDcx3
35w7qg5XMbrNF2UYOPXRhg4SbfdLy32xPgzZQpgwzaL6LtBvtEbKRJ9OyOoHWCHiQJ0sFf2V/V8y
KtvqrKpN+f7mjdTbSZ2A1qsjqGTFScBbU2Kahf97JKIpFCvy8O3UzBDLibHtGU9BNB1FAcUHgWzC
8s+vyuroncxteRnhYmzF+hh6MHplxxcDZmYnE/snNRvrrEDR2xnrlGFB+hcZG+NssV1VXyHA9AJO
KNBXZryQr79Lf5KwdF2V86gbJA7RkTD7gLUiPMKvD4YG5JusvVYCoTSz4AovpgIo7YZ9pgYd0O1m
zVAisYV7pRw07q4YqpcAv+7uRxKy14tuvtqpV+/7S9nfTn30hI54oe9ZumXAqMviznkG1lZqV83/
MTgCQRZ1vNE0iQMK1Ebjt+7gEVhPomhgFawNU+FLJ2llrAweEyPPxqxeWcpkOJHxvtgV0X51jo6P
XjST6V6eC40g6g1RiAMzO2LWeb2izz0mU/o51VqoF7cJDssUsUfY3KCnj5ipn8ONSJPJP0c3yw4O
0dKtj7L/qiJ97Vsv47ZySghtrC9YhfptzfS9JCVJ6prOL7GhnxF6YzpRbTT2hn+/3EAveCj+mlZJ
vgwpxniPhuI/D9qXskTbqCjkM/yLceaDPHM25IOo9Et2gYqqsPxVGQHoE5x1q08/RG/UwETuuDwn
GBq7MdlLHwGOlWneIQvUg3ekVcv+7DDOggdgkd4ytaE95d6nEl4chnZXq7ozbYW5Yzj4qdf3/tQD
Laq4wTTMrjnKM6ltVTafzSdAmxnvWkXQz+Xnx+r+3whTSeEgAfSf+w00hxexCgkEHVtlVt+VeaEh
rxSDZLa2mqBJNLVOkOnYbBMdAmAeY7koM/CUgveoeRj5DwjGFoN25yacVAR3e3lDFRfi/D5vrBlE
GSbU5cBhSWr+b9T/3vzmaBsfwRdGynMMDvbU4w5ol1LcA60SrvC49Dm5lZTKW07wKzUfPU4n/Qvn
h7XvwDCIiOyQVcq2I6A1uLxREphWfc6XaYni3KQtVh0V4OUYu33ZSHGDLBmax/REP7KJynVyKsfw
vfCGMwSOdwQKbkEYj7fIjrx0vSjbgZtZzsVJPKugjrw5OkormqiVX2RHSHMLz04RVrMxF12oeXfB
FNHmZQ8IyEmXzpNjXWmC8B346NBhAYkNJbIr6myaBC54osCWmGFcEVfiAdcSlul7QWnim+ffiWnT
eFga64V5DKqW+C6wFuY5+M6Gle+pJrKQCvG2aBdZENM+Z0syDxQ8DzWDkZiEoWD/uhV8Zy9qLhLD
fVLzH7keQJC9pwKadbLfBK0jy51Lm4XWGY5JFMoo68FtPNXJcV3rIax8X3t3y7zuhKbJeUCGBQ5+
UcCJY4DfZI0QfuV9cNDjQ3G0PonXc+Aj1nhn6k80vkSQXUEBieNA//Xu4azIVe2bC92AiHJxnw0R
Db9GEnHlJguz50m48U866OuWFJ+em2m12W4t/7noBDvNvYm1zzkzp2QYwqj0FY9FAwuK6Ldc9JfP
4/hIMewOT1fo9DelVm3W7Otfsr6VSmo30ejLU9gdkrLMx59bvyVpNoePD6WGlqs5N2Z1IMacZrYr
EJuI01hvxxHu2N4qr81J8nSz4oAo0UqUpXZ1ZzGAkD1bTYTxIfGD2wBUFxwLwkr0vfxAWjee7cA1
QfoR10oEhC87MMZh9kEZ/in7FOgG4Zy3cOSi6JIjeHfdaXsyvqp+vRrLoDHly3QAYfyBKyLov1Q5
htlv1wWkAO2mgSyl1/Tq9Jc5NqhiqEqEuil+bhMYKxryzQL1+7FOSKpUCD0PntIHQYJqvBJuurki
aTjOONzdBpSFzEErUoE0a/0Y3yHS1DRTTiJTWYwtMgQ/KlMGhVKCKFjBSDQ5cdTT9WNlfCMkE9o1
kn/uBJI+nHOWYVBuRUCkksmvylv5xemJKMpzU6PTQ8kigbXPjWkAY34BafoBkAwakjiLvL2wHGRC
frcObZSN4AgZVjkLl8vMqd9uhEfibf9dHaARHJ/+azKkHxkl4jyvz/TQ3swS9BTjkiQ79MgAAH/X
kSgUMjwFBiUUTXWes8XcTSApMVrcMF+p9YL/qvbUJ6hEjmuMx0f5xbQy7CdLjDRp87EqbRvUoBmJ
fT92/uCX2qfVReV9uraPLbc9zvEEZngEJBV2nfJ+KZPth8MQpvSUVRQmnT/w/1gPqk2jhM9z2/bP
Jm7rQ1uE/exHzg56xu2dknxt/gkfrUW8hr8408FQTJdq2UC/+P2Sk3G7YJmDJ54KWrP+7CXP0Wuh
6MFGiLpiSqZ/SG+eMjt8O2JcD3yUXVIMnlEtKxPKlCMrqa7LKnWlcSWP9e4CLyP8BBenHAbdGMve
d7uvaRkZ3JIrNzQ1Z9bjYtrsuiychh+I4X30nf8Pc+qLxZ+vj7juHiRRDh0SJqga34kSX64w7D1P
Ac2qEHAIX6OJUfDnfCBAuNqOmD/F39F5b3QxFORB86f+pwECUbaULtkeTSdUPBrNTThYo/nvF0rP
Og/oqXaAZmO/y4z/kkSX0dKP4ZOIQ/sepWkZM7MDNj2Gpi+8HlwRX4GPUEdrFU3BMdHpoEenIdr2
huKk4n8zV5ZOz3WsePPsgSS+zTHCJO76m/Aymv7Qg4gT0NBtHueeqJaVvYMpRUILweLBllqVSrVM
7Y2K7eVP6j4fI6S089MqMsHJRpgdKQhc8L40uKDrzv7LvTR4IxaCZ1yRT93R7GqIfsOZEFpUGGxN
mPYdXyoviG/EMI1YCAlDNjtB4T80eicXTryVWaGZD3QJPrw56/oW8Y7UACpLm113he5lv7bztrq+
zbhHN3IMhqSGXj/6sT/aajpkmnw7SwMPngGdgt75vYG2HiHCDFQ02ou4xkro0w73bG5YhqW0FC+8
Byw4JccLIoDQ41yaWQ++DYcsRiW8zxmbRHZl3LlD/u2Jh56bn8IdgBi5w724+bW2iP6mC1nzkDAJ
gTketMdJZ170+e6OndgcYg3t8EwwenrKzFCdcMnD/bCS3MeJwZ+DnmVrqxOGKIfAJpPp/t1OpyVJ
PbGHsxSlYdCCEublVy11DbR9HQE/OHRjY7p2vQmow1tZQMjpdFYkspM1pji1/xOzvSKM/xK65MB9
rAlazmXhkmuXvrVQO6P3j3e0CEu1KW3VtHTDDfzQokgFcVeOdadiOykZ2ffa5Ym1Asua4agcYORg
5e8x2aoYXhFrwbt4JNaINELhPUufj1uOFsEHfujL8RmiaYfdEqrRk7m0yh2X/YxjX0sUAV889H6t
tyasZOqhSQ33WNRJ8NF8VZ17NPGBLyL73nFd47m+RGns7o7d7yh2P5bMCoPK/1Ob3SV9/cTT0Nmm
vvfkgBzwXCdJwUHCjtZKcMU63yW3TglRw5sMtkzQ8c+CeYjrz1SqU96gy5wcb0nMI2PH1vPndNAw
l9I6TZDu1q9MbCIal/ikBc5nc2rjHWE02oUG5LUbjqa0DQE+LO2IGOX8IIE/8A5b9DwMExvs0evx
4qVJcTS3TJVNxbXdYFE8yf/vIz1SXY5L3FePpW7bYArnyX+ZGDfgaXKPnLXAfLZlX7HXUOR+nboY
p4VJkU5Q2ZFlWXRA5hear6T8j2lTh8P8arvKMFi47wSbwqiWF87YXeZqMG6sc7emqBE/wPeNq6UT
MwIlL+uka6zvAtRKBM0ZC0MIXg9K/6ZAixjHuvy5Cq/CldqsjvfTC6aUiXLmlsbj3NSzgyElgkG/
KMOHvt1TpaQ904wREYvzBS5IVH1SAvevulx3mpC7QPKnsOzmbUIpEfbB5kIbZ/WzYnA5Gi9qwo+X
poip454ee3Ku1Jpdc/bryo5ok7/ri/PCAwWL6ez8oWHKTfCjKd0L1UAPRiT9LsqArSM8SS1u/EEX
cGPncl6zMFhZdQsHaLc61jFi+wTDz923VUDVN+KMcrRnKwNNMn7LSLPgYibu6mhXTsIDew5Vc6CP
R0zQuuao7LOhj7fJTY/RdLvyCabh1RAXL6u3S+x/9A5QNA0MlOM+9mC4DUX0UeBB1w9wklgS5K1S
/yR0KC0nFEriutAMuMfajYpNRb803KhHI1u43ypWlA5SmYtYFVqphmRr7/l9DxRJ3aoO6IF9AIFh
oP57rnxrVgRaE1pBOZtNFWMhmA/byOjC2ORuzi+m2mDnkoVmKWhJ8aZcJ4GF/EX1KdNbiV0nwjYn
XlnRLUQoHQifuWQditS+yZ0Qbm0AfeVOWcJ/o+DWWutO4u8jNi6uLnMSYfOZ4Eddsby37wldPy42
X+FKIx8xE810f7boVnHOjFxFWKVTfVY50aomGTZfLraFdKL1GctE4mse8ZI+1jZNA77oi2Mol/0F
Rmjk7VH10sETaUYFhBADjhXOiV1Kx2YfoiAFfXKiPOU/tJWg5wpnJ12Ouxv6dMFKHOaGvVMnSaPl
5VloOaqvLTNC/d8wi5Q/3BUsw4weHWRP43Si7TtXuYDrkFwL/oGijEGYgukhdu5ChDusI8tO/IE3
n5RECRaDZAlkmtPp2Q0k6RyG/j0KpkfSN3J294GfZ89BcKOY+nr5YS0qeyuP91q86hGVm1u+Thm/
qBdHFqMMF9gZF5M/5IN9t5nm+6g9pKuT6VzLZsMOMa2o3c1LVSj1VySgmZX1NHRkZlKaq9c/Z32k
/hVN9rLkr8EP9+8E0/22/B9d2OPGEqQevP3FqVqwE0vAISs1BF+/7gA4rFiPA+O5I6/4Zl/1OLNm
71er7E8pO07rFPVJk4ytaSgjUikH1xKOBEog+WF6vwAJ204HmKol/yTsgWILjWFfFl/BXSzCGCfO
7ruSMUCCeRULw9NKJyhzx1PaCnu02wsw4XvMyvpK4VrlylU/qSiy8AYlZh8ZAfpBptiWZeP24Miy
BeGJQR/TaYxoATy02gURumivqLqIw2AW7XHEIC2V0HTYU6tC7k1fyuiZ8j0v98GMGLyRN6GQCEgL
U/w2omG5lD9tWFTHIQGglDSjdVbtZkAGxGaeMdQA67nkrUacRnH7NtWweDT3s0RxdynZdxZZB3i8
PAab5Z8I8h8mimj0IsOMVcALioAjEyitDkuEP4FuCiSnRwQo0IIB8kqTtJAFQ/BXp2B+V2T3HzjK
wnFK1wCg/ZomTabJkKUEU+b/UjrNr5TxzXtHhLHFRRuEBCjO8eZSDjiXkP/nXXqQcokje8iNObDf
4vcW92jdETfJEDrG9UsCVZrbXDrGkls0HkDet8R6xAJVRHt8iez1UwDw0hcvZxG0PyXE8mRBPjHm
H26k3S8PJpvkwSqMK+HfzMm2X7B5rGcGj5A7lQ45UyAZ3meyDcoAoRpAa3IC1vy1rb5QuV2TzcVO
OUwgqSy+EJvhkxL2UfY4STMiObo3riNIUsPnpOlZf502byQetIQCh312WC/Z4jXDEP1yAnbkDZ6d
8K8RiN865MmWgS9dPJsZ2imZHN/Ji7VN1qhTqwgtdSoGwOw0JgRw0pTlCevtYR/kL3xvW9ZE5jrW
jWZT3bdEZV8nK0+Rhdfurxfz9uOkQgqanTAJaKEFmhjexXWPZR4j6BlI9ZduTu7wAk7lKOMzakjM
uIV3+rQigSUS+hifRvBd5+HPuxwSmQSrsLLesu+5gu8XeM3NP7DJd4zjcRNpoImeXeUlnAoUBmTu
u0Nmp6oJb2oV8XhkibrMQtYBhU9T4rOzv1pR/Yp0vXu/U5aS/VOIW+vwrU/0LaMZAyrx9tz/Nk/l
W4AV5SkYUQknlmRl1hwnf9gYXSoBKL42vi/5FeIc0WTqm6XdAeNF3wwPF1WeKj0hqdeeh+dFLDZf
2BUaBj92q4kmxvehql6fP7tX5/7GiqXgB3WzQF3x7DkNnEFMnaxMvncMs45RkkVVdt3m6PmVugYy
C/77eNvnVw3UiKQ3WDC1iER5U1nHYetHkyQTn4YKZtb5xVf6AAkpXZSLwK2UyBCPhRh4vwPjjoWp
/6BUJTL53Ps+YnigUND0G7A1bz1tkO6eJAukt+9TuDPuA0/4OSOxWEfC+FjUwHUDPh0o+Pp4Gn3Q
W8zegoce5PVF354TZhVT3bLzeJ4boDjXbjQZlYpWRzzMPqUzAy1wReL/iAThNE4qOAZN+OKiHuA9
e6LcNjZUEGEXgn1N2wFZGhe3Ac+5KiK5V9mdHuwyGbQcr63QfhOayrbwte+Gd0kRSviWhJCmRsQj
iCc4W5mfszuSReF3pIrkn27AdIWoA3uuosEQcQwRN3xOd5MrcupgDo4OaR61mJFGTrT/SMUFPJZ4
8rkimo5heCJKqVEDhHiz76Ox/InQaX+OFy+BQaCX92OA9znwJ4BkPi1O738/pxi07ryC3WZUhTYO
ln5VZ7oqzjex38fPcaTQeFGsl1PRd+MyetH2shdY9WRlbp/M+OXTwVzFdvPqK0cuGklstsb4R1Yh
ZorNoTco4MmkimNWda3+LB4kwABWvwwQuSHgUqZHW/xuXBqej0ZujDgDh8WHEoQzEk09lL5eMy7A
/5UncmIqOP7AcRBYi3jAYGuXieH2RcHjO94v8Um2sa1t1h3A8b6JB1i1T3wuTRdp15xnxzUXW0V+
mksLxKX/6ltxDIi+SPGvhNIpfE2FtgFlaFLqAL7bQK8Pv1tfrAM7OyYnYD+F5/kCppa4fFrFc4No
PUf979UZBitCgTzYDCcKjXHAesPtMpvrJboK4AKb+yBl0RsWG7EBFjCUTArayyqzu6vma93OV0kX
1i3OMfHYbuzLpib9Zbexu5MD6YIvKEzSBs30+1VG0LeLm/DZx1zeLHgQspyr4gra58IOJFElmerA
ar8vEVvLImuLmz4UQ2tXlmN37pLXrOusdYXhwrtw/Tjc+Jj2Ny1oRWq9+KGq0YoamABf8pcmlC3f
csmWHmT/nGrdu1gNEBBWDUv7NGhLS9PW64TTioiaa6eOKUP3EqalaRWm/7TOIngrQuDwru3qFOJ0
8K6VTfaY2hgm2QheGyXZHotismYQGmyisF+tNFCLrotm7TVgUQUJoShFU5Et4c3MQ9OgkUV3ZPfY
HlwjMRUAYxIcvbJChunMyMf1e9S8opq0/lBbsrg2dTzyzbE8FxA+t3WfEUwbd/GxUeCMqM79vTyX
mkxoLKaZCEJP2pVi64cPppqEPaInTquwyx7Ui24gBanX0SJdojsSRLUK0NUOOhh/hFvRwDIFxIs9
cEBf3j83rlfc+CKplEL05lqEfIJCYpotBRtxsI9k/uWJLeAsMTK1Rrqqc836k+4VkDqoQLqmFnai
RG+ErlbQPDTAKW0wWFgIrZURbdIT3FSW5PLExMriiJ/RbicpBE/O95Pv6VdFyrowofU74CINS3cO
51YnkwysN2EOGxS9AFGGHQNXOsZm/5rFHy4ZRqyq4ccouXvsbYdUOZzuBBBJoAntdwwx2TP+x//q
kCpfEqc86MDH8luRez5FhR5NOSSnFH7qrDxC55ZLl+1G4dQ0gatB/05GmvXs49kUEVIewJ7hvTTJ
Twty0xlJUSmvcmXYyUiWDLuNGeeVs6osP893u/22ohLvkpgLYkJJuONtQ3tYkjZvt4F7VLr36YxN
HhzMhRWVisVABAlo5O0mtc9f4SiReu4E9bhY++EqxgKxp5oWIn2PT5dtmfB6+09JyPY8+gvJwTim
fydxQgPIDhcYQsBPF6tjc6ifLUIvcgrQZZRCWBz23XwAy0metNtuJ+REFyr4nQYvTMx0dMyjJHi6
/lX28FeGQ2qxaZoTKe1Q/t+S+VknSImceGD1eb5sVzU4V7I8pYKk0ItDVKFChdJCkYR+G2WYULBp
ce+A0kednRbwyliZBiz8NQy59c7DAIHiiEQ2jWYasXT8S2hZDVqrB+5hmUU4Ere0tF9owFp5wCQS
bs644tuy5Kn9HQSakZnuS7i1JgTLE/65fovoJQOvW28sCyninxsXO0Tq74Ge63EVlHlmHru/9/DE
nUStR1Pn12xWiE93LpHborDsv+V2KkU9JYYPVge982wOnYizA+wjWC7p31EEYKJh7H97yXusScKC
I3eWR42t5gumFqFrqyx8FzJiVVNyo1SnUt17GPhaBgvsZvaMkgVo9dJzx6H+KtlXeZpXiTMSMDXS
FWloyE8Z1te0VDNRpXzCyrUiMm2bfLfoX8XuDOzYQxHbva5PFqGeJKjR0Gj/wVB/c5Nfqu7sZ6Vp
PGLkAS5MfsvMCREmNGdvw1hsKy1SyMJRxJVC01aDhUhl3wOfQE4GYd3Fh+zj0qQNzsPM/tAVHpiG
2jZ+N0LYk+ktPGkZFOiQjfRhMi/uvX5zDO2gNOT0TgoxgyqgeqH5/UmRJ2x1Hf80ggjPRu4lTTtu
swI+l6RooSRZr4A5HBYY0p/3IRePqLEKjpEZUEoXmM79rCpvgKi6q+j8RWW5o/gvExPeSfeFbNyB
geA2olC3fPuHu4SL/O6OfeXpOf4kcjHEJNKF0y+WkPcZFVrP7I1AiDP/+ErkDKya8+Qo7kW/xxCh
lg+JvaCetqZjfGfYxXmFPYQKe2VHeJBfAEI4dO8vAkCncwB3FLwfKgSimWgfJRC6XjFKdisoStoJ
X9J2t9lny8saoGtqjbUoxdRqQT0yVFHq5YHL/foMrGWGI5EYj+SILD+xmXFEQZiJysEOs/Zs+pZZ
yKTI4d0omg7zfkQ6XgdrZCE/UGSJWJNEHtJRorJsQ4aMkgERmDXT9XrP+W32DT5kK/8W1Fbt2dem
W2EGfWpjrb6bdXREqS0RRNHlNF493v5IpBkMy+19CLWletO+P8R1X5TFxvcAQJYv9WyxPCpCdhaX
hwClbKG2SolGcEtI8omwxu6/OVTFK6sLEJ4NNc0IKUajnxaJbf31DzZ9BfhmcKqlx6nAF2RD8K1P
a4UILgVmmkP8bVUz6IXMIlVEDC+t0xCHIt2FgY0SprJW1qYKP4HgfOjRy07cv4N6CAnHv/uEWqdZ
MydPGFuBRlXYM/bWeBr0KtJjtmj2NCupbBob/prdIaWhoSe3UAfQUmdqsKmrTSkNezwHlNJwQKom
mPcbUeVnsdIdn1CGRA4S5Q+L+nd1pZ+SxPg6tyLj1cP/dbCPoS3FjoipnSjoAZSTld20+umJj9ar
/UGdCEt6Jg1UnrvX9T1z48Mi5i6BSFRylSVFCahoQVwLAzAddWqeJwfLv6hcW0HyAvWH86hx6LnQ
JA7haJvsmbmqnE+tcgmJlgbB9exY7q2aRpI21s9gX9FOVoNgmaXGqda7nCBb3kLSkrQ3kMkz1XVf
oUIU+Wp2pOVLnYOBJOEnUQq44ln3tN50ug6Qw+7Vsr2MeSmw+wbDDcT2PZvvCMKd0H/C9MGOFPv9
TJdPd2822ejFdUx/Tn5X6RQvlL7C36ZkehmaBdjixSThWY3jxOWHQDvZ3CTGmPk9ZO22NRhKwJ5u
7T5xvDzt5jOLJ5wKa/GQSZzg9A/SHJ+Ih0016CFxKMsBfDR6AVkfGQg6V3LpXDq1jniq134Pc/N4
SXuEVFeyK003lZImuY0+pJu5mwdILIUYMhpbcJ7gehAD3u+rO5p08GUjByQ5K/8RzP6znU+nMDla
aqDjBGlUltjltPvebtVMdkCemR9VDajUj6zISq/W9H93EUSmvYKHR7Btm/Wz1O71RTmw/oBrDWXt
jmCTzWZjPBSlUIQXHY7IyBThKV88Fq6aYFUgsvDhtLBE7MxMX+76Ate18IP94pouZJGiLu9plgf4
s7VuCiQu6yieLyQbzK6qdV+29FUpKOVw+ZDboUIOX2XnvKYs1Vf2Ia9osN6jCRIc+x5JdPFzVu4c
CAJ5tZdQgPdEWbHLmdCqdty/GyfBaKwsVG57VlFpwpOEwb7I1OEHMUoqtVyMGkErQsGYdLwN5nto
RARvaSDOl6/zdo+UUkIuHEaB8sRziyb+M3lheUvKQ3m9HjzsS/Pbhn1edrXmzTpizpiefYz1tFoL
o3K0wYipcyZQbEKmdboDx2vxJInfzn7Hy7hvI6RJWKKNXjcJ3PK2Udlp9gS8Pyv7WjS1JL6odQXP
XI/fbgCzH3cqTSKygvsoValm4ICGeJzZfNtTm37YmlTFWEeTuridVuD6TiKYQ4s+atujxl7/qlag
C4Lr9LqqTPVae/umH64h+Ghs1ScqioISN5NIfL3yQ0JUIGeeg8GDhif9m/h3J4NzQxmT2pjETiCr
d8BhgfcFGhqDSvhk+tG1AH6uB95roo/IF2aPbXyoGE6OMumPSbdK6Aa17BXYw0GHxKjexzxBDVnW
d0W8M8CUGqNe88fx0PytmpWTA8ZTjvTHYki0L7vmkCrlnkTZQ5IVs7tubNyXu7PebKEnS2RYCfxK
iQ4FLo7TQCWXBJ09bEwMFuAy6H9qFaFs33B9pSkpyf/KRGLWT5SkFjLeU/wvY9meFntFxRbP3mPd
w2G+v6X6axcfX667THx1cE1OD7+/GMzu6GO/yyZap/MO0EInJMlVDYYuEtkco+Y79oofn4ZBbfOq
gjdCVEhhsglxjsJeUHu2UPDCRoBqwF1SAwd+o+43JPOlBb0R40JRCj3dw09rYScX7Fgw4z0sPRv7
4H8uKhjKAdHDtsSctHBOYbKLnG3cF3jERYM+phUm6R535t0GGU2pHCmVN5w9GxPkxZxxDYyDHR9I
3gGWDVBuGR9YNvlYDSM18FXjA5HRpKLzWoYGLvch+2Q/qxeUPxYOgO711Opz3HM9SoP0C7Qnuzpp
f8Fqmvw73MTyyO8V3XfziqfpiAZVotPheo8XhiCfBDJRw6Qv/iD8+rbz/43l2Gk7sHVTmCjDDIqa
uYGHM4/U+q93eP30fmGsVCWTL9eZD0F3IljzDWFPjnNNx4e+GYO3jZT3EeZkWzQbh/feyWyf8Wxa
v4BS00UwToIsR+Fuir2+YSH6SiIgJK8QhCAt5rUM4KfzT6lnSWzzg96rcilA+dpmGF+Oc+zob9JH
IVf7LEUG17GATaB4PMFMGbi3lfMBUzlsNruh9SYbkh948/JQJasi9qeTGLzUmk3nXLOQLTiys3Fh
tmWSX49Ihzw5grDRxFZJtQ1xlRRpeqi+/G8+VJ9IdItpMo082qvY5jOo+V4POYkXsE7fK8y1CCcB
h9oGDZhn20C09wRlkaHg2EzAf+VSmo4qX3AJX7LJXwdzsCgtt1uBGuSjBG9O5i3xSZ4t3K4sbaVS
mtw5wNpzkvz5vD7Qh7ZhQBxIonGTNv8gR0hAoQ/lAZ4h6SUhNeNS1/AYnt8YhSXV2qAvWn23sCZF
oPSuE8NDE9n5LpvdrNr1/0Qc3u0iQCfX7fr2Ns96xXuhVMpenxHObUTgtonRFKKKXwpxfyQHD4ue
M1oOI2J7srjpSbCksFvzaTMvOuIpTX5w8SmHc9DDJntffBaV9Wy+CLDHl08Kzo6eLgCu7mvgyx9z
uHuppAzPLlaYVjX3F4vnLtd32hzBac574ZEeo+IAkoQVVU9vkr55b8Ttl8O3IqrDhisI1YbcSuws
A7QjteiHKC+51zGrPLrmIBKrHL5a7cAECFBvXFuWk6Ow5rfb/iQfspL5RIjwiKWMdoOMJqwdnU/e
Xo/80LjdHLFNl23N18oGNosVkFdod9JQPUNHMCba2c4als8vyWmhqaFw67VPqIOf5OUWldxFq9IB
7ZGMjUtvzYWiBfcythPnayDJsy35g8kMm00f0nUyL8skm4uZqOHlfR6tWXaIFk8z9Eq1omSLTiZi
pm4Ou9j2FwfAGgstIXLt0woPxalasoVQQyf5usef4RVImIpsToXJXwFQp6UenlZ2dabbeKKhl23v
9oixsP/hpUrqbLUCcUlOBzAU1lz4bvZse08slLw9Ne8cRLEMq3iaqaCxH98KNjDs+FWShJyT+ewr
Xlbvn76VZF0UvAOvY03p4UemHEMPy4bmkOBgiu3VXo6yCJ25L9HCV39W1qUz+ckdCEtOVUxDaigZ
U+LvQb1G8kVxw81YSAGN6xfrQsc7PO/3cguWERcU47GI+QrFc2ukR5X8SsdBrelshYwGfP7h3s6f
zWwMSjhIqp5HuThTtch/eD1Gy7WW5wRNSEOIwg3a7VE8XAgMvv8CX2LLWhU6JcelmYlAUBlXlIzD
Ven7Tr/uB5B/TYU0uMMxr1Xxw74BHvbE9FIBVp32s/uRwRRMHTxcVnI5BEyLvR3sTRjAhESOe+R6
AKESewhQqTjsYoT9j0zob5lRb1YDqgIHDBbrd24sZrjcn6Qedpl/nxhFwCySRm45osMiJHJQkoL9
HZ62AYnp3ba3c+Mmq+jKsAtk/NU26CfWsu/BuQLS8bUUk0340TrtIpkAX3MGIkvJR5Ywcxqas1Eu
23/gCdpxje6v6+zCE8fxNNHr63gO4Qn9kK3jYEzRfTWfoAdUHiVkpOw2pIcEc9JruIAzxJQ34ciD
+JKlVvqbtgDK7qh086mnG+R1+LFof6FRaBkmiTUCQjL2vnSYzJ/pMhcoVwsfWdnCSVewYGvw2xAZ
z6rkK7ECB/tckO7FrII/mTAueE3u/D9vdPjhtXPyavlresVi5rfG0l8oiVGEj9LB3rtRPRQBwpwi
ErdVjeH3imNLEj4VosrqIsqWvOoI1b8mFOvgq+3wEMf9lhqFQEJ9JMjAkgYfUzGNrqjHhZpTUCs3
4v89Gw8TzJPOrNx1oU4Mi+fcpf2g8MosSscz+8ZUUBXEzuzyopITNILkVOiHgcFv7k7BkiqAwh5A
qLHjpkq42XGD0hIrORuUYYZdz3U9NOcEaSNHQPkjypMhO5aFSGgZy9+8uqhgAt9MI6uQj6kAxYcf
RCnNr08l4ts540kassq7F+dqRjqnRCATQrPfv4B1mHPbJxYXMyHu4Owvo4FYda3lzUvCXnE71dc5
njEl0AJN1j/+cySlCyR7B5WcR6Qu3BYaO0TFkewDc2qQs4LY8msX19+UVfVHbwaDuSJ902LD32QA
ewf3/nNvUsLFmrLnjdZifFFRD4CBV7WMSgzzttLzds/gnWtHs2VqdDeChj/3LGfs+HWAXUne1bBB
Ud6cs3rZ+wCfdvdXObMT1EJu5/l+W+FQL4AgoIPbSBEMip9ptsme6Gde9XOMQWlfSnIxPZsuYt0s
iT6u2Z7VPfn8PA1eD9ml6/pE57opba0wgA8H6QUTCnPEPWkDZ/BQlDOmyOMp7ECoZ9UbgOn7MIbL
cwOHz4wSDwOl+dya66JHTRQjLY8RCv8RTZGtQWykrDaTGMcl4Q9e+0k1+6hHXeMcBFkW3yosLMrr
gXwmO5u5+am+V8UO0tTGfTuF85zn2paxhr6NZGidDTtjAfEiLIZ+QBwf2EpeORktnYnVdSJBoyzw
bVyDhq0kOQ7u3K9Lv9uL2RXpj9e41wqOtSYqO1OIhXPECLmKr8x8kNVdEdUSrKByR5w4zPMN6Oc1
QMk4OWUhSDbDkZO8MCO2IIuErsLasN8oQTOxg9KnlpC+rcFnO+FZr5tOsfvYp4j0FZXGsTuZQ5Tw
ATjrYo0tCMl7yVygxgS5vSLAIjsrpxRPaVCYXjIq8+5Yd13tOVXts/+b2z/okiJtmR3Go1FqN+oj
YYgrRxxZPO71dso8wUQwMpJSrwKZqBc6JpefhJq2g7NFIOtNtKxgjB1wzBwRYYSjsdydFP0p4yPm
oAw0g6eY6RiTOsvFCdCH2QjbE5crNY6dE5SFQT0iDpBLufIVFyTgPnHqtnOGlD9SmUZyNjzrRW+a
vjXfMDjmXl8uNcoAMJweJYt6FDNyiEnc4ouezfCDzr+bvB0XI/WCeMPptdmndPMYc5WwfB/XKYSt
5c7g/zqj3EmwbqzGLIpT0bVgngQf7LnDU8Dx47quNtmvpawWwEAplsR6EnRF5fRMeWf/5A/P24bk
lEne0jXeNgwLN01xUDJv9EM0SoO73fvhYyxKK5EtOH4aA5e+P3t+Q30HD6f8hM/YGw6dJ3PU++Xy
YoyGahnomSU9yl6SH9QutURayWY5YY4soEcTNLZgOsLsnO4nb6FkQV+yYHx6CRaLu+3xHtEG5P6f
xyZNhV9ASGjhy4SqyEhVIoV/s7w4rG5Ie1K800Wtt+8RxNEl9nCBTDmB72Rq5WEbg1KG/YVT5nGx
HmUlNvO200eewTc9XhCpVRj5SjfrXVjjzp+fyxqf4w6ArBQYT+1MCaQ1q9Q7HG4kx6Pw1b3+tRrt
IwQGsEdDb6fk9ptVqvHG1+3zONiRZMA1fBLppgbMHHlMUGrh1oBefwhghdqDdh9aRRKv9lOTGpgP
n0x4smRvbw5yHia80/idNvdkE44m3rBvfxWdKrARfbIZZjagATEnK9zyPL7dnXCJUZYUm9DrNpOa
t9Ii4+/NocSyCaPCN9mfJOcGKvggSNaW37jvwl3hX5bQluC5qN/zGH/asVfQKDB2Sj7eygojP382
Nz2o1qFOCKaCm+gTxIrbHLyD51Yw1F/5VP0c9fQvSsqeVC7KREChJQuhxEcmSZuk/kUEUIV37Ure
JZJAM2K92exblLK6LvqE5VR3h5utttzfSp2dcEfDw8Y2d6E1Vxv3X1KG7CvA3HQOXjhaGzhYfSLU
8r2OkMAZANqCLnxEmvRUzD2thRVrbJP5WnMz14Rdq/a12byRmE90SGlPHY+xZwj+kKQl8mWxPqeK
aO+0J/FDQrToigq4/XmkhhzZtXmfJagVbYnjJ/JFnCoA9F2NU9/CG8hmOoMDe3zGgzsX6TbZTrQI
Tfd9GMFpERi0Obnrw0qlzjRkYG52eCiQg2DGoxAgxiXVnk9SknSv/0G4mnIOIO9v7UXVD+XSMPTL
mW023izh+qbco+LJO/jWfuY+UawSsMclu/Cbq3FLAfG9aLx+7ub/jlCcgdKhkko9Mru++s6S9EwO
kDXAK0I6sVPzy8nc5t1q+jGtmEbgbhechPjmQ4y+M/C/avUoOtYtq0Cuv8vBGQHNPspILzjDJrJ7
ovCJ6TCPqv8L8dstl09ALFFSQGvQEUrfs/2sa3xcBd/BWi4aWr5hqF72pK/6x8vtScS53TtljLmS
BI4mHeQeNEaIVxm3jhLThywedIWDADyNkaUMo/fYHVR+OvzJVZNW4NXWRxcEzWdw6tRg0yYyr73U
lVk1DMWsKvrnnfkLjfha9t6/dvDoXGwAHbWjudJhD8s5zBLMI9IKgMPYwXPNv6YRRL9mxpSWSHAE
l0McqjbX+enLy2/3h0O8SPEcOTKsFllceCwbofkBVvsQj7NlTCZMiLXk/U3ftIqocDiOMpdtD5eF
FvcnF9hrOVUr4Er9XPndYUFASU8zCCaMbTN7u7VhgocxCB0AI5gWKf53IA8dhMnMWo7rSw29yxv3
wdsVF9FPn/X0Y250BCo4H4qy1S4egWq2MIw+9imdmjWkWSTONkKoHPyyeYnxj2+HIJFM/hs6iPJT
kRzcVRIxc7QIwxR0XBnd/vZAPJWZZVz3yfbA0mB8Yav2MCOYUkxVic/Jq7D2K96El9VzkEZ5YYdi
fNeq2E/2lVzfR4d/aXNcCI1GSjnVSZxw54kMEstOV8azidnPXHunR1E4Vrc8748np56+GvunqCGy
EXTLOxtxLK1vxV9Je8WOw9t6pXEVT0387MUZcu71BD+v/tYdmhkuTc4qAN60AvLcw3r45XuL2mdN
XI9rs4gXfYlS2mwyEYLTw9FK6BjvlB+XicgxrEIhd/bq/sw1I9x5kNs8n7XVnZEdJuIpK5k7UPEc
LK4nngVbwZY6Rl2YaV5lyI6PYK/RDJtexH2b6BSgRCsTlRW41OGHdUP7xFzQQta3bjpkC2UfG5ii
oiYnu4ok090aAPsRL/uAXmNZma5CMtXUrwNRVrKO9OeHKk9FEqGyIb9FMqSRnqJNKCW28sfom0Xi
c0y5dbRLqgcJDS4x9+f0M6qkL40oz+xEY/x3zqomm+XaAt3uszlfxfsG5ei1D71U+uYUiYKfWAyL
G0RmkwzVFc+px+QZId4hUFtpLThyUEh7KgPTBMvm3Z94CoryG7ASv6QI2i6kTr/I/gTCS6BVjKZn
H+pSKqPJAMN19bFh0lXgmnDqjN87uPTeiIh6dHJIX7RhqFYJMCL5M5vDXBsrRGaH+e7X0HRyL512
lV+DPc70Mvh5GQ4bHVYWsEwxFrRy3TMq0uUevtG2BcWFtXZeSU9jaxLUgroqBhU7d66uXCgtmn5m
IXCqu0oIavhS8d3jwc9rp4V79YBVNf9HBolnEL2CNGqKl67hWtiuVhmeefw229Ed6ojY150sUFi7
+E1cyKGlxu8Z7bQQgie9C7f2xr5wTLX+jNF4g8C6KOmiAEGnFyuYsIV3BUaLlscSAE9inBglfxay
vRUzvcA4WU2cxbjjrjLF0FPgg0Q+czYBvNhZhuI05E2u+H9npR7U2sBVbZXGW6g6ZkvthoU8bOkO
3cDNWau0sbrSENzwbNdb9K6sGysxqz7UmEsIxTW0Q1OV5PJnGkPtXufzuSCV/HhMlyhsxA4v4ejK
UleG2wdI/ToC4sehcEsZDGOnUAS+MWpj2cfhqZ1uFDLCDOwaml30dca2mcfvOpLnpRlQClKzSERG
4h5fkVoTyFB+yVLBXeCSsO+0Ji6qNhrfCBz7yOopIjCvunoglMrxPxKS28AMApeSqZvW42XZ0s0c
VyRr/C3sRjYQVK/FZus360rSq3P+Wp5YRETU8a3TZwhDMxjI3BlHYOs5M2PILS099KemmXFNNz1E
EjlJgOTRI3lhEXMSNx4DqcYpI1F8IRI+/sF44d2uPsQXlckaAEnrNblR2MoJmAcSJoWcMhIZ+O74
gnJtdUNAZARMFPCAa+KN5Cxvuq7UHTFJgT1qYREkn25YamroZ31QNHtKyzgV63IHMZ8XeSRB2P1s
4uO+AksloftmOlLxwDjFyf0netd5UhwVFQG4YFYl5iqPOClIOD6Or8wcqfl68A3mTUYROQeJ//yn
G33gCe/x/L6GJspa/ChDNCxbhi9jU2vi5GmmMazWnEZFfQCvJvz5egjih7Doo9os1kJFkwOY6weX
+abkOxMeJXLJ7VYLqD5eLuD0xn2fTBGHxW5D0Sv0WQ6J4tltgMAo9tSBSO0AYX5GNd0mZaS1GrcH
hYMyoPgOLu5jjVhKoq80+x/K/xgdE0j2jsH3/ziEKmyjoQkx1GAeMa0jQ4ZBC6b33R4MBxfKhTU4
EMg53gXSRBqckAHrfZbKjgXE/wvW+/l/MF1sxvXQ9+mVNbVBE9vEnHyF3vU8VVib3vf6POZpKhyH
RteEb16kbarRQc+2zMubKKWT+0kYKgurliVxT0JuoP49PIjCBotl+2zr1obMBr4ZrocJuKSd37a1
LQTmvJqeKBI09PzGyYSexa7blHLt/rqfka2OPC9VkLBRfdo7/NnUG/ESmmwbkYF1lhzaJdLV2TKD
/KJXWaS9trIPgSw8qt5/B2rOSzV4v7satLSrSwAfXz9KKR93T6Rnh4UzpnjZh3ueUSm4QNs2c0rf
XjBViy0I0B992Z3LlNriML0JXIUL+tys1VOHTBBAA111ti/iOa6PrJEJVcPpDBgR/YmHWOFypL5B
L3wFz76J+2SZKF/CAxQG2r2dgRfIwQOiFBXsim3556VcdInuf88YvIiMz6XmZz7Y9MSHidyDjN91
F2Gf8nawNYF92WV0hnFDeiadKx8qHgXQ3FrgdB7PIT5cdwvRmWRcgLwfzwb5avmgpVBBVsml4POm
G8uFadPGqw/7NmwuIt6lVn/Hp/y4AJ1VXN3Qvl1pg2yUHoOjEZt2K3UdG//uA1qlj2K7rgCSIpld
ZYzmbQ57jeqVHhAPEIEBYV48SSaprDyyABsezi+ud1HiSeLOQ1+l0pIMF5LVCTAPpcnTpGrXYfdz
RAKw+N2ETuCEnnFGnHUjXKuo2RW6a09lkp/l2rZqZV8+qqK3yXy/YzcREaCv7f05KqKp4/n7nPU/
Oo3k/ZujHbe5vGTfVMsPGHCcODyA0OqoWNr/apgaK2N7V5B5PKcdKuJpoeIUutMB5o2ASn87Sadk
Ya122tBOIZjH2PjpBQOMdO37ZKYGSmA0jlQusXkF50WtxiEiLiX5z2uifyRKf9VL4YDkmVBa2nC9
70wdDAPi8QGDEeosIp0yWT/EslP9U9nibdu9+4H95DYhLjnh1IJ5HMiwQy9hgE2YuDt6kByGKHPz
tAUHyDHy9Q4TT0KlmtlTFbvs9dn6ojGjfLV0hQ3n1Awlywxk1h+cZ34ikz1thZmg3O8lPXflKAne
+r5eFVkQpWWaHHns+BjW/dEl7YV1z4xHDr8VLFaWfAvG2uacIJARxFDCbDsQv8+x+lCrhXVBGIBf
IGoLpE3Keqxe97eqZ95R2PacejEyCm0zQvD0UGGXEfb3lWoHsDp8ncPJMGCh1N9k0QX/8ePuQUVB
OgvV4nEmEsuvxP9iVnFQJbD0HaAB521Y/ieuvZDV7tvn5xT2LBe6g2BQzK1xsTHK/fojsYke3qGa
l1C9bqDxFtckVc4PUDSVdAu+/6K+c/M3T5vtJrTvzyLWCZbd29lNyQINYbY3KpLb7C75I3ScM33A
DIwSW4jYk8sAjKFBkHHObfyeiLTwSJHfBdojTMwN5+8bShPZ+A7NOiDWhrkuhf9OQwGkOemZMtqv
gpgddNFK4CwHSJ+MCcZNCKL8F6F55eJu+9NzZ1A3KKDhc6OBu/Ap3LvkvjXCRgvjQpIZ7QrmhWmI
6P+m+MG5sZJXm3ZGbJ81D42dBRA9ryET9RSQLolqrtMsuU3EZgiDAk1U9rS4TILC9HvihsViV8XK
tMoimXV6AaxS6yemkFLfMDfY7qSSgKW/Z5B3X+qxau49yw7QrE2D+7RGJHzGFppz+bRJKNVirEkF
XDT46ilbYR/5kmOS7MOhbGbDF+i0RJn/59JqMjR9i/gHrj20ODpFT6U46K7vP6V0ePrGQqh6HMmE
V8JghHulav/VoGD4NS0i6B+iiQrqB/QY+EzaMRlVKCWhOinc1lgM3I0ixkVSH4nWPv9k1Y5UtX5w
Zlh/h0JPVOIp+CaqYX7WRUKnkP4vYGeguSMUbuYhM4z/VqmS8Gaol6kC+jaS3d27XLJ/rALd4/9/
pm4hHQiChU7RQf3ZKfayBm6ABWGO0rnqYoqfMiz5kUqtBJ7guXokP7aSuKim4y6GHAI/EFNW0QN6
219ehfrMObZhkhnzT6EjBWwH5/KL1KmyX6qFWK3GD/pBCx+Gvtq17OzFjanYV0/fgq+YogsXmvTX
aBfdmrvy/+hsLOUIBDCwvoOOgsxTQjZEBdqJCEwfEnvMGIvvvyV0P2BNQfs4SgY8r0kiri0cnTJT
d4E10ChAPysXc8St09rlT4PAlY18l/cY4P4XQIXqt0xctT90OZj0VJXJ5t8tffjCIix/JpND6Ukv
Ematc90bJP/xdIywhSlX8PgfXQPLcU1AYJk/cABKEuwXc6QXDs5HreUO8kmcX5yUuPba1OnCaq0Z
2XgkXK9n0A==
`protect end_protected
