`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pGwerY+4jWeIK32CA8RJTzg0ff3v+lGMdFo1SQEBMvXlUhs0TPuY6xvzazHlu2yvHFp2ifNJagZl
soa2ri86lA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
tjVma0VaFkbJwSJ/m0Wzr19tHIn7eCfqK1VRGDVC9lPuCeoMaZgnURFueO2rmAM7OiglEMaDj/2f
AK0GL1gmADgmmBbVZ/y860anUHzt+2gpIbqlwDR2H73OnZ2TlbDn1NbX3BWQ/aZB9CX4feZP+QGW
9/DwL0/tTW+jAH92bmM=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jab3FtEs6CbsbpFGkaGl/5ayuSTDn27LVhXEkSgRFQJQPcWpbNlPeMWMxv00vgLIch+GbR4/ri4R
F9J8xnKG2qRgkjNC3s4Uk/GoF8jNx1Vbk4lVwRZX6OQl+XpwR4WpVLcVd3Ra3hfHk6C+sGx42XaS
X+afsBmjsyw+98kCrDe92Hu2x+nHdoRnUyuFBFLlNLWdiFAjWthaOZC0Ot5ZWbvBE8BL9X7sXOte
MRw8jx3qhYhVIlVNpK0Te6x94iWoRRCRfbPtXzTzPgOfHcCWD5dNRlYkCeIM5LzR+S/L6rDnYN6g
tQz3AZYSC/N3BFK90J1bkSvnNWiJYBxanak69A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
K156ee21ACRM3cnAZM+OoGckuo6PbB+qlYSeze55LxNFLqCm3twSKLRvj6eBFFAZN8JXCSB/pOe5
Il6Ggo9zzBFUqJeH7O2GZmQSdsETNZmHh0YUl4HgTaubkIHpeu4jqvgqN6YMMUlD2/t3LYmQEzxw
6NV0z8AhohQQQAhSoqaocNZ5DmxjpTOe2ypkYqPATbQQqLmF2XCfaxSgPArmS3KoAYgpy/I6K27t
ojXXrV5a12f/I4+5nB8//y5iWvEsaNANN0vcVRiVzrWWFncblvxJBrqYuAwq76obebGJhzlVsxNe
nctRtjkfsBedhb6tWkXFuNpJQ2CG4/Ru/gTLcA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
VmS1TLOdl9eDuO6JJzp6RqpgNvoErDF8jKy/GnL/QeR+4K/xLN86hyWKrXFUpnUH598Ss9wiHew0
1BdHT0eqeuQ+LC4ODWj8FYRm5pQwboHqWMW7syXnZPP1hiSqlRp9KU7AQLS1uiVezki2YgWyS8Cb
bCPJznwwxhMzdvu01zU7hBnCXNjsAThw18yIcASxJxl6huVCLmdQxv8e69SEAVZyA19DWTL+Wavw
RraSG/4jqiSh7KDYCPMscNVKYkkSmpXkmrhkuNjT1kQvib3ZKqjtSZTXDJ313l5F4yLrQgPO1ZIZ
pCjWfHz6jb2uRH2LKrjz5qWn/6aXa24w2LSYNg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jOPxpiQQbt+/CMujsiO6R2VIzi8AIpb2xAYfGC55edCmbtT+VM7LbWCAHq2IIH2HFGeo3lClOVoS
HdamXZ2Ggc4JMvQRCqxSG+mMfBA3j+lLR792HxpZv+eH14Qc3ERaGN0DvMVAiM80cHUzNUIaClxo
no9gMOKu6Np4aIRnXLw=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
o/8FbYwRHnmZ2YAdx5IcS0DA+j/aCtr6Y6zkfZCNibemLmlRmtxbNZ7EqnwpqJDromwIqhznBAt3
/lzRvHnnLmrVmjtyeyMRvDP/GhS3kYEg3ZazXlcemtECeLACzKPRCGsZdpQ2w0iZ1/KKfAtroBs3
0WYBp1G+O0qgKTlG7MtPCSd8Dd3PSecHLdu6ZQgVrvbiBYdkLrIYsUbYZOMNBL0Y5A48G2PiwCCL
WQaR3RJP6b8HZul79+Z3lvw485DLH9VDr0Kv+vgKUCoFCq0Cz3muReorFhkQq6Wv1P7IFfCY2n/L
zbxL+WyfuAsRlELMZOIZg9w8wAv7bMnIEdVVcg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 566368)
`protect data_block
JxHO+dL+MQW4a9PlXIp4IOn+oyYQuZND81qClZMXvxlCoU8eKTAcuYKyGfMLVzzXj1z0DqyLTKUr
wU64Yfcz8zZXaQ9dJ9v92WUf4iLdiMpDRQpAOyrB8pFtCymdrFbJ1szOVgXoBR0v3xxF0xqywBz3
coy2HFvf0NT7JJC1mrRhEbUR5xsDPiCY4R5dpvaRH43+C0m1dc+S5rZX+TPmadW1m+t8LLim8Apb
fXRza43m7ylji7j65Y7ll4EPe7ADBBr/tagW2tBPzZInDnxopo/ug9wlDFU8WhutPwUbMGFj8ZIO
nu12plbm+cNro4mitZINd1+9NxzEwS5RKUqfrRmgGQpxE2kpBEYwtx133PC3rm0LAqTd/egQ9t3R
cy2lOwnyIZGgkRjYUhBH6rnLY6kyOrEYj0MPR5B81PPnMJwmijgEvPrbBnzlEYiLsrKP0xx1nOuc
D4Y2tePrKZyV63yrHp9PwOho06A+vYWyD+O585cKUqEzS5phW+mdGH2/8mOZKSFKKUXBmMFw/K0T
V4UMuxVi/hwrvuEURYbti6NpI/Aafoh69363zAn/1JxghBVHJcHsimerXM/AAYi+jSvr9S1rjIqH
MNHHJhVqCDpVv2NEYUA7LlS2PxZ5eGeEP2CnWFn7iQGSsod41MzLyO65x8XlR9l7hMmh0d7XSJ7u
08NhLFaIa654bHImC8YqSZ96JooZVLP8chkpCtB4/Swctm2zvwzmy1MLFFpsZ1CiD3dELWB/Tb2F
/3jgx7gC5Du/Z51OO0W836eSVNBoz0oXUMFpxhiNbgwABbcoSHP03a4dkIJkXVzSdlDw3W8/JCK1
gXVgcyhyIFxFTRsOz/OR4rBilVXFRzDbON6y0uNcelpssXgxew3PlA8r6DUDg7ClFb4JPiOpxErZ
GNqtOtrVwc7aVnRJTdPMC5O5l9oKVfQSrEOu/uf016Sgnv0KMIcuV2OugqN6C2f2dwXodkggS0CZ
wV1qwa4UTcpH/wr0buwsQGQqoVnWNk0fC6fWQD+cqZ8UgqlAOku+MktZHeiLlvSghKz9QzqUuTnS
ctUTFzAm7BN91QRVtWg+GPX5A5AEGV4o2b9vSKLdOD7Zajio3u/2mQPvV9vXMm4FPw4Gm3qEEZOH
lK71a4g1uJPvVz4M3iQc0+Dbcf5ToPSRZLd5NlrM1sJXOj1ApghrYUw6RoUr95AkKBgmNkgXI0GI
1AR9vqm5CN7No7ZYq5U3LlQz1azYgGmqP07h0I8g7vr6r1qJu4YGDOB/2H+txIn94NCLSzwH6l5W
fJHffTTzmO0qrUJsstoFIvUuRdYrABBMRcLIlI7WWimOsCPF+5zmbnspNLylU2a3U3qYJkNsB5A3
gHqG4u5Bb2bzUTP/TXqvxzRRla/KwRB6YX8fRjmFz4nvSGJZmlNVz4aFKzU4dxKNY7/6mzFFc9zm
6IawoKctH3xmiCtTO+FZZ4c54EDLzGqqP8aPTWr15V244CBnBwlvWKQfxwZ00KWBquW8OqoK8UPI
IKIjWoNDxBtXX72g01s1xz6BUihGs5+tD3EjOQ9y8BcZhOSUIxH117iGchOZBUCQbYKbszEromqS
xibsK5CUP/bGdX8R035MBQSQpLfFMAIWo9JKJrdZ22iEnXadK8z4q4jEOtSLUy2RhRtiwZfiCdKj
gPkPPYW30ZmrHDZ3jcLqTJvbyAs4L7iXlpLZrWaNnuRzUmbd7wtImkFzLe5K1WjgvJaxeJa2JM5J
cPCPB3TcjeY/7dX4bUokuOOTsBOE72X8YMO4b66DJfoik6XTFRcenfYFHnyJtU9DjhU4zAN9XgoX
+YwEIeRQZ5nndovRrj8i1yyQhF9vZwCxT0kt0IsYNRjbci8dZZDZ7Qy0jLQyGRQmuCnAjlKSL/nZ
9PzrpkLY6/hLBmRLflWpbMrrw1wtDayw+Q5LGEA8CX//LhmqH73JxK9KJLkwiGEXf3D2s2g+8JQz
L3IQZyPVsOnOqxvq/L9oFUWizUCr5Q2mtqlwWlSddHluCaRRx1uZrZyxhLv099wWIef4dWP/O57N
U+SZrlpO0BZ7sdVHEQRNhwFNj6ycZNXEYH8ama+/m51ATO/FnBaBe6u6cuthg8K/KifXvsRcc/11
a9vqoeNNB8mi/zTM5esy9s4NOlDrHYUJrMoL9ZREK5hXFiCdNcmtaEN3HfzHAIcB2E9Z6/GBpB1r
8vBdLqzpXoR1q/T8YCHzXBC/6nRfhlhRGxULuTyPtcAER1rTZHHajOcEfM7BhYd0C4FROCzCNznh
A066rSzt1wu9DitppTatUz7zsdGOiQ3naUpyvXnATfk3BvdBdI9IHU9Dd4YD/cE9ot94YQTD74DG
x+/VRcWabzamnI7+LxyO2q2CQ/8FBH5LvGc6Nur/tUBokOkJs1+w1+CLflO74Ta53ZRoaJ/RXg/y
siLPQyDYh4wMJbDCIgwGpnFrD8pW7bMu61llBGor6BuidWqIho8mXS2UO/u7hgvXXiB2/XDOrf8O
ADd/IJ7QzGLCo/2yShJfkU//g4/aWbBMTNYkhfUqntLloCBhIOdFtYqMqS23nRUO4GB8w6Ko6qja
43o/G+3cS0hA1HiAirDiFcOks1NsNTWJ0kn24i2ZvzTdFsVahqAivYsxJIAFxDGqRKZtg5ytZS01
sQ5bmaTLxltx39u/TEsa2GbJvP846GXFgx26K7XssXAzIm5EKG7MyQuieEELrml5OOXUZSnKMnIH
kjhp03pUWnRzsbZUBHoeCs9s/Hoo9H7cnjA6RHhB+2UhV6Hg83KjK4cPuAWwzcZveviojDszuyUj
X78gmiQlKBvfJmtUwol62UrBAazD7euvEuU3CFldkewn7rR+LSqq10oUJK7jAYMtIht0imwrRtLo
6goL1gmfZuouwraNkINu+r+J7RtJ/p5L1Sw5byIB5hZi5zldWb7rFHbRo+pX1tL7pl/qoe7wk7Nx
EpPiDjHwd7RXZNnxwMN4syoKNzA0n/jLHIEx+sW23kf4SkKkJCePsjWafp1XQyRiUhPvCrc/dpSn
9xyiXAX8PFCJqqcRHBXqvVFIEgJD00oaJi0436rWAXIeF3DZdum8v6K8SJinntFVGwWbaMGk7LRG
AmdJRl+kschHvLFkldV5SynvDFXZ33qHlRSLNgEJMOs8+JzpH+sAo93i+tU87Q3SbmOa+Ol0OjOa
Y/vgWcUMh2g+NsEuFVBTohFz0oA6DteYUIH2iXoa3SxKbgF+Q5PCUy/twTAs7Tr+4KhF6a1gOr8K
BdkjeNShBoVUnX2jXKJnfIaCRH1rc1XXor2zcx0RchtVUC3BB4H5Mx3Xp8uI+wc2gY2tuhR1r/GE
x4vghL6UGFTS/Y0HFSdkSF9g/yIlbCsxol+tpWgtc3HtA/RGsxdy9qW0CMFZ6/COoqBkuCridTl8
k2Uqwfqw5DtslUu/fdY+m/CjHaH1f3ty7BzzTD1yurCMeqX7YaxeYZ2L+owtGO99EnICmjZHzurC
EbXGK12FUtbaaiRmFfwFWa+89MWDcsdCXxiYP+DnbXJ+3CeXJdOZgr1XyKb9mAwMqRvOXMqXwqMP
KbGnJLwrPqj4rzyz8cOa4pOEmVUYZ0fO+k6qt+OzpZVeu6lyyVDE9EJw6FLc5zY8kaJ4kg5NaUk4
6OnBlbfHTjoWkHHD+aoevRNa4sMQwe945JfInhMMY/RW6iokIY1Yx5e6p/ceKszZBsutvY4rVYFM
jdGlmaYCLitS805S0bPySgJx9VADzUayXpqCcrB/O5hdPg1wMxXhQP912U6GcB7QVM4thYtdqDJY
j/NsgNoz9s7iHMqeZYXG+COf3EvZ+bxtyxxl8DhSIHMgv7e3U7mBXgob8FQKggrqyfuvKpIHQYat
vmXM/34ixr4Iew+7wdHFAsg/MIox1A9VfSDIjim33Thgcgi1dElNZVlt4GZI8eE0rjDUr6I6Hgxk
Mk/ol6YpU04/EZu8hFVtQswjuRXUEGA0MKRnhsFmueckQMB/nHSj24s+L60JE5zgOizbUKSMV2Jf
v4hZRCeYpZXgVw1FM37Oi8GfmtXdd/Y0d7Ol/qKOIW3D1klSqYSrQHJIMlBfYTdoKV2ZfjnGD2ff
01VGPr8t2yK/bsAecvU3xldXG5g69tD2WpylrlOAjRB1E0sAB2cNCAam4Pqg8qZrCSGj/OvaoSvA
dJR7cH+LNSnrktbvGb2R/GItF/eUZaYZHf7im4T5ektyUdxkmo/yWTqgg2hQvvcJxvies+Wu52J3
d2IVeoQZz9HAhlH7glk2U4mQT5tSSMfAE0QkymLPzIOXjrdfLnqbfg6tVPhmFYCwxrXUOlZYdrOl
s94ic2bsy6JMXqyEX3/jUmXkGs7t1wBiJ1vQUa1mmbdyeZLBQAS8UNvmNgAsMmcM2Qq75h3nOvtC
X+oC5CT8teBhz03JnXG1sxvnIU6ViPu6FnpuBaPxjqQ8d0FRm1dWbHa76XmQYErZBdsWFA/2FYNu
T3GaFvWTiKGEMGsiZOSbueu+EdPPkSU4pimwBeO76J3V4J64gtw2i/RpsE/jafB9w8tEzwth+C8i
U27jdJPJ5VDPpQE99txrcadxJ/9mWICLlyfDhBB74F35ccG7RqrmrYfnHrDusxFwyFSPmSVni6FQ
0PlavyVeyK9fRbRE/6cnJQlX75Y5A3GP443OwOGaE7yCR6r3A7hoZxLb2s0u/RB/oEso5jJjvbYM
E9OPQ5JNk6s8Xa9DVVuJRfY7Y8vGSkxJpP9KqT2KIQc7FZ4/A07nWdAvQXDIf8lhNlPmC9xL0umY
/+I/vHyJQvACZmj27PHgvUnnf9reCZ1wqX03nr2V6klaPQvPG7E3I2fwGArFKp1caVN1hfRCn0D2
txs4gz0hLfkQiYqZaMrLXXa5bcbqEU35Wzpn8VPQMMgc7Xmu3Xz4FF0L5UG4GM7Vm8bypV4n8opI
dR20mhUrYF7BnEmwpkNo1nCxp3O4ug7kVTTz6zFbiFVScqQEwxznwMXXwkfcmREiPPbd4ZyXRuyg
VbDblZgEU3LzNyLQffe3Ox0GWGrC6XKAW+pCdEIJzUm0G9q6Hm5EgMZp8ZKHkxb1eOwi2irmeG0o
fMHBh7Hb+NgLL5xdJ/N4s0O4pBxGacfMhN/vGsRhSbPE9xBuSNvcga9eptK9OH+CT622WhJb87lN
owI5/CPphSv6WsvJp0/07P1/FMv/gB2DeNlg9IZuhqqbVP3TaJXre11GqT/9q/0BpRiS8d9/vY0o
TTwKDbCyi2Qgmxm1AmmGcAQqDdNzWIh4DxKlxGIOo5AYE8nudSR1q5GTg1lQHcjM3Fyu6rvmoXUr
bDMosSKYbBLcwKvdM8pMjZBZi13gWVmS07Btje9/ok7rSwbx4YwQ4p/ndGPxBJwW7AZlebKhTS/F
r3IsoQIXvuE0i06dN3HhGrNwdOeMhlEqUXubhM79dUG4B5Znj2eQD2yZ50DwJIuxCKB5gd7uNy8p
Up/cdxWgNrHKM2l6UFInEfZW+ZJGSzBWqvAul6xnWdQLf6GK7Xpnu3ryrV+I8HxpUdu6XCE4tc0n
/AfsYxPLVh5kwhil4s1WNcGaF0QhMgXGz079gJZbLtOLu5pULMSVGpB+8RovO1hihnMYqHsSQc2f
iDDnCnWXeK5GOJso28qjtABYSaocPInlz+DTXIMy5dLhANBFPhNuub+jIqxhRq9Q2Pm8CeJwLZ6O
gga7t5fI+apYWWmnC3FTr94rw2D5Wd8AffyxPy0+MVloGcj92oRg2qc3/7Y4ZoiEbIGPn8UnQ0RI
r49/5+K8oE5/K/DCOJ6RW2OrKba8E2uLzUvgiecUjyd7rR7NzmoGbtasKkWws8zSmSvQhqaEZKwT
LmayS0jMVqtlg8TJBWFt7kT5SdmNJ4lEy+Wbgrg6+1GN0rEA4+iOW4YKOj1Lk+dTgC62H3VXG9oc
gEUBJOUNSd1Gmp25/15UWjaN+Fy3r7bEL9mXrBH7lacrATNyG6I69qJdpEnSJuJg35v0oL/KIure
NMb8F/Ep9DFbswXoL2oc7gNUmXokV40ixUCV15Ttpi/LP0Tw53vf9msibSezUJJCCotvK3tQWBpb
ybm4oby/WqQozVSBlpf9PmSb9IHjHyz4msoa6vtsa9m/D+GtK1gvSwPtbrYkxWy8WQXJpVfizeKp
MFD52Wxw9He26OLOHx1xI9vOSrNJrEOAfsPyuDSdGCIFYhz3HLKHdBhkU74YnFrFI+7oIMvGhFMg
mepfeh34soRdFZzC+N+7jTf4pPA1/HjDouus5cQARBeA8IEpghevk8NeQY1z8fo9HhfwuaHAcb2x
4E4uNJEnDsdXzhkVNUwI3PT+zW7hVCFbWvFqoI4WGH/WQI9OHiUjypr5qnzJS8WkA1Zqm8Mo44k3
RaLb0B8oZIfhizdOAebWj1spQnmpVYBnfG8Cq66pbZilwccghRJSpVCb8uNue3Trwzfgyea6KDHk
1Z1YUJ4KAGL+cM20eCgnPSxkvgCSiaHaklW2LJ1H5xTeoU40jfYy71sOrGbDYl0vxbhYXUTZvBgB
FGWvEwx/aGMB7V1NouTZj++Ffg5jxOf5JzzFW6VFfP1bxA1XcK+ylI0C60RipPmAta8KzMsSmHYN
C1GfWihhJ5Y6yfoH2Z+i8h3lsv4MVYvaazBdhM2IlBQ8XZtZb0piNamS2vgrhI445BFMkzOzjA5O
+JMQforUJm5AdVc6d+IAepSSyRjU4HyjqcQG/rdt+KkhE1jhTEIAifRBERjJWTyplxzKoztPJ43g
RQUdvbHZaSfKyPi7/6oDLi6xW60+fAzH+vrgwFDlcyztuM2N6wRbERiMXdpNY6qxJ9Ob7kz8cZ4D
rlhoOwYZBSnoozR0oBiEGOKUWQ/Md1pvhkQINr8hatrUDFrXP8PgshnBKbK1s7Gln6UA8GzEmNqQ
4hF1jCww2ZJBV4ETTJnpjjHDZEIDw3yZoDjDm/k6Ma6/wiW9IHurm82ihf8X++N0aaBHIHdeHCsQ
zZyJoIUu60o4Evb8Y6Fixm40JEzK3yethXSnQIgP8Nq74RS8XOLJ2qA/PCyoAlJI9DFQlvdH1HA1
P8eGtxgB/9O/GdOo5AzZnKF47xnZ9P9aEASSLvPepaSVPrGg6+iEZ/OrYxVOeSrBA77y2adwPZbW
5JSHpKBSolXiP4l78da1QG743HgcarUg68wnDGpPfREkSyiRC6/RthEqY9tm5AVsXgG7xxe7ojV7
CCWTL6rwBnCHonVSc8RhqbH5+eXDToKoh/2cAneHNrglQGGsqNK52c/bI7GJ6zdd4SPqN4g/PxS0
PqC95Bp1jvEKLaCpem4eIEZQ5awZb/PLKtTTUuocFMDgyYL9+cOIcZ2FrxlVXYWROJgPIVDKKCoE
tfT9wx22FgIuXi4uw3yrTWTow4QJCjeNlpbFtMr/mw85rl5/dxWzzmQph8/7bwtmKAxmOkJQRL6K
Ybj5SM9lHQ3Ibjps7Gb0Ry41dqFRXptpJBF3IlLlWoadh7HBF+CiEFKZ3Yb0dIUOkVpwcn0qN4Jk
dZgFvF2qs++V+8GM2+Ugh5sD09fBg9KFac+JDwmhm17j2oyIEmKg7R04/Vq9EfFqCxfugE86OEK3
Iee0N+VLGMoqw8E5re1GbQCXrTWgX5WunYYksgslflOMnN/VjK0d1tOilyWlCgyiUCE2TxcW/d8K
TTYV+aZLn6/DLG92RZxtP3iHIx5nysYgVe45ZmH1f+aJQWFVKFm8ahj15AoiiM7FK/BSIDfe6w4y
UK+5zDuPznWF76xm3sinL3Pj8LsGsj95AXlGFekQ9MPL5lRZF9cyYKrCoI9zbcC509oCvaoMCU0h
VBE5FpGgAnQzYJoqP9rZwZbm6HoPdH+wWjnOW6rgJjch+fkKnNjpA3HVy+ugJWKrK/M/SLDKKwjt
m+ied5/uz72AWHQG3seG3qqVfLUgudTP964X0h1hSjE2UNuKYtgjvbQ1PKr9nsVCxCnuJjcwHvhq
xS3TlKn4k6qsD2WS2oeGq59jJxrezBYYgL7i0Fs1BPf6/rAvjXX5Jal8InY3fyRS98s6Yr+5PvAY
6qQ7fohUpZjOU4KddRPNTbPDdLs92vTsHdj/wCjJh2K/8AIQ0/CuXgdQVxJLsktjdej1u2KsVH2+
Sf/hiDssEEWaUwqAKqKjhMGI9ITNKnibzvHLSQseyZjOgUyscAjWIMcB/sI4OvUOV65Dv9oijRX+
3zjkpud9xjKmRXNvnXCE4eRT9uaYjwZU2vI+/Pr58B31GzkHOgYUic/KPtVmGHw9EtZKv3BZIPTH
kaz8hmagn1yNLVW93KspXTgcEsie7lzZPLanWGivKb5IsZRjSi0SBB6e2XdboPGH5bDmvqK3ojMp
G1zeVc6hxJYleXXD01Xhy0kPi96t04bxkpIjXRc3u7JKKPVXSg7hBhar/XwFyXsERKrGTRLxi6Rj
llG4RBALun2ioqVmPuf9CRDTgFQabRqoXuNDzU6AqwdQd6nIOX3UPbSs1m4YJk8NpW/Rzp6G/maL
Y3Bg0G1cUvYKS+iwl0si+uCR1KnbVpx943c4Io31kv9DCiyCbyLl/W9EMBKd86oENydWvHOFCjE5
7OcoMdmBnFr/WvPSzvK0ARc2hOz4FqsbeutOWkgcFiCnP+H1zlph8AzNRkcjMfzLWRJAwGp6ombY
BE51En8bo4kziB6VjN92CwlfEj8TvfZlS7YXQjv1Ziy1/VLNpEMFPVPCLUktXK5q+IxrfTX2Dm9b
LDzbMStVqeqLqP94/4QYly+I2vn5ENUGnbHAYgWbgrFx+x0MLXJn2QQ2pWAzN/DhbGuFE3IVb/rH
HizhkSQkXnz5GnuUlYFvOXZQfww0o/JB06+rhaR9HLIManbhe5Ga3kgTW1JRjjaaa0SvSJYeDzJ5
xUwS0hoCBArSh57lOmVuPH5CyMup7zAvgVwr418h/YRxocSjlXuoPuwGZdxJ6Ij4AR1URdiA0B3y
JqRImDixqFlXuN9wY0UQXnKIxUGMKp7nL7P/Pyw4m4DoaStsulF0ZgRaZs3nZ3wpYYOXZxd7Cd53
SNS4VU5bFcMiMbdRq24mo+Y64HhaFW/Ygt6V9eBr8OurdC06VAibAQQj25i+Ul/ThTsiDpD8wN0g
/daAscSE9KG4niPbuYYTTtSgZ4tU9ADxk5OkL4xttH67GdxNRLop/1pREQRO749hBeoZIitBKWR4
/rOSIj86P96DgYA4pSFUZytDMDo6MWBxRjukDlLIak0vyHgbHYQRsnMoQtAJHO7cXuNXGta9hRfz
A7+jwW72lAUoE/n1/RWG97ONZgKUBBIPps7fWHmrSVhfN/LDledb+CvKOzWN74z77+o5CBCFhGkk
SrSBu9DkLeiqZtuYzulNfw+WDIjRu3cgyc6yH7mW8RcDcjdvxitlD+bqx4NI+AAsxO3M2+DLldbE
eSHuicrCEGML5VLGAL0ronKIAJ7Dhvy6Wzplvo/YWTSgGn8cY+RyLq0m6uvvkooMu7UGbBuLeOjA
7hA9I9/qgb4XbXFFN4prhPK0+OZ1Pm/2Oa9ZZt3Zxpp1WU6JitNIOBHC76xOs0Nn/LGPbwoRq5uj
e7KB7Qd94M3/8Qw9ix7VgxAtu1LoPnYDuHHSHGPuTO3f6a86W345DzzSgwHmQ869uB8weNOFdGrm
6sGYBfvHn21s5EMu0DbXOGMv274EP5sxy86E9AqyPQFdY9x0xY3MyDS7vyENwge8UX/ORSx7BArn
8BWUWHdEFhg9vZkbIHWPOGLFgGELKiuza/zfAUKpxIvpIYolWuqSChc5+j1ywf6tIRVPUyUXSsIw
LEMYsLQwrDyOcIF4RwQd3XSDIZ1bpe5uW6UNnVRkQPqCW+HYfGT8kDr+S5ltFxIaLbvVt+TodAzB
4rg9iHadr5fOLMVoKVF79xUeeh0wxcilWsm3Ror4C8u+mA1oOMtTi9/GTTpzMd3Zpm7HCyRPtE8Q
lisVMW75wu32SJf7J9lO0QPZMEYm8RJweIykmmTP+s+K5g63zJ1NbP8vnk/RQNEawYfc8IBregBG
ruQTt62pEfwx7YSJQcNrOVQOA5KPW2v0QzQb3pbRveehyhUd87mQ8y7V9Go8N3XRpB3AVrzDySyh
5NVj8+l0FA80r8X/WqlUEy8LXUuJqFrLaN6DpZwx2QAoH4hHfYX3YcVnQKAtxP7uvZRkxlY05c/A
cnHaTJLNU+1vjEB7l7b5MYk0nXVzHcuH9VClijYYaCbeIumIPQcyBTkBk0KdrFWNJkdWEK1VPKLJ
5hVOeJzC2Fh4td23+I41wlnrXV2BzStX+mcasjHo0oRmAqJ9WTZdrg7ovcr/0Ah2YRxC5TGgEoui
dpVuY+C0NyTESPcm6TbJHEnRifabNFexTPMlkNTbOcOZs3EAewq9tIhFGOU6gaDaBeTnBzj7Jr/A
O9LN+xK8sDKG2qa+Aq0DyPTxf2LnR7Pts55bIlhpYKA+T1qDDQHAhEPj4liLN57SY1BUMrlWFwNk
peP2qrXml4xOsQ1vMdgAtYqpTk9Wh4vHxb/gl5aDu5y/wa6Zz7Q1WggLHjQ/z04CSPrQ7peo1p2L
6fbPBAeQcmgpUE/jbHE+84mDPFOhvWCULbobKQQhLJOe4H3Q1qIg+LVdIR88svnDtBsOf2mpsU1A
b1XpLglFfz0lk+2H4JlmedSFjuNNrl4MS/9SlKV+lLaJhJB/dGQCxiA2IIQl7uWylYUKgqZLote1
yKPDA7oGYtCrE13MI0xgctbzO4QhxxTmpaBJk+k3UVoSTzdKbyndElvYjcHoE/io+4zlsRuqLHfE
ODdCtE8SkyZLX9Iaw/yhXO4zg9GztKSuc7Vw3sfFBqUDa8N9Sv5V0+SswG7t3wF5B26ahocwI6t+
qtWCb8kIwhTRuF4tsA2PErtFEc2318GwsGIXhIe50aoge0SnO5DLNGOD3RPXnhAQlpTTW6/xhJFG
CbWfuKr1H5clX20TrAbqpGm9tlLFowjdZ+QvshDZ/RzXUxMurpiIKmhzV4mrgox1zmW6HwIRX/Oq
PSwXGMpsHW9DAJGidNyWzes8Ep5N15a0YLiRdhp2ELZGDb5TAvFd17Wy/DpDihWx2hnDzBIiPV7L
BvM4n1pjzenTr4bm4KUCfC5bBcVnQuwHCJaK9KJ5sgphJJC8TIdvuvTnMfPOphNRJwKvTvmmblB2
W0ijjz19FwrPtP2pyj1JmwJbi8EABYNtqW8w2wDrWZvD+vli2ptV+ATgUaJF2JCpyk7qqBZg1QFR
Sv7Ubw0OvEBZrMeR9qkQVMQqjhWfkgKh+gL2C2h4atfUdK5bTkXq7hpCr/4RMWplcoBP7LlQ0tGN
6JsmnClRqVaEv4BK5mQhd6qM13MsWOnNXpiLrbA9NGkh+GaSHsOwlAb0M3dsCY6K1ESLN4bPUzw0
8FcY2gyvDAJQq+WVJrbzzjwQt4zFCwRlakHMxmhXkpVptr014i1ASuGTHkcvSZezIwChhPQoBbWg
lmoX/0rCACJpHLpUFeelW1axqRJdVwqP+5uBX8PCwZ5ulFz2nA7tIhkzk4dpYsjpD5+iwVkKnEJX
OPlywbwTP4iaGMx2q0D+21b7Wk9UZ2t/9Vdz/TV3/IdYS+RnjCArBy4MrKwC10JlKD4z+WjapkML
lTFaOSOulOGtOTgI2w9nt831JWDrKBz7MA0v1e6zeqix5bjiOEB25GR+0tJPQ6q+45wQ+x5WYGB1
Sg74hjMrY40oWlJ9eb+JAkjSHpCoQVK98g7wBCa1h6zpKuyeSCmngcAAIqotNa0Cfnb+wfVi566m
unfY9TXoSYpYyiZ0fjotRLcTRcuU39dP5zvq34d4PppsAJSpTYo+Fon+W1DEVzKSd6+8n9CF2cvq
KUQ5F/+yEhlhBOPJc2zIiU15/s3n6tKx1XhTRtuHkhIVdWbzAYdkQFVsnPmSBJ1bSCCBIkBCA5Jg
+ie+i6tkTyx390whXcj7Pve3lZYS58C25BPHJrDUZlcCCBXEKLckVj7E1heFyUX71H8pGlNQ2wCw
oj0lZElSkQyeHMsuM/J7tO1g2s+jVCgkfkaZ/uagQjcrEBNWzZkOLjule9zn1d3MHHvDEvBNUNF4
BmDzu0ZucuhytdJb2BsZOJ8mlSHm2XAl9jdpbieWIvx9QzQkHghPOkbR2n9K4LpnCht6hB0uouCS
HvsvUmlCOoatGCVXXMFFlC3Nu8esMMYT+u7//bx6Jo87AD7QioVO9ChDaW2eHGLhyXpws2IjY7Pz
aTTTFTicXB/85/ZrqypklZH35y/TbGFTwhMHY8GzYjN72bcPPFvf2Z2ThEAvkYoeCbHU6kiDMTub
jbZfqb3mHrY5hxQEcwiGiQUU+gJIlPmJHQv/x/pmlTmVksbpHaq1Xcu5TQ3KTTwc3COUf11qI2SV
P/VeNn2yBlxep06GoFZVQiTzF8gBaV3mJO5Rgc5m2ONSYaBqnqHjLmwxra33Iw+d0AYpe+y+dF0f
7w4brb8ZN93f2GyGZSjza+zAHkSPk2K+HCUgYqhKnnb0b0WVT/ivXhk3k7IAvfRxIk9vLQ7cEpon
mDO39soJgh3YhFHwr8RNCuF1bs+AOLe2sWPvIP7u7H00DlABgOzfCLq8hvpoNhNvbx08Ls74QYR8
+f6BMklkDZ8k/MI3LWiwjZBH5Egj729+b1dLlPOo1uiizWN0vdCrnZTx5aQJcJhX0gumrxOx5FXI
yeQGztJriO4EMqDN22aNqBXUPHqCoe0oW4vUu2xqoSyWl37SasWPZXO+qUPQHbQz0j5R3dsCojut
/XXch6EbXvVIAixsxLJIpBTMGDb9oNTLSIwS3MPE6Ww99xo/jTZzduZcXVxl9o05dZGF4pfWAjmF
7fnlAvaw3k+2s4QDGHgm4Kkey3EFxQms3sNC6fl9jos2m4c8Cmms4VNu2XvMR33IJXSw1AO5UUv9
72Gou1/AgLCtHsHUa52h2/1kWFqLdz6ndKukQsAx3bGEemQ7YtHeZlNUwdB3NXLeOsOTVuPrqDHS
6Ha5rnExS+ovFjy2GKN6ehOy5eAE5GPAVhIDarlzEdfbzCYzU45jU5CmG/QHaDfLDYoyfOSU5jdU
zqYc9JCJew0q+5yd57MR0P0siwvmLPKHTFwYFJnOzvNHKatYBw+XkpRTHiQhxGCowJqvQmc12eAU
ajozslQBqFmBpRVb3in81uVnT0qQ4VVPjjbW64bQbtJQNDBTFbdyK+GhsC+Mkd0/p+fcP2VePciR
QajgeuH17V5Wzn8xy1WkkQAENgZvHt1Y1XNh4Tbp910mjSA+2aIMumQNsUoxzjRMChG1m/eIu/kL
ifBALLjPBI9TQhJURhwVzCCkY1yqxBojv4swRQduA78ZXPf0kUh3gR0WvRF2xC2JDaboEKboMCag
XuKkoWqFlO9hTUFnGo/0Tlwy7mjgfnP8n7olEwJkM2wH6jLutE6I6D/he0+X7xDsqsdXUMye6mON
OHVCtxU3DoPcEnZvO17w+7SW7FFE7rUv6Yc+68vtRrVYKkhGIDMAj3ZTev6LbxAt/ftJr8zrLyh5
FNoAl/2hNJ0FG8Mx8XbvQl5n/JpvmR5r2P1Bwap0jxt+/9VqTeFbcfWr6p/UiE+n90jTbiK5FLwp
VoqsneYFmkWkB0OL903TdEQUcpFgc/NrZKYD89uDRpG3mMB0gUMza5acXppOrcPZGXncovBaPCcj
dpRTSEGwtGdNVz06fhlLkR/DEFIzMaZ1ZpcAzvDOkT74n2HSsO+hwXowP49pb2Q7cCKTKItkILNG
HL+Barisbq2D9o96yk/Uqa3WKOePrTxw9H5UgMAxPwKqRdcR+DlfnBI0/L26Vln7uetSySA603/K
OtIg1ILXtghZxPiowFPGLE4bKdS8sE5mGRulm9Qtg2aVlkgXsh+aL9TdyI2J76fO1vReDaz2KOA2
NdTOc/Xrn8nolwCjsvdlAXWARXu5aB1LJV3/wCuyr7OD+KOHiPs6uZlJQNX5KZKh4voAHRkheYWF
6zSMtVy3z05asgpTwbvaGpPRAGbMfIKTwHkOrX9gn5McEKMdC0BKrzy2TuA0oKMbkc+xpg/dOT3U
h1XcfuuaMb4EYeER75T2b+v9Q1EVnMdpwLvVuBvYTQ9vYkTwrKedYvT98ihjLaO0MAVk+l1gA9UH
yxUOOiOQXiDwNhdicqDX/fNZwtzRKFLQq68Qemu5GVzl4774qCKhmHCAer4VI+bRlfXo5iZCEwVk
c3TVP+UkrNY2h1w+IOu6fChTApg+fXnPMXNcUJiHeWFcNOkYIcRTArCpmOIuFFjes0zhioZvwdE6
DWJvebqOXpBu2CORai0WaTzctxnQci55El6mYOjNcnuJd0ZV9A9dTzfWdW5gp9nioSNsXe28VeYs
27b7Uluco65tDCPF+d0UL/TJ/6zYevankVNfCJi8nJw14MlKmZEAdoWGOzOqHUNli3hCEdSM9Aw7
TPsYos8dEKuNQsl3kFcHmapwMW6GLMwiSoUAzKah4bWgO3DMZ+2+PWuJ4EV7MOaVzhvdxmmguxpB
D5JHQWwCx/PyfdionknrDuomESjs55uof4nAOXYUxYrx+MuFmEFFLZV8IaZnDaq1XqG7ZKGrwVP4
zrX9KXDbiuhEYMAkA3tWW7Xq+k50J4RM3SAYLm2iM9wkwGveaAhoVDZrdBvPzNSShVxYV5nhPXjP
vKpDGK0UzoR2wAbU0JkNGIaahNwvmZwS/Qn84CgwFDcgJtSIZD/C64wIhqptRUrbhKzNpCv3aEuQ
/+i+XFdqb/jRObsv6vw/aIH2kybx1Kdswugz3XV2vaIccacxhwhs4qyg2saVH123DoXvH3/EjaLv
qyWzRWB4ZoLDbY+x6JpyxlZqQm8ZXj00Wbow/V/ziW2AvQaIdH7bvio2LwV3ZYWPKOTsTaaYs/Y9
ytIjOeaKXZI7aWFcYuZsQnC3LX8YIM0xtRHfY38sow0SNxbUrxH4moK3tF1UC69H1s0P3plR1k1e
sAmZu63Zc4h8o/rjTj4MmwmDE/DrIENcd0vTkAW9Rh2hKhk46QVSBDZLCWQieubqYVHWqvBjDTiQ
3Rw+2dKDq8Dp8dlCgB7xPZhifOFpq6BTTzOYk5MChcCmBl3IqBFCUNeeHMHTjH/NBO8BoYgaefvb
i3tL273pRedcg0eynaUBoGiXfJ3i13g7wiyxarqiTWBaP4puZehepAZTC2gdqtVTNDu35ipajstL
tc/AdEmeJJbehj10ysAREDEEGSlbxAHmyGeEJO6u5VwrWJRqwiXG40nOmno+AC2hXsv3rmrA/iNJ
nbDF2DZyUl9eLVDzlOQn9S09KbJRbObpn+xfxbjjg0LJ+e8EjQXcKG0+rhfiT1dcTjGt2XYQx8jI
naXaq4ZLYFP6zOI4Wj+qj0P91IKkcTFcaGPnIKJlIABTSben6y2fTIPH4brDkhboMKAWW5tUVNNT
RABJrmaJrivlMm3A4IXDFe9H8f1QE8ZlNn2KUR8bwqrOiUJ2413Cz4C+KXTSoUFnp9v3/wP3jca9
5B5GLtoLpKD5IZPRD7QcGM3kJOpR6RUhrOxlgIkoRflXJRi4r40dhAbuynPfiir9y1WL/7WcBU38
DszAj87X2GJAwtoFo7GkIWGASIRlWwZSkuSwMcdnJXErgItgwvRPbezqxyKu8K0+JgKg7nZLhOrO
XkdlImS48aRwiFxlJJyjT40YRkF+u+5DrkxA5jzT5i0xRHsAswi5NrDJ4r93Bp1+VWLcgdJLEoic
dpWk2+UaPkGMdlc9c5c5umFl0dvfOSTyRxDUhFtFheevS5eu4m0yd6O5h5WOdCkFnXER5ZqUQaQF
AYsZ8eh5vOQYPXzCjSbLh5r9Zv6EF/EWfl5OEfTKoYLtqZLvtVv0KHXZZoTOI2qiGXnX1gWT6nPK
BJS05jLBv5lKO610nPkddNlRRj+y70VZgZN3Fhgwy3ZNoXrkiYlSbG+6UjDextVwOw8l8qdnhJ4s
rExfNJJ/zd45ozHq+ZK/NBlRga+keAjD5XjBPpHzbWmbEcNhFVfyxe5JhT2EFyaugK65MyoQegf2
TfSMQkVkm56//x+bSPh2VE3zjYenqPm8EjQ6fcUpsXJ8gRMXdW0ucxdIKHjIkyO2b/SdXXfSFOVR
MeHV4il83jEdW+u/rb4XywdPdE3SxUHXzCm+CzeJ5338WV8DJVj9KxMS3QMbZxS4nhnOMMC49anD
dBmJSCSFoZE31OewADqCrY8S7nazKBprGwaB4A8Rh8xDIQx4z0mEWSKqzkeYbqiG3CT1UEfmFE4k
tm2M2LTGQ24MpPqQxa6HL+mY9ZI8M6J2jZaxwzb/y39huokdim4XP29rP+EVdf1uOJ+z/l6XhmKD
RDNCPnita4FTtTK9aBVp5FIh5RkHGFR9b/sgHjqNyjYBjjuxkJiF8S8LLhiVeCB40DXfTa1CIYBI
zS9VFM+t1rlpJ8C7FWx9NWMBT17nOQQDllAEuJhkInChnLVi0qMHGtuSs3OQa+F02UEwjMUbR8NZ
3e90VutyUDhgsuO7dXVM3pKxJ4CSjYf5RmjS54XDMS1jhIZBy3WcfIeGltESSqr1+70Db+8w05eY
UTaoL4S7jL0hVqNgAR6LLv3RYAVUFxkQF8NYtkO8wCH4LXYNMVcHfS6q4iNayH2eGlpQB5xKFPRw
B4bJHl1mhpbCAL4jEWMrFW2sbXUokEuFDMemCa1cV1HEpB97x08CbiIezMyD9sQj9rgriaXm8TfY
Nn9mYh+jHh0e5BJkoZPTilGi+zPTMlTdE9L9k0KtEc+DQ7MgN5RPoMNlYHKgQlyf4pg2NHnjpKpv
Tzwb1x/IgoHCn8EbwnatJSt3otkZF1AAb9afUAX6gU6LIVbRzj2vAbGvWjtShKlZtU3X368AfkTJ
YVJACVLyEutGcDO44xro66wpS9CPxC6q+gm5cOskC5JjABt0eMZiXhFAgQmJOCQX0hBzcu2sKcV1
nSCHQQiuEuNqtBha8W0lz5XOp98pUGhB3vYK9Pw4vNvileDkrBt+QZAl3J0nijprwTUphFq3REkY
hpM1L5KWxvzrbgdh2AcOb8olNxN7KVSYdi8cCcY3Tjm+i2IbLA7wfoFTyKhHM6aPvJ7WG1sl6t4s
0hV9mpmMXga+JQMUY10QiIWmzIT4CNpvX3w7prc9//Ij0BjXXr5YTgCRuAwEvCwinXAaAZvg3bYm
+xsZnolV2z4lsrkzDyA8vYTtKoyPUer+WqTO/cZjVbQb0WTe3oReZizWJhRheT06rtPIK8eqt/er
87F8IFhnOvQqV6nYzjhBIfxAOjtfT151hCjdCr/m6EcITAz6pt/T5s0ldpL01r6dMBDSMjI1egC4
HYpdXQSC5EL9z58cXIE8C2MNe5l5vpLyP0etEZEDY6rzSDbL6Yav6aPjZuG/q+18yqoyDe8MJg83
DFHqIcxpojJQW8O0uzfdV9MugHDpkVLuJ1yDlIJ7Oob7Y02QuZ6TKaYT6A1cdjCYUX8BbNvmpLPI
6H1omp/uQoKWjA687yZgaR1DOEQVVMc4JE+2KDBWWHBG31N8C0fvPk7WtPzRPG0p1Uzq1yWgpR0h
ne+a1ZzfcZWzg8NROvQkz7fa3uc/izd8VifiqZzi8a3Rpyp57d1ojXq4IF4jz2LuwEzMDgMgw1Xt
jgCdQhqZsw47cq5OtsHnACt6fJmdoYUjByVWHfxbA7wYRYkgKL+Top5Hr+g98I1m6g+juR30D0QE
WrpamtIBLimEl42IDwoa0+WiUYwCfuSGry3kzUWpxSth/QM5mvW7SGQYjAaV2DO8g2pW3are2Txh
NxoKjiJCCtoaPrIA1BCThSmo5awiZpIR5KIDDFomc1SbF5hnCn0gDz1FeIbarJVqwDKsoLG9xh4W
dUTiD31JotdnqN82aMgvRFoVBSOznJaJPvktJ1l9Pc1Igakn5H7zMbwdV29oJtZFgmUNhXzTYnHl
PkXdw80xe+/jkiE4877mZBrXLUZcpgdDZTCq5DTO6fz0Ql/74AkV5dpLT6rJgc/sW7gkApCIrfuZ
L7NTNhBM4pWTZZbcgZQKlqo0w218+v696n2mcoDLzh8nnbeyJiev9N7v4xUoUrs2UWUsOtBiYmWw
dZwmYH8XQsMwmrwQNMOyPVtI1pZND5wFfjQymu6oIZtB7iPXXWyQveyabjaH404gx5v9SJyk6lKk
NtqOg9xmO6qewZFK/ddZ8uIme+lniDi4hNtVrC3nU6NcS18t0Rj+epg6e6l/rkOgTPdTiV6MI4Pw
ZE2td8Ndru2HKVMtBbNHHXFx8P2WPUXpqYUM4j4fyL2jylV95nAx+eZ/dPV1eVrl7GA4EHAUo9O2
RVAmog7jsd/cD8awvdxmT0udN3uE4PHYalE/zh99SSwEixuqV1fu1Xpxd+RJg/rRUTnFVqJiQoZa
LBILQp4CIzR4dr9OXJqRGYtQf8MwSghpCQHhTLBmbQ2wBN28J9dzb9TGf0wQ/4DkI4s/j9RPfGbL
3bH/0HOafJpLRq+zMkYx17R/0NFaosHNCo9xtynd9NmSWChq9sCP2POwgERUlcGlRhnHBXzZ36/3
coKu9pUQF6PcJm1DzVIOb12p2SOlRAadVu5rTTshKkXfZbXsyrxlIH81MHz4PAYDuzR7lCWjM8ve
XbCqTL3k7ZIc8F2Aan4L0otVD+BhNSRahRZrfT58oVQlipYD2v8vXeneC+mYjeZJYcL1tb0pIAst
w0VNHpOOFnn+3tQyx4ZX+aVGjwnCwPF5T4UFd+ZElCiEDF81vaOtkp5ZcVhYqigPVz2nTHwz0HQq
h+TYKYTw6IDU2OYb0wghPvkK7kv1ldxlm3QKnz50W7n7mww5DM56PhsVXbTrhbw8NmRt/5SPXPiy
eg5csGJ0gFIZPCCA8O8ATxYMBwek6cpwxlsPWhuv+1K6aGcas6DB8bqbt/l37y3FKpGpr+bzsfCm
YTRrIKjnibZjFU8lZfrnGevrlgB2n1aU56KDG71+k2bP9B55bTcxDzSK5TTnJiZaAAVmeD7ssrLg
D/ruCBstOedmYGBPD1noyNCPXgW1l7y+X0P1k1C9Mcz9V8X8Aq5B4QlU600DxamaLAVeZx5mSAzt
tZOQh5u8ldz4dHui1ByHQauec2XIqruF2enVJZTavEuQhfc0/So3REruNhDhvIT0xrSrBtImxVzK
IhvU3xnDBtiMxj5YNjioOZ4EC3ryZlAuFodzArThrLrcJZq011RYrM9LLIaYn4VQ5un8zXbA1bny
xL0JAxHG/5ZOqwl5LygRY07wqGWrVsJSOaoyTN+oEMQuG2ItebPwBWSIZdqtuuzJgrkwBuYJBN6v
Qq3EvUZqe7/4qk6z7KxBHVw6cxfes0/By0nWwCIjEk6KP+N33rTLtiZVMZCHQcVLqR1ClHGlICCV
1QH6i3qi6JJlsj1DxkPjFE9zQcdLs8dUw5c+Zw+YTZqZLwGvQ3RwOaQJicMzzSqh/ofy+WA8EkVz
ynV9g59p/IjhpkbT/9Tt6WwxPwYeO1ipEz60q+2pwc81NFk8Xk1TeGDUCgWLUmZ1EYR3PUGb6tud
/SL6VU9epmsui68SKpu9smOU7sZ03RfhH/lSpe/mnyT2H6ZTlHOYIiJw6KSecHIS6dQ8RIEiFWMx
ZSkPgVtJhLDfnPlPv/RcLXx9IjC1gXpFv5cDU47uEVugPSpWt8U+S/ACzlDRuGljtQndRW9KDrbR
TL37uVKZ0DM/zZ82LADJTUpnzJabE5ZH1BB/hrNFYtsSejVQoCRb6+Nv7HFa3bpMWrB9+oEWV9iJ
6oRqmGtwzeR5982ebDVuJZNQDiA6tYr4vOTJSm9fcNMj4CXIiW3J9CWvmabgyAADNiA+HTK0TX6E
xU3PNHH7q7QLFdNeaV/dg4ftoO8gWCo4RO+uNtCItnqkoSaBEEfaHEW08djW6eUVBi5g9TMbVZJF
E6HnA8HKHoXdKNh5LW9maZtP0l3+Rs/0AKGRWitm7Yk4FzJhYxHKaTV937zsTYPVga0QEV9TOGqg
fqK4ZvElKHawvGrGtseNsRFWeVT2QSLLl96XRdS2dymgndQT1BpPh97piDPz1X4qv+cu1Zd8ZmXE
syBCSeoJYUXbEzm0JPK4Uh+5bOjYDe4A6yMGB2l7LTrra3qvWoXmbtN5Xp/Cjbe/kYWEldqrP/FW
k1b3H4IrHRHBNPUh6pOXb19W2NP7LSA8kp7kRAVkCp/wplX5wnnWVXyzQXVHbT26KN0KmJIgE/eC
95rwzyd+3nqD3bEms/8PxLj8SCRO1JHXonlyMZV//RzKAZT/1d8XrmUkmNQKQxd3m9QTLwm/z9tS
jZCZ40SfZvedWHL+KkY1Sv/6J7zvmf5G0dgt2G0dSeY9NqZc2DJWKG1WB2jaDnLCKB3fWsM8TJtE
ztH5vayYAnUbMoOC0NLm6KlT965GKfFaSyUNrjMQUMbmcK3ve1M77krjqehTNBVGisfo+joes/No
6Uz8oR5aHVAcceFrKyCSyLH2BBQPoLS2EdraIBVCuyN4rpr9Jk6f0WA9K4D3mnrwCD/Nra7jXBWv
oiDK/UTTEuY2ypPxXFnpohQf5qTSGoWjb7U13tI/vIatgpOghtHiCjYLDm5rZtrcowzYDbmaUxmQ
x8qeVPbHzPVJ1UUlTMalpZCnOqFW1VJ8t/is5uuWYXNArFrSd7n/LSYgBycApsgZE3wOd9Us/ZzH
fl/Uj4XLHFce3ZRWw8NMMh8x8loXc6D7FV+Vi876SJswKEsA9Q36KKOt7yX3WEA1ydJHYHWhC6sn
iemE4IyTmRWPVax1vhZQlgc5vTiBpqyMLnkIOAEAalMsXRRZIlGpQrqfDO7eiiwjWODpIFRmZ13C
lHSfxvKNiT/iytam8NAmjsbSDise3IgTlx95WSNx4RI+V/fC+HaErdHvAVWYXJi4zly/EC34nn9o
d4vxwtvH6Y6DXkrA2RISyxV2c3i/LAx/LFJaK+EZnhgYNZNH+Szvs0SWSD1tCPcCAynNNJSFBdcI
0awBXIBf8F8a/dcoqLS/HSFxMsRP9qzLBMFBi/6asQcbwm71BDrQJAjZGL9FFdI9MeeQKrKxCqEK
4XfVE2RgDOyRxLGzfBoCTe/J2AZsvsMlyfppVVi0D+8lyz+pO5PJqUrbSztl+AOrdP7oJkP2VYhu
gA5hc3IP3Eh5wiPWf4coCbnbKwAORkmJ0vZ2v21MiGJGSNMKPWEzN/pyqQLfYIAFrdiLy3Cd+y2Q
WDSlKO+jXRDTBN0lrDIuTdDPuqfizc61fwB0xDXzmW8OlixyM0pmfkWxloQBJh0xI9HsHsjfQ4Na
QEc0O0mCHsknyWReOHQAV6hW5d94qTbDxkhBXttFx/kRs2j9Bw5MHM4kZ7on/gI4+zMvvAsuGpzN
a/oEna6NRVeh9JuA7WehSMJzXXIfkoZ2w1tZHowyDh5G6figy4DZn00T6VMgbIoCg6+4hz7wbG+z
k2TXSmXXk/XBUCLNyp9NCzFKxEyL47adSOjT3kz8iT9uLyKX+i8gcluAC5xpcuZbrQRVkoUx7u9s
DujD/XjYATAr/9JCQexyjiXLvXw9KDM4HHc05x5DK8e1A1skrPmJC0vcCkFZn2LWW7grgTaJXp+3
iYTufqYwgOac39/UYlXia06sq7xIMQyisWWgGHBC1sHUzZGzZXmciic4LMeXVqp8cVnd011kwxsK
cX8nzs4Om3XRnYW2mZFV6OmO7heEnPR2wAsmKB5ay24JxoFgGrI8YUEDwqirut7TStw1j54rOX88
RMyGfGPFWGAGv1xRH9TH6gHINcUBe8j83+C/tS/uLGUwJvLyDMzRUheBkCPU7c0k12vjfX4gfGh/
KgxVxJ8D++KMojTONbbKRMPMCRdMq4wtmbgXCEAtrA35Em/PWty0BlQfzSng/jM5sqqHue0w3Kbp
Dvkcn8RoR6zbqpVAg3OTwWiNRjBYbcBtmE1tHNel0y7n3ann9ggaYLYc0oWZ3NNpmKodUyB98/MR
fsQdbWHX9vKvZc1MXSR9sepZPi8ip7idcTtXkjyOroSHvhCkfV9ECaASu7uNg9Kz6IU6MVIta5hz
G93GD9N4QS7cmQtvq0Rt269+e2ox5lJCRR5PXbdvUIQ41C3UHgjjoUwBvpTnMB7J95AkJl8p/oIm
P7CsLZu6wp8HanWR3/2+6YfsLzDGjS9A9VOuT+wBV9J5Zyjz75jF0B55cB3TMAcYYVGGO1zR9WYV
gi9OVleIw8ogWNzIjKnK9sszYLevea1REbHyXGo0dh9KMTx/3PS/6jkcIhmLq7yuBZHylcSDkoUb
dj5kRuSf+0DMzryTAWmigAZZGf1rsK7YAEOZ24fJUesdwxrGQmrVdlwps5I8lW0v94qvPGG62Pn4
c2a2oLMSvOcuS5bXhkWd3f9T9huHSyN2kdQZcXKQh7XqXNSShTwjBKmuLXImf07UP80QKBsKdPOu
Z5ivn4Kg3BOFnAvc7zQxxqElEjNt5icv2KlDlVZVy4Rhtr11MaJ//46FqgCbX036kG7Q2pBR1g9z
6dFBmj63z59fOY+Y5ql9G6u9XKeC4sFz1IcFZSf8JQd0UMf1AUSJNVPlswdIp/rDtxaf+gwL2FPk
DgDKgPxPNMVKrM1zIoDhvCouU6zDe/LyUsRIZVABvWmD0sakXx+b4zXR4jSmzZVhBxN2m3CVmTt+
eh+R+Tj85Z73yIj1Xmz56YTnMzRy0HxZtw18mlSpmkgq5ollckuTojcuShgN0Q/yQThynG9MLqwN
qQRKliocs/cl63s5TxApzyUy+5wP9XB2ccVobT3n096qHmPxLXIvpfPf42noVBc19OK1okiAnAdz
QpFu7uCuPmwVMDe8bc7nIsq53ybAee4dXpYnPq+h8m74S9vA5Qat/Ov3pgQAaeJkHztIpLGmCvUg
EiuaQ6x3HLt18MTR//vFrVcYl9+6+KiQUN9Tqa0JYsNiRbMA4DkKeu5lsElTFmbgsHUzvzrcwRKE
LN5Sb1S/BO6phT5eJLaYD30fMW1q7pKUULieEGazFDCfsg5g3KtSSifntwctRYAv/ouWVlZPEqNr
hPOYfz7qvfEqH+vZMc2cZYv9x5GernBZpXeIX3t4/QiQpm5RKXjQ6jBpl4BEJdnibMw/2ENByorP
uPD1O6wLHgwSF0zhhBmFfr3st5x+zP6yk4OA5A2KcHaN9IDYaQ5VCRMivlah44k7IVCgTXUu5MMf
0TnlmoO2MT3e4aslgmn0ss8tLVptOKuUIaNpvIOKscAnH5uXr5IuaJ06WIqQNAjaJsn0a5DCG5/T
zLbrFHLueOKLCwg8cdMYvnhpmcRzJUiMg28Lj82lY/jzwjKLte1wzNY7SqyzYyyDwhLdq6ZfKEwP
sqK1Lu9rloQW2k4Dg3Ht/h/UR+3SCGrgR2F0Gpr0wO3apT8CWVngpmiiEGUDrFzIYlq7luHiMxhD
uAXc8PXpmEtD8tQ3EE24T//FJcM0QV3VBnZV6LkzpxeiUXT632f0YMCRY6dGHrQXPQESeRBu2kkB
rFZNRTXjM87dAyu7ds5jPkXohSmuuy0ahpqkguMJtZ6X2pA+hizzbOTWqxSDQZhWblL98+RL97/V
uhK9KEAJPZVRkxHQxtK6VhVAgs8+rlIH7zH5IvNghxDS3vyYasBPyK1uvCJLZer7nIDYvBhORNDl
9UA0uvV7B33XesjI+H6gjwS1ZGc3oXyI7WuGK5A0dvX+N0y8sKZRxOXI8g+SXRJoyHjAK9988CK5
Ow40YHIysqrMu2/AUUFhOaU8MEgRkfgS74k7SPMCMqo4obe74lCoSWYkUcGdqG/aAY9EGzaLD9XL
JaMkMUJ4vpnydEXfei2Z0Tnj4ZW0MvuGPGHrMiXw+CBYPiaj9KcRPyVAqw/p6tDpqLjy78KH/tQ9
whTeY89GGaPNv3jWgkqmwU68XOiAEHCzgHO8inKrF3gdx9Prifjw2/iKnaQvOLvMaSkmBvUqTsgF
d3o6KewaNUToZFzCLAj4b1JA+4Kc/yfwBxvedvoLmXp6mMgSxej8IJonk3AXUtMzFVuexeivMliY
Yj+g6GrIWToqLCb+AJ5P43743v27dq2dP88hJrshvBdx9rViiETemOtm2Jv1kO+BrNGn3n7U5G1B
mt5vyS8NsxWcTLBJmZpFVh75bXDezGRTDFNqR5yy0I2LJ3wg403rK3kWAO9lHkVWCBIbE3PM8zRd
mI2PClX+EukDApAPNcBeRHsf5mlcHeFxPJCuD7vOHHpTRWGdAYW6bLxq9SLbUMcWe3Q+8aSnApk8
aeWvJ9SrJzZIgLcgzHigL9iXe5mz4fiPFhloDyZ2TnoD5rL2/sUM3++hKICqQZ7CQjpbY95aymiE
Gz1jjoTV1KsDcru7A/0C1j595bwIfmZoothr69f02aABs/j5fCpONMvRP9RCa/xJzYIeggQqCTwi
kZTLZXE1QviZusnD7cRTCjPdtWlCdd4NW1ingjtiWVZtPRvNhUG+0OD2dY3IjOT85wr2cjW+Igjc
PPWc0+3uSNDY0sekKxIcMZlHBuVDThfwaAND0UsUWOOWrY5BAKseqX+DsF1bXtya2yGPL82Qj/PQ
qndtFjoerxGx7g+OiJu47103KvoiyFqnWq12wElta7nnWSRW6lTbaUDElunDKV3pjBzMu/l4yhxS
vdO4gr6jZTe8dhbLTcMUGD+ScuWzDdeoDfYZ9CGr37oX2S0u5/oLog7e4w6gwv1R6yya1O0E32kU
gT5wjdZaX5z0214kmVIlLFkKSpYY5GNAhp0FPtjm7BJEcrwJ464GcHk596r2wPsfi6tSHjxOQ8np
z03sOFdW8inifwjVTwXSAViq5rDnFS2mXDI5T32GPdq5J70fzHFSt20MrruDpfAh37m4++QH2EPN
QsNMNUN2pTIERRkmODyEfaNr2axNLyorc1C6NT7l61HpFS3e1vnSf4JJkwI+cNHtdX17n0DO5VH6
8pIV6z1Ztp4EtH6ZASVbg1xkSHkO6s0btmlzJ/SzUP5sITfkicFiYlehPeEuA6FlIagvm2KJUsHd
Q9mXnm3KzVBg7xQhLlDAhR6JKJlwTeoHyU9U8mXy0wpcHFojcUDkmF56wDapyT/GImA0bMzbs8Wn
Mxr1G+eV5p73Tza0EmhpmgDTnvLM12dolGJuEUT1/4VlffZwaSPuJgRWMEbTnNmUce+RNW0mx+b6
9bI++kFk/ocGZ2UN7Lh13SOzJSUEwubKJKuAi+vTmWVSWApWCHzKtFvGgz2Sk7NGXiJuDMaC0rAU
HaXYTMqrlJcyXzPVf7FBv5l6XgKyyhdg3ZwrS92/toovg3DX/6TcnQ50bM3/ngYp2uHNceKFju7i
X2EkYpIsvKA/Etsn6Y3xSe7Xn72xxQaq6KIaX5ByVWXqVIoi7nZLyBxi3OCCMU8sSckuBcCCJAnf
uZFgKmyyi+KXdMrpj4upcKntiHTKDPi+tvt3yaAhD0t5/h0kSBofXPtw3UbXUT9WjLXSwxbKQJty
hjH3C2nktdWanaTlh9TVQ7kXI8ObterpSyu3HT7PUqwkckENBWEKevW5Q/6kJMN03DDwYddif7fM
9HfLbP4ulSy0CmFO9gUuqPu9rg+wfKDqa7DczTeqzVkCIILGgoFUa9/aY1aw8znOd8RTzM8AYxvw
ciocvEHTia8HdGg6w066tSbE8xyxWDg3T/OWak/vKAg0iMT6ja4U0l3YZX5vETkjFflYJ0Vh6gNa
Mwswa1oKkhjCJ5SfQXadS9sZZNEnZxrYmwbOEQM7SKedf1MePKeHsp6NYv9BShTnwVJfjI5LP3VP
uq5jUha3ru0+lwdwkD6gEhX69Y+3eoaAtKiEaXCmbUCCIzSDFGDWZJEuqAAdi0EgU44wp+1ZmGYQ
V8lMAf2Xsx21WbLo/is1MND96AhhOqXLtp+FAyWdd4ReO1ZCs11CDfD3T3HVPLX6D9SsXx0RTvoz
/PVKPBtqFbc9BHUFOF2ulIpCCInUzm5Mpdpr9ec53TXmGaXNYa8IS4t10hLjiBVSJfwPseIHLqGb
6S8zxhf2jbvjbpiwMw3TpQbbc0Rxd5QjRZDowWsKRZqWfP697VCak6FiSlPSEgc69pPFUasXz/uE
DRaT2PtWyywHj+Jjwwh8Azz7POeHznFQavIjG1msquKYdgIx2CCKeuOdTOXT8xTuQfC/UQVDA2DQ
iMjQEo9wFReJwwI3R5omdMapqKFAm6HNayYDeSAbTa5Su0PnzkhNZeJw48zhVTLpAUAXiKhlReYk
o1FtPvuotk4kSYXJ358Q3sDMuHO6PTG5CGgJMXibeJHrewEaheH5OQFzbaWvUStcQifBHS38yCOA
rH4OQActLT2GKrb2jVhm9/rBp6qB0OaS9ceHZHbojxxTA97eVSbVFBlPdqHQHnHLM704IEnn3hPL
L2J6wTVh/sWHN/SmiR2D3anYUh9icchVQyZhhwxcccD7BHKFfNUWbuAgGh9cJJCk77/5Q0iENpwq
lSFjE9RYRFbBOAGUkl3Z8Lf160angtRIkggobgDggAwuFPQngMKiOvKm6ulUamItlr1N8Bau9Ofx
vTUyK582ypAj9XZ35Pza9PbqYU5aCLPB4iGeSlAMUUlOJFLbNIoRr77PF0/wKtEsiJEzHXJO1HIF
lyVTXJQFjtOFnoOiImPy5tPT6ejSy5gtmrikj+5ixxJ9csi3Dqm3C9ba4iZDg+3FW5yEe14cIK9F
NX5zOaRNMuAmP5N8QGyZ0UtgYaIe3DQedAqqb2SeaTtmdcmMloz/wJSwvo79F3dpzvsvLOS1pPNR
U8R9wgmPmBmIOhP91zNw5XrqKivgFti8D8I0rqt8dv7PiV+zqLS1LQbkbX0NZCajYBle3yh70LAm
ui9N6uPwSKViaGbmOA2OIn5htW6fiJ8mY+l+u1Nzw8aF4G888bT7qn8W3+3dnnXpAlPQURpbHG40
cveos0RgJ2RkqZHn5ptZWOrqcqiTSGy4NVzFWL+Uhhz4Tvn2d7/r+bVPPJNxcV9/y9KfsyT4dj03
zn3KnSaQocg8GY3gVc59M3y+L2dQoFcn5Xb8CDFWrtK9VxOI5pk2GJYJdFvqeeLyGL4b6c8680Vc
Bn4TdrinMJ8Aw+LXzgAwYml/Noi4s3JVcnlhGw6OdwffqKh4Uc/cMmTjESOIoKYJiHJx3nJ42grI
ZBQ9S5ZdwMGaX2nFaN7BzrHbe6UrGNjELAPUpTo//EjseKzs7YcxqLIBlpXaL2eitBAO4wLTArDj
al4GD8X6Y/oQMwJmusCUnhOKgKxTnOlblCpgJdZawWqlbV+UNkCivNxYOLw0e/czAfw7sriJFa0j
eESGLfdR47bwPM+Ldp03OJxLL8rh6Ljzjj9xnnUUzggTPITUO6p6LLCuhrj0aWXZ2w55CCZKBrb7
dpfANrrtjCy1hAhMt3jrBitmQmqsoHSDXxcDguTleUeiHmpaelu1y7Yd14OJRBAltmGQL41aJfWv
VxMzAttL0IhID/0bTO2YnXJh93pfoTZRQGw0742k/MWrpfOoJvCQtTqCGPwTI7vdhSrXdQyV7mpj
qG8qNsi4yaX7OIT0/0fhL2ye8TJbwdnWh2HwbXCiasZjQEwUOV8S1WW47AflXKUNkee9UFCVGvva
PENHP+OB5fIWxvI9wQi3R7IM6AOy1+dnZfMnRQTrF2/mo360r7YzVekkxUgWRfrvnocUaOqmkE5k
wS+rSaM1HAENVexYXZyN5gbi1NNWXV2DfsT0ajQ61FNuznvfhBhPm4MszuKrd3chrU0Qdafc9j4l
BNSX5AFBTYabXszwOI9UrDpgKWEjJXZrWopykwUyUL671OSbH02IGxn9GspbR6VNEBh1oVGR2Bdy
IS12qKFLxcu7+8+FxkMKy2ezrAzvtgNDEcXEWF26A0sl4AvPubCVeIdsdEgzyD5oKhOTXl6ooPWP
tqG1X9KMEHsNCkzvdwzSg7Aqlw2zS/qsuISxpraV3fuWBvPzcRXJvi4K2tT8THXMou+UzBrVpDtu
4oNMVdWBv4NziXHM8iJJXITiqn81i56AhtGGY6xVPiDDU98DeoFiTgGudpq0nLkdogACdZ43pOfD
4y04FUFVkLc1vKmcZ5dLoVogDnTN+cRmkkrK7gEHUzy2M6rYj2owPF8S3M1wzFgGylPj09jkr0Bk
osiUDQ7A2qgZSrNPSdBWC+pVymOKIoU4HE/VA9X8SH36rijve+Uf3v25LG5aLI7ONvxLo5hecCY7
7RQDJa2s1Xl/WnQfYyAKpwKRf9SguRG+wu/SjWoIjRjGA24YwBdjF/7ONxYJyDVX1I1wB80rgSZr
i60Uz0oyzk6yh/hI+mMTrtjTwmWa2QPF371saLGtDdaMTZKU8pe7ur0hMqQWn0Bx5vu+gAuDBxxO
6WP/2livtSRUKUt5JSIsAYKcjlsYQ/MX2GraBcqiDHW+yPnuRNUNUEtrENdiShD2hJLKUBtF4XbQ
KWQVkhkWQj8Y3rwubPDrHnD7e6BpbdLimViewSOugH8KI/45yIcXT5NW6HxFZd42cvVmGtUIN8si
PuJiVMMcX6qXaZspOVwc7NDoqvgZeLr3gmKbmGdaC7d5Xo2sZS7uZYUImZU+dgIfHALZYuQuYxJc
/ocaSlx/TPZ5C/5qdWT4A1JNACUHtSEzPG1ojunlsONa4Q6MkYjUuYIbKhhvMNTlzIXZjDCyShqt
HkgXspGaa1UvHSDu6/1YFiVwJoLVzjxt9PUgYI/NrsSA0Krxz+Ti90rYghm+0IMRBhaOtTQaaIU7
e2keJHWCx5Q+aKEg8XhOan49fnCK7JLZXBcFn/W4YSG9ZuhT3gR/PTnc+8hky6Ftl0wm5zuQ9RGM
tyLiqueyBrkfg84vKvgifg+r9v1yV9dv9pZ4Rxc3Qe8ER2SbQN5AyIwTTO/9rEGIHa1BG+S9F6+z
fm6OyZaY4LxEaZPge8bwRVH5HLUbB0tjWxNkNNZwHHtiAFc6CN/gZ0K5eEYUhmKII0Pa6Be8xe0q
Tcyo01ShaPxRX8+Es4f1+KC61gYtbvja4tVwLqPRmOWqn/a/rK6EJzTu2orDhj4IExNV5ItgSeJ7
hxS7/x3+5OSDV9Eee2Fe1I+V4e/VieCs2yoN3n+jduqxE7WDsr7UlfdEA05wkv/fnJWimA7eOvzd
wLaJkec7fJRnF8vd2B5JGdr7QmvaeqwY1bf7LuHtqTq02X5/cvHmQO3MufhnF0fzrBe6waGgkfbF
Yk7A0zNBfmU1o1hnsK6Y0t2V9nyWJLcvtcx33WvFFkCMzA4e4dygjNw5Jf6229cKoeDwU+uj5PLZ
pGJtQQcpAffm72CKWnNHYsERHAfTZdlTjHrxT36fh/i973awdVCnN49gd6DGqkTAYHoRWqfA0yNW
LFH9g9kbWxhog19VYwMKQfJE81NA9kzKmZJXn7OA/jtCz6HXMpkQ+TjY5BYmdfjP1QyZt5iFjUT8
qKC0cW8La40GmaXUXV5/np6V6oBEEWsDMrm6nckzGt5PttwglkuPWRJKtVeLp2IDHpApvvjs197k
hqS7YKcZvPvjeKBRwW9QJr4E0xeOAjiJs0gZ2epICS/L8J+FS1EYnx01+d2w1wDDNb6f9a7xUNEt
OJxY7Q+mweVoDNI2QO3tua/G0LpBfH7TRstE+xgtA5+sYZLR3ZepYHgTLbGoNLamTDwoeKaZM51B
gvwe60ieIM3ZtC+jgAiq65V1PjyBdGpS2rMt8Niol4KhHqiHnL0YulDiAbpXNytPV3iTIey217Qm
ewxo14gEi6z9cMGJqIPglD4BpB0k8FVsujM7K40odecH89xTCzEFNS/8mF77R1vKNjgTBNR2QCJa
2oLqqTyGHv7recZ3NCuu2ZYJMV8czT6B0WI0f8kEJNh2eg2mN12FfsmWocUnA5OEEf/ZY1PpbsTC
WL+GUUmo/cmoJ3vCwScE6aUp6Hi/Qq0aspTI9VW4xECVz2EAF9ammA58xI0tjnqZsWF2oho0RwBJ
Wa1zt4YkmBg8zPT9dV10miNq9pQohx25PHgXDS4RMY8qo0j5LrpYVimEP1LTnWZgoaj/HO9Tv+Qd
UYW5OYCJCeftZqgLwR4Rbf04P02TEVFQ24emUNyxnV/bGZuAzUwQ1pg7UTEdfxPdDYCCQASTwf3I
OpvLcr7R/i3Q+ZJwjMIVw/tZtF2JFlFxf5EEX5uwWeMSvMtWQ6rBbeu1AvZX2PXtg5d7lIvHqaf9
v/x3hsz5DbG2nI4BGXUDl0SBCyZoXWwvXN9xfXqegmRYHC6CZ3SyQoFEkJBtuwulGjujOxFIR5Yd
0suyiih/SupIVY0UsUf2aomfCwMxOKp3kQs9/bcpFaLomSD/jRnSszQ1ZN901lxzm2Ii8NynjMI0
c+mgy5UF3g+HCFEK7Ls42COBNr073Jzl92IB+irGyfNVpy4ylkEZwU3P4SUlaXHPnWXXcRX1rIVn
Z+4gV1WRf9rUcXENfgoRpL8KwZGAs9vTDbTnxmTA61hKUDOHyyjnjzU6rrRKAzwcyoKFz7Ft/Lgw
MMuBAzI2OTWjfFISgYMOzEAihtM1vqp1PtdbzZEHH8q14TnwRd4ZUTvj602IhOUU2zAO8ieihMqK
FQDxLWMp7U/6PTuINXPFq831AvGvUDZLVjiEuzEbV0MrPhL5mnl6dFS8hCQIJIwByMz7VRHT4O2I
TSVz/E6n7waff0hMKO4k+6XIUKQEUTQja6WulKBN3OCSUNTByAorqltRjCpxS+VpK3x5HqpcaFKE
suQOOHs2oL4GI7qdFQG7tQ/ULcbI5hS6Na5j1HvcEb4cSLAjR8MWX1xBcdK87I1rKecoqXeZz8JZ
ut1wMClVbV1+/mLOAfV1asEVmG79PvE/KE66wo2gMHQ4GtVcH+P8DSaTJwvB97dgNVDk4hF+5gjX
Yc9b+E4Q70Be0sZrHhibdFZxjKJJXQfLbXVmjTa3SA5tTdOPhmuQdrQp1ADBnt6ByPM/F3THaVWW
O5isDGdGUnjiDsFhzKBBbPTPoltyYY+KuIdZT2jwrvg18uJo0AvdTOCWqvMMPGKyTYaVWKDTXF+P
X4q8839eRZomiz871yUNak8vZeW70FHhDXy0giu/tv1G2akPIdgwn352Ssxnl/xKT+PJ5so6vmg+
wO3HEuB+a1MVytPFjp6k4UVxgHhIWEQk3G5Jh54rQxPw1PcfSyktb2uuoRlCOF29iv4HFvJlM5t6
8w4NlTZlPGArqCdNdd7Jn1oCqjMJkhl3upr6HBjcsZN0z/prTF/VThUQT5G1VHnBZvnWyeE2jbCw
WEub+eJaqtO67ih6yQw0BOrNJwxfBhILpCy/AVKD+p2fdvV7/3jAAYPeCXcbHK6mG2DlvScvDcF5
kM95nvL4VVSKDQciUU4CAm2YmpPkWq++OnuMRghqXUn7jncqqdwoWSgOtmkMQTSBcnxCjp1G0qC6
8sgm6yUBOoazUVfvUZECBFnYZErs6entSzRRtHOLDVl6xq5OUtNaSXBAo2k+W/MtyYHXYIRlLuN+
75pLerTwIu2bqrDsg23s1rUMkV3TZmBuyJfm6WvkpELfRGZ/1/9viVZeHvoPakKreAxW38detQ10
I16IFQ3/+DzB5XMNUXfw75x96ok84inr1i+mfMzqZJg3qRVk08PS2ibZQe/J5x//UzJFKjbUC+CR
idADz9aQr3mZs9wYQB3crHEZS3HsPw4YKKQAlMDQjmILqaL2wtIWlywBXmoOsTLJa79x6aSK/VhZ
9lwbpGEcSYX3V7fAnZXOjXTTA5fewKTUsuZYzCtcsd6PFI4oGMHro+sPb7EBKArYxJWstyWM8Eq7
KeEuj1Mv9w7OntCyyaHOvLHiz1RqHfW4kW8SIL9gIwJ9J5l7pS0xkJzsgQ+6SRJhrwGsmaLCBotc
VgzYWodJ4NsBYQM5oX6ti0Du3pUkptt/+WiyyBqIM4QCYWmV6JBH+ABqw4kLkqhPZ4zgHLz8gnVM
TlJ67F0HLsbg09mqAEOB67C/OBqW79X4tRAK/N3ATvs0RDR4P4Arh+ZTCwVmPZYfz0uNyKQTcInK
GsR4CFWtFfqA3fna5EmE0ALiSd6TUegoV4WNNxUkxDt8KnMyFYSbc5T+r+aMeVM1PlJx8l7MjfRy
x6a7mMTJtGrrlyM8J1BaejoxC2/v2RsMDxWgBIF2ZJXpPXegA+p04KxDCE4wL8PCYhRI6Tvf5+a4
wsJKQZrI60aWZM3zlh/jxXVIVNlauzc2Lw4WIpcF5t2IwnCqtsDZQzwAGXiaWhGDu3MOvv85KmpN
zP8ILU6rMdShqRuacw0R+10rbmjHzXiNPt5GCfwDrN72U4axyFQvvt4DoX3+H0wk8MUasj9XcKhQ
9gGkwUScUG/jBvLXCF3xc5Aett39gikxGL4t4Cm1dersgwgOCHmSFABtcDroRyzPo3OilisWirOO
RW4NiJL/lMoU6zfyujNclGAePTALl5hL65+Oh1EMtNP642UR+hm7tEy07jhlf9mQayq0aLc5vlA2
nB6RUvDueGsDKvJCQWCXbptfuGsWS6ZPJ3o8lyYBWz8hbxrz3IMXqI9XnaPSG54eDNGMg4ff3Qxe
0UJFPLLPRDggSJvaRXSypDl4zxhCNlgx4lGaiN45cnNRvV8lta7kFDzdewoqddRq0SmDV8JFegM+
6Rf2MVQ4ivAWDFlKxB9Lyw4Qoi13mWsmfwAMeZCxaZKJ+dsz++I/cDjEyDP46Lx0/7RHIE3Afsyz
ArDjO+Q9QtMvzAoD1X40ngBqaknRi9Hsgr2lTJhfBV5kspM3/SkUWyBFp69GKy0AKIDnps0IqMMo
mipG9x4YIFqdeO8lfQQzpihDDS1zb3q1KGOK+GkIuD4iETRFmpJUklCvLyK1KOy0XIT3N/zX98CM
l2YRI2SETovWxNLFN/2EH7YzWIqDxI15MXyqZpY0dm1KXgg5lVAWSdZ8phACk7QqGQ8HVjHGm4x/
36KBicV0HGP3QBxULW0Ytss3DOBsIeaklpm3U/guwSMFa44UPNm1T9nFYzMYCPwLGCD7tZObJhC+
EsUoNDo/azKgQzM+96cF4yuDHj4IjxKQXrWpVjmtrEUW2cYds+7ONorZxiQE7gTlsUTwrWlyrIgw
YR9DEWBmJobFp3e9NaTwTGAdv9gvScTRnZ2cQ+Q2d5cpH+ugeZSIoudjUMP/migwwYY8ePU7Kmso
RIEiSV/j6qHxdPNeGMgnjYyiSLMrt2bCsV2PXLAuWqQX6aHg2+UH9O7QlLtQM2pD0qWGhf7C462s
o0a2U4vmNVrnH6G755WPgNCAZI6S1wmIX+2uQdDP1dZApuNJDUMdF5GhRB0PP6FN1WPac69D8v0l
zXE9uQ3rEMvQ1gwtnfJPIYqRyc65ZzGVuPIvu6VkGI3NSorks6cQLRSFHmO0iTRiYk/DVQjvsjyL
oLWbUDlVLBlYMjsumM4oSGECLUuq9GAOjpwMWPuLvSsofAzPDH/XScEEhsWkRM5Bactky7SZSE+j
o9VXm1vXxAEeJhkrEdMNe77Wri0hsL5abMf/TYKXlKlujV5N4RNd515fn6OsFZqkW4TfdcrDGfVz
LJgfv5D9b6IZI7sV5PDFrVtcrTGI7p0yw9BiyA1dYfgIPYYXYIlWiJaRlP3hp0oGRCNkvDpMlkJ4
XeSxnISnqkdcjplbeVGH+m7v2bk0ZO+pRhJHLlYNWjivt541KcEloEe95XnZCco39/jERKzmWhVA
NzcSH3PTYWbSRHZLuJU0qxIGpfERnPDCiUq6LWHoX9WyORII4YbRyuXP4iVMsZkMZELqjh3Z6U2q
pntIKvtiwiCWxSSIyRiuLr9lxzrXN7yAFqjICGJQCdm5bDebxMX8v1CMmsO50gPJoFwJxKhYUS6T
wbF181mOsnclsv44Dmwowo4IwVtbSOkCm5GkaoX6nxxZpb9ld5rohgzz+Jd9rdtGt8ovrhZy0wtD
DBZCxg5ExKrDIWE+Bv62vQbhPyvIeyUk13GCfmaUCziEw6FDtD8DAmdb0orZMWpbX+JIEHupad/u
0jK6KOPNTyK8oUdais1dn/nAPzQCbSnRKUE5fONvvMjR52uw4bFyhbYTud2QOZjowYspFywygJXS
dyjC56VJ9rfe/n0sn5uwji5ppEHrCqMuew9Eu9KzQeCAs6nkItYy3+6Vh8t/i9vBOcfpe3xeRN4U
KC+Owu23l872oualkoxmNUqyNUb6BFuPtcU1B0TzvQgBquKoKc/AoWD1KLGrYry2riyCQHlpcNBZ
RHgSviGDK1cdHW82xkpVwYKbY2xw/EyB5GGcOBQEKHiAdZTQW3RsOuxCPG/w9g2j7myULDhO6vST
I/MkVfhq3A2udErzoSGGVqx56LqgZPh3prY8hbah2YWvhM2WWyz3opv4gI6bGceKsfv5q6XBIQIK
2NDr+/cUJx3qGStMvlzpX+ULJCFVZsWVlS0ilIq3LhtbevncG1ym486bqkj0EU1+0+uFs+tbvzd/
Miks4PIp757mQfeWe1gloZc+nAw1KwuPE4LoVEJqifRRi9ME9tCngxJ+zMjqt4WJF8N82MlsyCq1
pL9Q4Hl593/WlJDZOZvycVys+4TNdU61l/TNn1+jbQSa1g/AgqPmXIE7BNYFZ9rMM7e8OC6DXshf
6GJNLMXYNlPco8SM0zCbQUzuFcBW1pZ7pb7PzlgTccImJqaDbWBtnnJtIKKK1jxhhlo5wBq17bZ6
RUlUqwp/v0b+n6N674fqd/NoaDpfRBNFSpNaWwxotmwkOJFs3l4Sk7vZWyp9nQjUTxRpiUhScPv/
BhoUtFwVZhDfLv2P/hANK6EmVF4oTMngA6Xa0iUC/WoU0E0RnUF4KIkl3FQgmWhluYPLfDPaedYP
2pQgWQmgdGdCf9Ty8QERk+r6xpIMOtKEg89kZ+6xKskYWWy10kFQHiSS0YmdfkTA+gli+Nw9DedT
ejhOi4LKprgXM1JJCgdwrOiKtwzGEv+s0Oap6jY96uTnw8vqK0iS4djsTgTOztSvIFX8AawHry+g
ThGl7ByBGqIZPwQcUS3XruWo++7aqJlrX/WVZvM/CazRZcGJfbVn9KToe6wLh83y1nUkmhmg3pVq
jaNmI9W9nN7chpBB6sdkjO0DyLUYXzL9uyn+MKGmxRoOTbg419+yMt85UF4LiSQvZgnJLeseptOp
C38AGIwY/lrKSVuWnVdWi5oHKdlu6OihE8PgDm3jOF59HKvIHic/tOI0kxVyJrPgtK2BECJX/ZOq
eCLBWAxW7wBJ6aukMrNXaiQTJ8a5jXGQWaeuvetcFdiKZgLe8P52UrbBSvnN5eTS8jA8Wmmd0mcw
UYOqJhJnVuCmFDyik1IaZAJd5IC/W7Le/UYha1jbZF+N48uGKOP7xH1cmILcj00SJXkbv7KZ5/tl
PP1BAPXj20rptlOTC+Ik2x7mzIYCA7pHhC8FQm1B4ffBVse1/q1Ys8o26zeC8Qug3VUIe8Bs7uNt
BT7W0yhFaZ8XZyeWhVf3z4mztf6BKVWFCTN7jludjUCfOdYVOoAav0JiuRmn2sDnJ7s18v/nzeP4
eCH8LUq85MEYKDesDqIVmeRwon8wEdADWZDgBkNdFUtUmx76KcsS+T/Lzuso4XL4TxZ2xpkcOzmf
x02d1JXvvRhnwjzn6rOFNrG5v7GlTJEnhEMIfnEAzEYKQmFGGhVXf9pfsPVr8873pE9Sc85UkKz0
0FKsxxy44eTdS1dOMRzAGHYQtal9AmI2aaJqmCD86xxcHLIdWi9NwsxoZ+euYBX2HYAlbyVslh/m
VD9rYfouGhDNzG0DIy1rojV5kYCd5GZ3bMU7NCLYIu8luJ4mE64lqCbY7ckUWBFo+zc3e1fDb/n9
2U0H5mRy+pr5i7RRdjtqOYmdvnWyWIofBl3erVPD1kou6KJoak6YSpFBXgIQfI49QN4X+Zg/vlvM
YEhyPYiaJ5V7HuH/rhSaHQkF2cGQGLuukz8+z+BJ+i34V12a2eS1HeqoVQNc+CDD4iCjROgkmMPu
6lXGzHDR2MqcENcrt6TuJxV5S3GO4Xtig1Bttnde8gpYyFka9omgR0QqrI3cmBUVx+479NN/++UP
y7jgiDNpA/HHFZho+uCt8CTPsy8h/p7EP4FefphXSkYDoMdVtFue7ubk6dcCZxsmDOwMPiy+PMlm
M7IKPCwlJN0L8rxpkQKcoy2D4CKKIRlETNGK6BHrvbAxq3xy0n1aMp6VjRVVsB340XZr1nlKQBh/
FO08vfl4RLjpHgX2eEL6aOy+jsqhkp1oJMGhnCi0FCKHA2nG2DK+I62g4kVWZbinGpYkefLa8w5K
245+w7HvfVCgp5GhWc6GZ2GdhS6sqtWhWh3xBwzxEy/3GokQXTOyjx+XUFug4RSR39FnKYAuxxmN
LZ3g5VOIVLaej/zNK5cNekMrc8QrRtsMewyaQNn0j9kKddYlhEXgfsZBwKbBEaikyzXKxQn3+IuR
+/qgD/pthU83EbzAnvceFbPpoI1ha88KSeDsqJLVamLLolQfLyud7QpotVoUUkKyUhPpl9Hqx7uq
Zpn3oYP5YE1ZeQKocChxT1cfcg5dBPNxrfa8q0k89NcTSXGzLNxfJq/CU7v5d7tqQGmV0UBx558k
5kEHeUg/nSt9fEh5hfQnDk8e4uyHHXGrhwJgTUcL8mc690B2tDKHWDhGEKwuNIWa4dnxastI9Y6g
bA14PwbI31qVXmt6ul1QO6RVMrSAGhg39KZ2nbfebIa9QGuq6eIMoierb91EK8KqyngS4D0Uzi44
fXMWb09f3390HDxMG2jNBj8C7miqAAS1kBPNLb91Wc9tmLT7Aw+MalB4DHq6M4I/A4Xy/Ma5ol8X
TJ6cpmDEAyU52zYlt6qvneTxvKup5G2y1bQ0JDKk85xlkYJir+ggfHpIdPF+e2H4+4rFlngp/JL0
W15GFwNRb1wd4tzg1Cghc+ij4X6VR4OQhy7x3gGvKet7i2/q0f+cvtwi4Ht3cGrF+7P2rCqIoVn8
MY6ABKJ8njd5kZlx3Bf27HSVNtuAVEn8f7MFHJVVuiJFwASswhI1CCPkeo1njGtLLjNdNitGoH5U
XnV9QyGrGIGJXIAzp/YBBLoJ+VkRtBe+WlB5u92XFtUPLn6hQ3meHtKbcszrvul6GdK6r2EOdbNt
dhf7fGZrjwtMY/f/jA4D5taDabI1jhQqUiG5QAc1ChiZrjq+5MuP9U7LPUYfwES8uFTPadc1oe57
vKlk6W1k7hORVvg0tQEbqyvOVLg3zjc8gIA97BYExCrXKwQRkMkE/qy4VgXWwKsQrth2O0NY+wP8
cYMGvT+Nxtp43LmA+3Ocir6GiwpX58PtFz7VZRdQs00mj7D77AGR0O9BmpxGE8F13WS9SwIsUzx4
KrBgCeIQB8ZSCYRfwhXoN7rA7qpcGiowHpcNZVUVOJdRBI+oWDb/c+bCUdd67i7XIwrLjV2vqGkA
BVh0N1JUlzZeyPnAp52V+DfubmU4BWT0FnjNXqja+LT0pzux/zKqpvmNelUcLTpGFlwRElbjl7QC
4HATx0KCXteHdwxOoVuSf+7iBzPaoOHYHGSBadzNyqiZ8poKvtMTPrPs3FKKr6hTiW8+OfcrjpHV
IEODe7/kMVC3gk/m9RXTETY/Fm5OthToWU1eojWu1qxGHAYX5FBPIdhuU9UngMrWzKaGTwEB3KYp
BqzpCqVKdlRLeLbsN2HKxPNl/IxWEkX/qB/L2oEzLDntEBHiAJrghAkT8Z27WqM/YwCbgkG5sp9L
aez0WHDmYpUmSP+ivmOLGjcyj3dL9P6mJjmR8kqoKJIg/GeAev8812PZMcEr7zpW2BCeE6ccQpqY
gwMWcIeK7/Osx9++8uQu5Xz2nd8JwvnQHM5Kd+Huvseo3NN0/bAy4k38vQrW3sJaZ6+he/CvAf4t
pPE1ok0Ilf+zm0L5nIyjEqIrElQi8TI6HSi//fsOd/UvtSSBibJFEjcBkhOXRIVkPNJ2IiyBhJQS
WK9ptgIq6Ay5vc9ADc0eC5shfhMfK6o8E3jcCNviJNuDbnfoZJQnYVnhwkxfVRnk/8749/1r3Zeb
P66tE7jmp+VTls8EoNIeVmvne6nM6waGTOXrQeKy4SkOm+wDs3Ngv6nkawnP1z+dBNfTc8swjJB+
FApBlM/upFkpXDUDGEZhn+tDNRMWJ8yJCLuGJ5XMAJ1kgi2sgvV+evom8qAFIsSdeNYLnv76UBAa
IFDdDXrDrWPtENStLTpka2jejKA8Cf4iX1yWc4BIQ0VtgcO2F/Yz8YWbLB7DopFNB/dCWUffrAPi
2eYUtfoICHZA8xBNCTsqz5IPV/IPuYjMSwlEWwyh0Rx+l3Eh7IOw3FxQDkqoQPObvM9h6HqM1/KO
Haj+YNw2bp1PlKlAR+Q2iYxUT6TZY28B3UVLA45e3FcR1wBBtKkd0CgYfoj8jWC+UDUbRu4V3eLw
Q8QgjTWYxApuuQ2J5fk6zvJc/EHMRyK5nfnaQF/jwynMZsmJfqB6UM9Hju4U5g6mfbJa+2Ku8lSY
NE8IMwI3bHiG2jR0lSAbS6rbxzKmkahCAUvk241OEMgEmJ2H4gYEQQ0yaFIPN0ArC7IGinECiPVr
jwF5DEbkoSeLy0JmFPdbY7OweTyUIU1yC1nNosqqSdYpSPjH3N0XqP3TcGerUVcPU9UF1Rwu7iC5
vhrcbUqVkxVaCt99gjcYjhfOdrGdW2ArENZoe2HFNrn2+pfGUk6YB2r/8qccH/lXBro7boqtvF55
8+zUQUzs/TaOkPFeUryK/2ykXzP3eBDz4mGU58E7v7hq3tMbv/I+5R5xETiwWncu5LZ5ti3bkqlI
UJWtCX/M+wGYvTYoWLmU7IxV2JR3DBT3bGa8/U4BXA+q15rkbAflybeF9s2+qiEsv1UEyGAONHcR
qk4a8965H6SByl9fnmm2v049WDlizfBq4M/WFjJg3Vu+kiCGHmOK4uxUTIurefog/p5VYmWGQ3s9
Ff1CcZDikBZWBOG2uab3LsNTntcmcRA9L998nhroZ6r2Q+UP11XqJpSV7lomf7FoPe023wbFWM7v
pYjd++uPOA5MShkKvuegg/Ic8VnJKniRhQ2+K+HTk8K0BCj+aCwG33JKsUSkYT/Yw63HxntmHDlI
3lcSGlz53CGzV9oeybvNgt0WR77odgVf6S3LTEy5ZNEY1NgrWprEB493RIAN4pkonYEJ5xNUbuJf
x+Davk9cQeylrfa4kY0w843c7N2MOYoN4FCAw0Swrpg767NFPH2UnWUJvr07GHkUv86j6CK4yWQB
/4IjYCDsbYHIe8q8TmUI4HU3wgh/VYtR8kK3q3CoC2s6oG2ee/gc3hfDUlTTXy0ZJ6LIfjWWsj/R
EIk6evU/mkLA/ZePHCkbr/pc0GX3FVqyAJOyn6bWzdR3UHX5m5ccXwaNaZQj3WD1wK/HGyedL9DW
/w15gJkHSXlD9Y8V3qU8qPSPVxMHeEZ56gvwUtUKEohm2G1nPp/AeBNFAmCtDNH7n7Kqkk6xdmhI
RtER+mvk/LhLJUg6byuCI/mPoOAWFoa6M3W1C/mlW9n7I4ZLsgZqBHkD2nHOFEPTj+2FnzQ0cm9Y
Uj8I2et+8gt0VBTVxysaJpU25duiDj8Kl1VzEWQeartN0YTOkCjHqK+BPqjAWz8/0rW1cGGde+lX
TL6Kbfas+l6ubI9jFavFxcVMEwt/x8vNk+sb2ZHqoHRz89LACiSul7n30uReVn1ZIqwqi5c/kFpS
0a8Gss9X64PpYN6SCmkTFafeT2apbwDfrtG8+jkH4JScFqAEUuKKYn4mKNw52ITME5yRfjYN4cer
ZzvnBW2kxfTK0zSbn1HNyHhgZtwpE0W5jMeY6LLmcpEKZaJUuvSls67r2wHk7IgcSjliB2zJsAgT
yz4pfu3UlZIxU7CjJh+JuDe6AFQSOKPstWFdscHUYld8wAle46odcfxJ0NCmCzZFzlgTRdV7/0Bj
KxvpLH/dyeFgSURjCaW9ZJYJFd2cCoPKWEng4HVQr7KMN5b0vKSQu5SU6yTTsnSnE5gn2euGmHSp
PP0M3taw60plLNvFjKB+Czd07DJOzCC8cpUZQ+WuI3tUEURfmoKJyhpa0uqofQLq7HiHX94Uslo9
BFblX+EtClAcq0LUkhMUpxcFJh+014zS6skwosjHQQqXijpr6mM0wkT6s6fQqQvbJ8+5DyObdn4c
fDpUIu6+16Ye6j5LHwDK/4ZB5+Yg59eqOJJGA2wI56u5Hq3H0BYMdrYJpx9eK+uNktkvIYOMVpBr
wfL3mHQrxDFPGj74ayBTcp1oxvmEF43+yfdNoZ/OgwzmKoqskSqtrDu0XLxsx7xXzMXO/SOJwBYe
oo6O92XXVMIgxvQ9h/w0CtmatlOttimABj0BBnT7PW98fGyFXr20NA5e/njd+/rAWKHXPRyYIg5c
dhFSsJpkzanbZB+V61fIluDwqvHD9ea3065nwCTsHfLzX/wxNSigHYXNbw84z1RLEc3tOAHTi08r
JlXJ2P8QbsLvGit9pRhRDgfIRVeFpohp2ItWIWvhX+GqWjjU05fwwOJrSSACbE9lJD5xQ4AMLaq8
k6HTOwg1YE1XIyjtKmLwyXDvGJjMeanEKexaUZ+tq6RW3lcmlK+Be9ISxrRIo2iTWg9l4pKMgYfW
kolZ0taJ2a3vBjmm4A/1brW5lD2k9HHJpiLhFn864/zVwmw+bJWEEHXF48gpoMMmb1ASQ9PDIMSo
bI4Bj6PUj9TOuifYEJ9VBxQ4DyjA1L7DHufCBb171RQbBlV5BT6HfT8eGROuI4Bc0CsP+tT+21ej
WAvyoTExoqDuo6nYXP+MpUDCws8zKZ4PBJpk/YfMCgBXI8JUUcKvXXTJUPi8aCRHu3tcLj3r68Qy
0zpHnVcBxthcM5ivPthDgLNgSj080nwRzWN4MoDm4htjxSMjU7nos5F0WRgkPivPEkjb607CB8W8
ClmFY26l8t42YiOAelZxm96pJ92MxAJcW+DhePfKVgQhXkeAW6vKsUj/RueIeLDYMT6WzhdFW5FE
KNcIF2dEYUbKhioWiFAg60AZaDoj8gU0WPEtQ11aST2971knShB/vyDMeosNNf+tZ5l6/RE6gUhZ
VQXPjklJphMhzOveIX15OcLa4LeJIU+A1bdQnP2Bnb7hdoTIUjQxLOiut2Gm1KT5TU3MGVZRs0Lo
X7em+hHW+Rw18YoUamf163tgy/L3+ehT/KXOQBs0iP/K86NDnL82lXb0npTrCFsHsykjx/y1rR0Q
H5o43bAHN9DYwGNpQ6EefoUcdi9xiGtdxv6OAOYKzHthq3VqlAZw5mylQgw3gLFxnDxieZsvfUeY
He92tKj1ZeLRibvzRh2UbRsBs8UlfioTdGjayY6VHV0JIN9Yrsgu65VZtzZCrGa/Wm3afjNRgDeT
C10c77777sOIUsgyUMEcb4qB66fQG7NucVy6hUul10vfUZwyj8OgU7rchfmKj/AptBxfsYxhK797
gFsIfiGhxEFsIS8YDVhIwyW6Ry2c1CfHezDMMQnz00a0xLF+GFYfrTLAlr3gm9nKk5y1Z2Nr4kld
S8v+TRTtsqzs1cTW9So4gowTpoDZCWaBfUXR0BeRjZH+xIAZzgPMqZw/tH5DU1lNa+3wDzjWy6yA
4mYAEFCPqSHDFlQYmK/v6RZ8ldfRcXtWvo6YfU5/g9eMj8Z6FXMEQU9XUbNKo1ZMDbjmrekkGeVu
TCKQmn10FU5oWDNyXKKLL/7LWdIBBUc2WLY08pNfHDW2v5aT9kR+ranZQOZTxL47dkT1ON7xREuB
8LBowoz8Cpxc1Q8u7D0Y4AQmsxxPtTCPuvzF+YoSv6/v/oZ8gUXNVZnPp9TfAAoXE82ka0TxfuYT
qJd4R7DbO8l9EQ/wcPj79W1LltuWKURWzXzsoKtah59ZruS6titVAy6l8JtGIP7zZm4SznUTvHjd
iQWnDtE9OnEs+tofQTnU5sn972PENPbU7qSYT6YYzs5ceoAgqn5xJtzbiLzMgs5gjW8tvq2u+zXM
AxHbSqRFs/XlPhTjGDPbR+MV+i1JlwrIa/deF9PlcCUC++q1c6nroLQanTWLKO1zoLy0huehlXUO
PPUR8kXMykzWnuFoPqUFdmy8flA67L89O82y99R65+k+4o7sPyv7Bow2gifagdM7lPx3rJTLbHiH
mttyzmgipLwbAKbB7RODtrpMnUda8WHt6/sDXbwgPjFuEQ44fSjw//yoIJJaQMlwuhm0GwKNAbaM
5aLiEJoOmDaLsc6HSUbF13dmXXD1+xKv/D5UMERIR8hEZXuzeFDwVMdVuaxI2px/kWVEfzjP1W3R
Tpt7h1Svgs9rMPVggUS0cQyWQrfhPCqKCk0P4DpQFet6OrYx68TIPW3eoQ9XXQfuFFrwF0ljLfkS
48aKxrtGP76FEqYg6ikvUx8IHA0E+wET3yAEPl6V2CJwViaWivCyjuIJKZXD8bm1doXT70nKtt0h
qDcpxk6smqYdpIzPO6YJCo7jM6RL+CZ8dnr6C5Uq+/603jHt3rMrRIN+x0osDA2Ke5moNK3UOdW3
iUCC4rzt69wYdsFJHwNzyPwpELGXlMugFgs54S7bkf3D3w6LBGwZ0sLroN/QRz/an8caqtdGr0+x
NXDMeADa0nNOp6jS+fz4EMMDv8EKKMvSgTjHE9m9Q/u0v+w3XH/HngyqeNa0qmUwD5V6f5M0crh1
GCCIAM5zKLO1v20CmpZAtEk+wFRUT25ZIIx+kZv6/LQMAbbLr3jg20fV4q0/JYAooA8oJzsjgICp
AT/bdwhrAi2ox7KAZjz6Eo+6vhf3Xic1a1qp7cWQa5jA0HEMFKyTsiyPW6fHo6L41G+QJkNDUDG3
7GZO1iGo+88vfQ9lUo5VIub7j6oRrk30xzNiV817uHbxC0ifmbU/WEdSO6s/rZrMjj24mtHAq5vT
boT7nw8wBjp77kD5VHRlwqHZMWCn7QGfODn0RjXoKApTYQEuBnIC6s0KvChrreVZKmjaxHDEA8cE
zHtNu96/Tu8SrVA74ga3b4x//Kdd1COb3/OM/H+/EFNVyNjQQpqjJrtgxPwoCwiN8oL9+FpcrQIJ
vdoF3WrWU5lXHpB+avRrCPP9C54xq5uZeWFHuxQMXNo25ySAYHgVhDA+2IXJlobK99mIo2+nObPt
tIG+BV8ZWYktXp3vMacMoZNsK/yuPp5lILEie2ac3AzThXV2TIp0NSi/WpEoG8Jj+HFosJuBZxBD
DBHCSWsCt73thUyrk/dwG5V3+LNKAzMZw56O4d2xXdAk1LoWw6JV71VGpZ6KZgT83bFwpkZgXKUY
B2Kmsqt9/iGD/1nFyZ/Od+EtfSUPqhPNXZeaEIHchYr40PeuZ5tH8/8vsH0SMqOM6LVMtTv1LOp3
jHYwDOKwkQop0z8xTKniVlbp1LM2zO1e09ETWa0JMoeK4KbdnSijEEVKrfyFjLyBP/RJm1Nm7Oc9
9YBbAytjOD8x9nLQ7Ubhal3x8UQMVEsY2JSLRngRLgI7jOtQoyv/zZCnHCan5wiVB+x2JluTYC0F
nTZZzGXvoTns0dqcdjJAoqmotzo9Sc8h8d6gJ6bq53rcknIYEqRfIRSgGanpreWMN2kg0xdiLuZU
sq2Lj5/EozVHIOXyQZzW7+X/WfpEEhl1Y6N8thMYWa5u7oYQT8c8yT2fgFHO4+PDfuLZ/4e5YUkE
G3IvWzwmgZ1M4j3mDDmD4ByM/6Lv/C8NI4wtLGiwxTc71fBm+hq39ewT0sWO3ctfr4luxdW40hlb
75NsMH+ILVP9CirWtFxU5r/tSD2ohLo5mFg/KM1IMPgYL6F0PTL1GnjJ0unSLPL9Z1dQa6hF6yAW
ZN11mTIoMq0AoMQRAP0vp0Clp5cSSrmQp3ubJE+Dt3I+hWla9maBo8IO80WOoEA4dlL05vY69+ZB
Oj5f/3tB9j4G49skWl8UnFvkl1gWoVBQtrxObcm7D+x7jU/2EOfilA1TMEp7F9mFt0lbNsQL+mxf
iOA5mB3qICvPN4LK2AIKUk6w32KVHEVOmCveu2S7WEXn4S69ed79cmPSlAfp7AwyIh7MsuSYOs50
hMf7OG4U/3i2iOJ0xl0B9YXa/PvG9JLtEzfl594obUoU2+UBh0np/W1ZqeGn0rKg3XsPh7QpwvMz
4DGfXCIYIWi1JK0WO+dHXaY2gDg5+/OFooiKvDYytJKE/fybvasijlCHKM/5OkHQmBskKIQ0jUX3
eaZ2v03mVZBJVZhuIHAxsTCFMuZC2WUzXXVuLlT95Nb8e8leRp2/Yhvsy6qWzFcPA07rhfqSK5sn
ExqAzxV/pX1DrbpAh95KeTukkU1CRC1EwQKdYF1ymH5i78Z3Q5ksiWXpVZHsJivJJYs58va0GlSi
bMyroUYK9B1DtT7HiKI9hnrl9W5qTNDY2AjdRTTUutMcL1fPBXg77B5Vr7Kmge20HtDv9YfTkVgK
CeM8uD8NW9MfmZ1AgHwDthAnx/6jbpFTQfpaHgrYW/NT6rYV10Rx0tx4/c6deHIdjJENJAifj3HC
FqS5lRN+EK0PRFht5tvghazsrYE4vwBfAf4d4fFJc6uyBXzMn7LWRzs642B7yOhwXeP7z5jnwM/F
tv60on9uRCs+5LVjxcEoxCga1lWbAAglKhMCiLuuTLhbredNYrulaYjNVzgOb4h+XuuKrJS9v9oG
HtbDIdBCWssLn6fmHQmVZFSmHtmNui9Tc3W/lEf3cveYXRIXD0Q+xJR9IbhLleYgeIR5T7L/QwM+
+fO53p08lP7yGV5eU/2iKU36+Py3h2b2T0qBLdj6Ks6J7cXHPZ6kYSkv/jAHagFHPgtKGov5xqck
W6ig6MAu6v3oXflUdhIVpQrGaLjljkMIKwk84px4G3gSltxMGqW4BsKxbNdt69okGxp0/vsZOgla
AKRiIRhiVkLqP006eXfPi2Lc7NAq3hKYUwFrzpRKIukfSFzsUuyzEjfKd7EmR+mrjBMwQgcq2XIJ
1bUW3m2mvEcuKvU35DTKR3T2frUQNoKgHovia7oDBIVq6V0MPZ4gF2glhI3MPJgd3wkXg3N0f1AP
1XTINvHe851UwKX+i5O15nevSyGLzpFUz6y8pV64hk1bHds8RerqSl9BRArFit4uG6VekjOszPQM
HMbT3Lx95ZrtiIZJ+kx+IIEtjjCcQYLiHRo05i5XAPLQcQI5ZDgP51P2hpbZueDW3yFQrXk+bkIe
BbWSSvgd1NLyaku6HWhpDHL2CicxB8Wa4QQZT+9tSEzFLMLdVauw9o98oiE84v7JYoYe84CCKKNB
guBelJs7uXZsednhGae55SJI/6hMXEapY6z8NW32Jg95DBCWz+Cp99mNXHnu8alkMPoNzcOVev1l
SMImEops2P5lNIq1S/7D8koDpWMWcP1kWfhJhPYkyHg1HMN1EbuX9VEaWDFphCOFa8/OnzSb5ze0
gXqw/HanoINHsA0Jv6NHiA/J/FM7xNX8Rj/TfGzX3RFPV2xQoYaFbe3utdTyBNiTOnZ7lJbH19e7
evS8rY84w49SVoRdon+c57EHn8twrKbVNzGcn2oYP1P/Ci5u6Dv0YK7QoglttggwA4+hFrNcOeuq
J8UASyL8keA4HW8+F9g0qIB7d8KyJ+xlvqqfdUAwVDlJnDjY9tZ9ZSDvnzoDm7eH4Fp+iE9JZaXE
apPDhmJ6uFUb/x3MpUnKM7LGFp6UdnRNBuklMtktOUyIEV2zx/Dx0Pl6CGMmnRQTNhOvmSsB/rjg
tQbEpCtav80Yw6MR8+nJmTZpyTpBa84Dxzyj5K2l1MJhBNO7lxZevAVxVJGxT3OBiNXzA1pN3R/v
PtEfjgNIDcsC9GokRMFOiAgG4vCw3HGmLtnurnra0d3BUp0D4DFstNw8lu4Z0alTpkvwOF72396g
B8NR7zLcELYU/QifkvjtwKJ2gZCmmjY9c5wUY6oIl1raqiIWKwbC8pLZa1XBs2i1Tz34B0oYcpXf
bXDWqKcDvTk0EOvKei/HIClXXMLi6Uh2HyVkPima1ObrqxvaINrSDHhoLRqT0QWiA8b0lkBD2+ay
XJpKAnaADOxGZqTUv1GON6U5Mi84ihatrgYFDj+ViqupphWcnUs/dXstjt2mAPAwyqM5mv93pHVP
mFHoMmrmO4CaCIiyQmxUR9sMuRE6XCCVFODFeWqHF0B7m4W3/xIXZkg+9LmLkl9gjZYKdAUoy3Di
Fj7JIs80VloTQZoQ1kp6eg6pB4ByzrUbSW2NW+Ell0crumqI5MWq8KKW7Y+9qy7fes5D5na/OAFU
CzI44rY77hqOxhT3tbDOSEdcnMu0L8vzwU8SrlIoCvrud3S3HDzwuwtAtQClIrr/tw+++TlQzSRv
WzS9WXPhRNAm8OCl3yERQjrr69EKx/+rKiaGQA7x67UXN6mkRrPHzfd0bh5kUkm9x6Cu4yVVqS+5
UovFg+D1nf6Bjm2nKIVUnpnYYZMH7xYXyAH9oOOFWjxfsjxQZe2qgbZHM1JXq7aU6Dv9sVG9qOav
CrqeKBOqLRgbWd7tjhMSIsLk82BZLM9FZ9JizH9Isese0TsetnyDmpkVG9ElDtTRmRZ6Ttk3I+Uu
SJR/2KWLOjRuF7wi+2Pdf9/6E2wsdO3uuWYVy9QuB6Q3G9l6CEuJMbJ3rqHl2ydKfdIGxIkQFMGs
krqTbxr+7xst4NbnbTf7qISgWBLkWJswcj5PQs8kCxE+92pG3KwlfPf6Y93bdOmgwUx5Xiaj+fCY
fTlXVgxklNcNjqBGId7yJnZhShTl0F/w5JJkaJz1BAxcVYuDliz+8nPM1of6BK2vhcyzFEoJAJf6
6KcsraJB6nmvL1qTBgWjzAADk8MQFgo5oTLdsiXOcSxU2/ouSHv03ewDRDqC+p8XjdlZb48rpQek
Fbk3uurbzwPe0qO2qTzxV4QD5yziiYIUMvRHLMnoM81Fav6Qg/7dzr8txoRzmicyktTqq6BUHMJT
4r095kLFuGs0KwtKm5nsZw4rmRbgFmTn0TD0ptduCKNoUecjmqxS5ePed23iOcRH0KTIqoZWnJ52
iLGQrGdvrc3lJqg0R/FxPixPmtNcmdsEYJESbtV+u9Pw6vSd+SiCevPF1iv//tmll6zgIrFeUEhl
tvqDYmloRlr6nf/gUGqbvvd0piC+MmrLWJR1xGRovwF0gKatcA4rple+CwnD9GjDhy3bfWvzGWSd
aeFs9oyxt8f1dHzKrOVp6fXQqPotUAsVfS9BePsJBVu8rfYgVpvFUMr6RbRpLM0rts/MHaNE1C3E
izjw7xvJuQqld7rK7aXrhML5yhwx/BqvTIQfUUH42SSb+L6y3Kid3na5JGUZDbA2ZUnKpdr/jkEp
TmEvqeVWcCUxRg6O0aCNpYnbq2FQWG7VhAvK2xvcPZSqdNAnQ+GPCGxdyUEShqOjwiDqkXB2Sey8
IE9S0EEY4LgEQbgk0p/bAa7oti2wRLzg9pkl8k2YogXn2anKBOpEoxb4qJgjZabJ1oEqt2/krtOu
vIXeSYBYABBZRhrR7GblHD26kHh/ZztlEnghnv4MnAdWaLij7jUMP18RnBs9jQRl9tuix65aXThZ
PrLlhzpATYv+ZpFJ+UGUiKipmEsAWIQu052B6njk1KW6FCoM2X+CBNiB9wS+Qo84NQr3BV2ID7Of
y08RErVk6zCqnIiaHl65h8cyChb1yvJw2bhTQqZMGNrZfMaw02opPNuPLutdTV7lT35oSP/BZC5W
f10SIL5ANpDCi3a2g3+D/oJrtZMylolaMDevHOxP/S4b+pxTkChdNFghLjHEq9k1yYWYOFZQarrc
n+vS+7qIrPoIXONBlEzTogn7HF2cCUX+hlTrgQAy3yiIl9NtChMx+IQFcMIT1JrdF92xjTIJhyYc
xPzdeSWJFbTlsHM36bA57Y46kRPn2PRCmyeBwIcp2KOXxgYreXFzFnrCPsX0KmtDffjg/iAqOrR0
R/bF/dgjg4RXm7m+OkNeixlOf8konxGM4lgK+dyfVJqTwqnNfokOAjf0v1dHB2AxCSBM4+rSvTvc
T1nSpHvDkeTxlxTcmZwVaHNfYGfpW9+pd8ia427SeysHe9xZer335NHSb5RJiZTjGN7ao1R8cxAB
HYxN+aj6re09rujpZyMrzEaW53dGDZCGl/s38yD7lOePn8pKpHdMHMo+mLoAGRDh2brfmxNlSaw3
dmoKN8DHxPYJ1Ly6dVjYgtHvfbUeQvgk4azf8jQRRyElnhtheUvyDAcqrKt8alyphVsCcFpEaDFt
X06eIoy66qF/T3Z/pWKHkUdRWKsFOGplXIxYxY1KijC8k6C1piGB7KsyT3VIfE3ll8APxCptlReG
W1xEKGNL4YVw0EoMJ/ou9B/b0s4RWPWujZfOZ4NfK8YEWYPOMv2NgMEl/s3ZX+oTtgkDbN8KEyU1
HyziEzovn4pBtonn6eyv5LhycXsNFLFrC0L+AOKLgD71gpX67OIaDVj9z7pSnkmtgh8N/CSco4y0
23fBNIUeFN6S3qd5/ZAMjNEip96/sAjmdnhcWll/AAA/wFcFFN01H2OReVUQxWo2fQo2k1oeJXya
9xZAXGlG6rzJC6p/keqDYT/P4CiHWpBgJoA0CUmcRIVamH+fX5TZ2hxMx35oKUtvpxc8jVxWd1Ue
QRbuadfTrjHm4LVYX5yDYkE78sKgK1LgFMSuT7CDd7g5K7hRgtorH3oxeQV8xzmnajQGnDc0MJ3M
isLWKZmJ/TTkLS5l6+vVQWhk2s31zLgGxHF9ikR4YC64iKcJmCy1COF6EGMWUDBBDq9UZ2G/t3f/
X0j8amL4xlrUwdjDe8qxElrNd76+5l9Be/08sg4LYUpwArJiQrNJhva9jwd/McS4dVdpzoegeYZx
dho0O7IcCr9JGL6Ldcho+t7ik3trq1oL6W79GzNyeviL/4A4FsOIs9f35FsKFfbCXCmV7R18t/p6
rIyKOIK+WkXLQyy0Wgu0NyYih7XC+vy3+fXUtlnhbiaiS4jR0HEC+1UGMx0WFzJZDfIi4L9j4toN
OyIghRJQw7wecxtLnKFeAgmYLHQpavs/KM6LwEBbiNCbqP1jO270IOGr3jWYrml0WHioQLo1eH+V
Yu5pokIYgSlIqIT1T36V2igRRsq6LiS82LLzO0CKc2HLlBRy1D/ccuLqu67JIcC/dmg5iJDPm8Ef
omB9+4xNRwYXvQtcFfV/6xjuWO7O50yGeCzgqI+mX6GC9n5wkWWZFCpnMkcnTYyh6jnPaA0gaBhE
joqbNGKaYRa4OU8BXbxIhhb1G51jy/j41K9qik/rsBcTNPQoqthGroxNK6mv/+wIj6mM2sZttJpf
WgiP2W2IskL0sQgZS/6udY1+amazp6l9xO7+KVtlzbuAamq5lHeLzCf9kLDDlHNN3NBDds8g+rLj
W79L3PvnBCu04mM4oNnExVQN9RH8fQS12omhBrlpAth0okIU8G9k942BZnjwBr/3XxU98Ofrwahe
Vi9VNJ4ENFfhaqs5nMWpDIhCgMH+GdRbGer1rM2o3Usl4rDZnz4VSrtr9nyjrkW8OGWcSNwguenN
qnBGQ+AZK8yzH2/FyiPZVxjRQyDBFpGm3d/UlttfBp3Sr6bpJ6OU9LC6F9XQmxazu4Rky4cBrQ7d
hywW4mbJXZv1t87MiNj4n0H4UpMFL8oJ0TvHsaomdByIzIJOd/ZYWtijkcDMWg7tKiY4wcAOGO84
wVLXrFzVmH+e8oqJZBrFQPRG1W3AzTqz62DivlqS/1OuWXsumQxUT4Hdqkdpd8akVBzWxsVs81Lp
hlHVz4ER2Vk+UkWNh/cySqfRGBd+4gCAq2/8yb0n1BItEZrtFCx5BP70GUzOg8Wn7yX1BhP4fYZe
TEZvbPfx2eQSlUwF4uULAWp3yzCNBnMg4b5TZ5w307SOV+5YFeoLJijgTayidzS2Lnr8IXylAGRG
Pb2/zrkx/vXu7FYjk0HJMEzgLGEKsp6lBKPVoEod+BQrDQVJFeAUw9q4VabMzVL8cUMwzRd0GuRJ
viW921IAkuW8cP5eMyYCP/P09bunKwqbPl0rErl/U4ulwfYyLMsFPyE8hBO4c8b508MxSzJMq4Lm
YiqP1Bowy/0Fav5w2wSqFrApEmoP3/0ISis9IiX+e4Sd3yJs6IecrI9ZyrFUdQhsNXTKBx0N3SZD
TRB04ECqDB2mXVgr7Lc9ECVeKnv3ow8AFRmiSfJxhRSFa8lxK0IFyWFcbONrV+TFTlMPOIRNOdKn
pf+6MF4SSl9ET5b0tvDKTAB6wj9cSgNsCCTwrieXngKw0sQ+lYC7tQ1qD66jYAKm4aVYU4qTKrXG
6KbUOo109JmOe/ib9IpCOw3oydlvq6f2RGOyxetFnnFNp1oAJv4Qi/h+AWCTM1GSXQkB0G2D2Dvl
Qc7G3vv6hnzL/HJmy3SziRJMftPpE7npnBSCv52bBA/schsXqgcu6KiX660lOloiO22XqT/OdmrT
8n5XT1ys2fCQ1z5ZJn/BTgoBRtqExgMmNzmGfkbX/YUdUH6ZKCY2ZeIeNXFTGlOuqT9R7lTS89Fq
mpctGvWCTmvGU+qAYBMgzIYcPuCBGkx2Pim7KVKLeaCfSM0htGZ4TbAW2vTSEgGY/HELTVOg70h9
F/BdBcGr2JrY95kK8F9iFxE9iH1dQMpzS8KHOufbv1VPKpl167neB399ZpikuUwlmRj4oeIu3BhK
N12600P2S07lQCiaPyz16CHhSS5gNnCBjxqYsOehmn3Ej0xFWPvaPTsWubAq/pRvqzpJqDsf1Q/X
ATAt98QNUeW3CmaCC1jdS23XVMqLLXGQVJ+D0tFMN0gTZOLWXdZPDgJzSj98qQuasGtd9nNkD3BU
t33LVaLLSfyNCisjkeYhr3pKAlOWzFZiPjl/44vcOyDBfEXDgTvefjF+9Nazsn/2yjAkeJ2/XJh0
0gGu1Vo1Bo4962sp10P1o3CgX1A27ReyNBFkTtkUAN4BxsOLAtzJ+gTcwOc0FeG688/bjT42oyEB
4P0hGLQt+Aq4GhRP1zbyYbvrBw6xLOh1AF6HQwZqb56d39PJ3DrPmnhJLhnkZq+K4vDYvIvZ9wfB
oDpI7Ysls4mcr9EFnDxjOGuX/pIGFqzp9wMyBFqbzspn4BZVZv4Xe/oubU9nwtNRHEIZPdCBuN4V
+WlnLSMIzgd9UyreGhuwNwOOwo9KyB9asblI+S5CC7PFSab8zfDpaixsuZGEFLKx4uD6xlKUVoGY
G69YdSYAzI4xK+V9j5MMgghmf2E5I2TaYx3CtxZ/l1pcf/8aa8MytQiOlDJADYpr5523UB8J5VgV
TXoiMhbfgVDwBRrcdM8kaSUKX3czZKNjZ+JllSBep5jBkl3C0MobQIo+KjSy/ydpQoDAQv4ftNvT
i/HIP5G5ZxmB8VL8ZOZdrp6QHyclutrkQHZLaJtRBSIaLcwwZ/Prn6i2BFkFBlM8pD8wAWLHE0vh
5EYy5swJRseF1WU0oTPyK09fBYgUqeg+GdokkwhZrj6DQQ9Hjh3GCtgxySUQmlUW3DLMdylcO625
FVpzxgNhP9J4Ppal/dAUMarc4Khh4mjzeSmgsgaEGeRp66BORwTeFnw0v5BUeto47xs2or0dzyFj
wL7ywnvIB55B3uY4LJMHhmlRGqOMDHCgCcbzqM4hfMQbDVeUTevi/ZpgXLrLQS8PkY13e+oQGqYK
YAfHc9TS+eGRoOxhguijx6gbEM72bxH8nGh0RqyrH1iyDKO+JjQpyv9aMATP+m7svJgzf87BFmAm
4s0kJxzLx1F6Z6OGULij1xpdITS8xIb35krGZN6Z0U005rOv4gCO3BbzkKFJY4QHAWaONO08U2+7
lozegZWirwW8QMMRZz0GoXRZ04LxC+ldQaodSuW3YHfF6oauCYYhm/76g5juvPvUDo+r4xd5JZaf
rrprnphG+XAEpGSxmgwB+48fZBb1UhetzjUlQ3K0lQR/VgwoJ0YHCvQt+D7Q3wgJ8kZ1BhrjWYPh
p2AOIAf8X7X9VJj5pkOAc/s4HPX7Ca4P3LWoSlpnVW4puDjgiDjbAQvKm7ck9ScIEIHDak++vcDH
3qQYCMnxh5/mqFK8MR1efwOYchxbSyT10YBKcKlsDHI2nRni77zUmzaQO05AEDWiGinfVGvuzv+z
8SZRCmHwKyRyLl2on5ZhaktCX87gtYjyU517iIEnm5XvIR4JqjgZkIUSNLETcJsbaftMdZX2UqXb
Eyiy/WC1zTyCS8+/AKPheI2FJVaI38h+vMlphPcprLDY+KTwaZnSIrD+pWepMrBi09Zd+McPeE7o
uROBD+hQds8JQztuFODdnyNN7HsbrRj6hXtTDBkWBenslaxJ24utqQ2NJZ0721lVw/SrEl4jGGfz
4Ous8QaWCZvTDJcJ57YWIQqHzQB8/258nVfJvzGmcqRkQChW+sR2ghmKpSnPKpo5dLoNC7sJ0N2Z
yMCj9q/2/giml36v2rACvR9G+ruhb6ezvOBPGogqQeMqQF5RpSoECn52uhdwv+NnqN6/q+IN7Yyv
F/Lw/1tKhsfQBc9WiZOw01F3MoIuffQ4RFGE7cRuI91zi/j47kWlYR2aU+4jOjpTmGc9a2JtCUOI
/KdgEZj+1U94kxpftY8AV8dUY0jvK7NxfV/+2Ql51sbZMRmeWFEz9zemVHjioFkT3kNZg0gU7JKh
oiwjr39zBiTZ1qN7E/NcX5OM91qVy/F2Ltl2vrzXdB6Apz2woeEq2UlngKjnkgjOapnc0Tge+SRi
j7cKsZUqWiMxM8PmpWxBP8jRN/USG5iKIhJ9qeVZHW0BbUjfpNtzCo0B0VJzZl/XB760niRib3BV
bWmSyzLSM1xKLZtQRtYR1bjoVuFmiXNfH5zO5Yo9lVUUQ94/hkdK4XNGM1PPtJPbfRqYIBZUhHAa
toauvjgIO9ZmHNubvWNmH+75BkPRcfv6jNQFY3b15MwR7b6bktcf7m2hXhqpUzAa2r9E+lRKQn8j
vMy+cs2GZ9JH+RaLBi1iOtFlPrtnv+0yKSp1qghPAtFsmK/iQ43CArJVypcQ9d9oAT7zXgmtr1+3
d2mP/gzfUVFbGnxSeTiFfh5f+VagD2ru0E6LFeB/3X4nX2Dig4iZT6uLIOHnOcYf905PDSTZo+WQ
VCObKUMES01YsIZDU+ck81Yu6tf7nW6mBi/YOkZ7xqYcUL6XoQpRIQOmyNzsiaifeiXEVtj9sMWL
DbH1p63wffqItan/j/bD5CwHzT/phMs+IWkNLxNjmZj40vel5fVPir38Hy+kP28vuJ1Q5yVklz5i
NstpsWVUzki3GOj9zdBQJfVlHb3gzb7/EQyG+NqrcYJoeAOxhcJ77FsPgn1F0Z7uceF/QcDllmRj
WIcT50osn2wwYKYrvSXucdPXu2s78NdSgkxNCepV0K6BcV/tJxhPQCQGyF5zVl57p4lP5ZYQQiMx
54hCy898+MMtz7GUkOn46RQtlOsfw00HiOKbGXFCXGzAofPEbkuWA8QqoMZMcrsk98pISkP45c09
TeB+c75/QzMOgz9D0LuyUiU+zJEmIkkCEW9vPXfL//p/GMPNygnzx4csdc3QHbr7yogO0eSuCk+6
rxCN6yzYxo449N7KZWavtFYJSRaNA2ScM34BJ99robYcmaEcNuNfvsmWaX83VE3I7bngglmz7KF3
fhzVE4AsWwgda4K6ji6lDHRB2H3kau3LAU1mGlY+JIskrgj3eKTf3vXguUTKEcXtL6HaICDpew5W
MqwO45InLasUq2VA5GpLqI8uZDTR/7XK73IyjZ3XidKcf31jkvbfMOJGfMb8+Sf9KwUr7HfljiLM
GaW6ogU5FJSYE8b19QbOd0Vu8TYmDcdEHrDGoKIOiJN452ppaBZC5NJPvUBhaV3RqOL7VlNeO8Ey
JV6PRTvOTirI7DItoBy81tH1BuieOg2YvX5UrqAnUp036nq2sHYeZzthh5bdszc2TDHRYVwbocgl
E0ldwAu4vHUfFh9q+JkVd4eWejJuX9y/0tFA09Jw58kI5vD1pMhaP+t0X27t6+6dmz6M1Ja7Sbtz
Xty7R32ZyDInaUn3wXRM4GA/vat0vJ7b2WyE3u8ez9derRfgO+kLpurk4F41Utcj5hiuewwWm/5c
qXebtUzTAQCJ3J5Yf/idGwiEN3Q8XIQDkIiuhdZMdqPGLSF9Kg5qV5tMw/eS/4FDJhLk0aLJmfuN
YZ5cBhPzXqtwFNiq/2j7CB/fJkbCkmalpnrbXCg4l0aOjR48PclGs9MDNf1UHyvyyf8ceL2FGew4
4xVD+7f8iawL4S+2aivDNurgWBG9wgBlhxf6NNMmvTx8y11mas7w0G0nUrUr0sYKK5T5uZIT820l
nGYdqe2wSgv/gca/DdiKxfWtNp3K7z0L9K36Bty35MjzpbE3vX7Mr/OdrIvwYtONwONcEyoTi84A
7vGZxA4IHZRDgxtwVdv8fozAZuadmRUokgzOxm1AXRxUqHOx3NPI0412FhtXdtrMs2H23eF/CFsE
3npArPLTQhYUkWQ4YAQtA6rxElHs9eyoZte8tnUxdwdYCk1xyWDG7wk4y2k0WBT/ca0KeHV4nqDb
fjDVSE4y9qDtvP9lACrKPHyNmGI5d69bViog6pLw2zVBDacuUCVwDVfOp8+4m7Am5mdUcFBRNd8i
l63YjsjUkObb1jg9DanEa0b53wJIT4vFXCbC+Y316X2pPShopn/LtbhjszY/tH1BTdz8gQeUwr1N
2wp4ok0hot1cXPO7rrkkO08YC8F2aOmVKQ1bkbA4VGPVe48sYZyJ0c5beSbAVPR7DAKpjuXQ7/ff
1CxF3+QwOpdwhvGlJ/y+trNK7Ste0AlyxCf+BI8bGBFWatfimR02f59kIPsbvg7JfVQukaoIKt4P
F6lVtC3mfjlX0NTjfYvuyV/UB0Ix3HWUHVagAXdJej7hujBwcTbMxnk9c/hzdPi9YDSXIe21jlyY
uGbJOfF2LopPZQdT2gdtMQ6YdTVYxGq8hZVCkNHaQcSQAx4r13W1Pui729taix/coCgMeWDseEcC
OwG6y/1It/uYjWa+bCiiHbErTobE4YcF+klPHXMBA0kuzIfxwMxI7s1exXqkCDNyj3hd3cjp1TuJ
xTw76SeNcecxDqQ+Z2x6f+UaqEPZZU/b0EEd3emPRLeozhyf/4Jp3wgcxn1BpS5VQKZuXdNZ8M/0
LcBE2qtlcj50pGYXKnjSPXue2B6Ov+QvXDm/5Ku79m27SDsvrDq1q5f5puc3cAPqju+xMFVrm+zt
MJi+eLjQhdMSalg/DVcRdbP6Jj3wlMLI35/0E5CUIBc5w6exPoc0h4J4y9ADSCNg/uBTSa4qn1dj
TaLTeMnaR4ciCuj6zNTZCsB2Z4oWKYxlDPJ5o2OMXe29FfeG6oqRiRUa4vAngtkESHsKiaN+mK3e
IMynibbOe4QDD5PCrB2Aq0eIixSLe+bUm2h8UzKrHmw92Db3WYmVfMwJKYEhqcJsfLmbWuCtroIt
UUwWdjbAeJSiIDiigDQwG96vI8/DqX1JLy+C5QBR1hzV9JVPUH/8e1XFde5ZMUqhclE8rAHsjCUX
8SFAtjEcAoAMQd+EqKUyKmSC8IDxA+tDu2kK75Mbuevx3AeAZGa1lbKgzaUXWXKW1C5OUm578gzc
ew0k77AqG8u1KRU1q9lLYuFQXht1Td/mbCM+ujKaoZFaZG2eMh2Ytlli5nmuxXXlyeF02MS+vc1z
3GLIyDNkBZ42201WY7rDhCDy5b1TynbuLzggH9TDvWhEnXSckZjjiXZRx6A5CoUD5Oa79E+0s3Xq
uKLghw60kTYhnUSl05OhuOHPzwUZDGML7TxvV3CuFgRzfbbYKKWf1PKc/EoqWcFZx/w6mSZREr4C
7rf3wwV1tyJ9+JhR6Os5aUAsqcZ0dM0iFFSRPyySjLFhkg9L80BA6dsTQno+TQ+X6/aHt6zloWH/
WHZkFRLMTSnjP6N3PkOoKvSrJqfSzkVV3A0qQq9Ob/Mh6PVAgpwtPUu8M8+R6zLxP+HzbYP42VYe
w6VqGo+5uHFCpprhfTZJJgsZI3dA//UscFr85ct0CDEzN+vmgT6JgOo9QPQRwp6qSRJzsDJatl/F
dJGwocfE2/48Wz+vg0Pbc/lzUComxBaPVxtbh+wI9TeK9zDB5DqnZUFrWhkEK7KCK/pqE5HWccQ0
hTEqeoCFQGetLgZZN8teYcIitS3mUqoLs8fihIxD1giMinfpVMSdAuEQ27QhkG3HSOXOAE8nymNr
rfPE62aSZ4OHiHtTZRJ5toBDyiZgx4q1Vt4bXE+TRPh1JhlEXswvyu+4n9u7o0GLFHUvlQB0Q/+k
zO0fekX6K91NAHzLTIGxIth+rIQHdgeyKFP4bpevRiEcZpDdLINAM/OeDfxpcMXGAiMkkc+DsEC3
cR3X7k5GlUysq4xI4CXE6iNp/bxvlU3jCZQBrUUHye7mwiJr2gy8tQ14pxVDQ7FIMdpOhvL9TeDH
OA0JX4iofLUAI/Pn9ivx7yMZhvxQbAJGwYtnv7Y+3r5Z7H5rRkDxuq0Ii3KrX59RBVgcJ0w7eXNx
FkqoeAx2ngA50OTuhftIAi+IZzVtnTLlUXn3/Mu4y0EVwStCR9/u/R1VO8C424mTf+KF97ZfKjCz
zROIJbFr+zpaDdIdOQO+2gHur6FiEepJbJMY1WdNaA90ybmIGBk4okCfZ7AEI0M9m+EOv+8goXxK
DSbGo2JXq94ehW7yL8EvaRkcjanTFKKCu9V4uxfr3ytcbGF/EDGZv+zKFDGG5L2HWCkkqxAAUnck
nXpHKg9HdzsVgdk5hbSsKRzY3JrBRICzOlOTQymJihqKmucz8iVGMiUiKydAVLyFV5BqZX5s0b5l
8cX3fQ45ASevjs8VCwW4o201BQapN2cac/tCEN3tvLfBA9RvZ2EEcFBkr8yXCMaq1DTjlXVnR0sU
dvwoVeDtnASA42GmtoYA5cPouFbVBW/HMOsUSQ9+C9/WJuMFOCPB8X/0CNt3HK9f7kSgAZiLSiSu
Rk3oDzOOgiaHVFpTomnXWAuvycu11BGzfOvRVasXkHdIVBcxjM5GI/plqhztQu/mH9rxIDYS0IFh
4syGPjSIDVtDFBCCxNnI4m2e2KmwfMJO/dkceVPCU6icFgHS1q+cI5PYD9IRy1JqEBoxCCVvCiWY
k8q3B333NzcpemCx2OEv2N7AoT1/XYf4aGGZF8H6YJFl+prfkUtWUrMwY3L2Y5wUePMloO1FVWZe
528Qj2UamsSz7iX/tPZXg9YnqtTZ8zznzEviE4yZT2Oqcab20XYN2lY0CwhGxM199ySxKHJAOHRK
2i+MsCZus/5w6GXqORX31YQPPMOWxtksO417BVN09Smikb9tcnxr4Xfqx2gnMU8IX10jnnq9F1OH
NQiz9pnWLgiu3HFrlSyVXoSmUkST8/4PR/KwylWCWbUK/29NhGXBu+y+ZkqS65MmXLJUJC585lYu
s1E3APbYN8FAnZmO+FrgpJqt2P2SHUFSBGe7z8uq2FBSWRmDcHc3zcxofVVQmlEXWa1woa5cMoQ1
/BTZU5NHOh/SxTtiekjXe1xos4Gz1+dl+TaZX4vLyzT2bk1Uopt3BU4EsbmCoxfE0ZXfRYvPsYwn
/EjDvTW5oeYfUVOCGA4cXN+gkg4OHJJzdm4MR1rMDbPmmT/bLjFppRaCvCsLPRnoUzI0AjWU5OO6
lM9L40jAlU8Bno3zDbvapVhImRHothWYpmY7tVFjLQBfYut93iH3x288B5IjMaXt5tvkaIrP8E/p
u4RKkzGiHnVC8KcRf7hRIhd89MHcOnvTeV2Xw9EQcrU8+OvLJYmPpApsWYePoEzgKS3a9tCn4qjj
KtoHX76SXE8fyf8bet51+MuPWpnFvd+ZORSS/duc7BVCnjPEgifWrnd67zGFPrptygLKNUwBeu+5
Fw1i9haqe1CnZ7ExK+gQy4FqLl9bjVDkXXxOh/QTEyAnKcs5XGCamR6hUzmf4qM42Aki5oVnqnXC
TAFWhdZn3OKG69tdmrCtCEN+SsoUoqOx2BjF5h+9wDQ75Y9qFxbJcjtBmNpXnJWsqrydjR8LIJRH
MFhaNZ4xDp/tOlr4oaaAb5x1jrhaAnLCZqLhQbOKX6ODIVjBb5AOV8EMy5iyukz72VHpn7MgCxwB
+7xDtpRHSalu8t/XhyHB8u0tiD9qPSwTfi6/7Vu5B4wvjv27onca6cBpBEHzCiZJ2rCr63qsBOps
vgJicIkdNqAcoI6JIvZhO1LGia8gAFKJj9eXRM+LTV3OkbwhdVD1mqeyuA9MFVA38ZyH6/dcRm04
iVLPexbSqwSxLB0IreLHvvXI4rEgF0kR7sHJW6qTbM8QGWk2RxyaY3P5tFT4C7qnOiqBfoF0Fwut
3xIWdiUNRl9lXeP3lpcB13eNlowhQwIFdtcsGEB9pIA3FIK2IAaVzCHPsNmPmqm7pu6rh4yM0gZz
/4eT5YmYBD6PYU2qW/8jjWj37JQsHUv45rKCZA/OdmzIoqjT440hcvSaQG8tBJ09tpKQVxfKGO+0
uXX/cPrNKHwP42SqbTICcTuNU7nArIbUafWbEzTxxxVWI0LThz2pq+WwLTWQ7zhU1zZBIdKsxIHR
tm/qYlLw0uloE5/AZUVGaeRup6IQehKcG4NgoJPmkvbWRlHDLctobZ7wUj2JnoYQ7XElEQfM2bLJ
d0gD0nN59eZSpDv9yh/n0TEk8Nm+iviOoKtpDf8UYq+CumotUGsWWbVbnxXs1cLS5GT6qbyORL7F
ZYUdeCWoPsDgJ0/h8ZNU9xSg7S1/ab16ek2dg2msxT58C8pS/em+hvUq7E9id+R4Oh725+ATRQzN
/12E0mJXpF1QmIy76quowuW35dKFIIhUb79A/WmMF5Uz8M4if5xKruSROapEhEVXLUnbqrqaSlVQ
0PBVPrcnYm2Xx3LRGLeaORjl4avM/N0eFKcJeMl3DS9mi4B4a3mGZxmVlM96D5H0i7CSxUldtcmK
dVeChWo925fq0nsmk8sinSljstLA1+w9MlJo8sRG+H65l08GmfaPP+2g3IX+vHSFBZvhe+WsAyI8
HP7Aq0PqoIcqBB5KZcqIEmUr0pAtkesbdbDUadDXNjDFxn0AVPi09Q40iuNn5MQkjWOOsZIRSUqM
xy3LepViDStk5zYt9GIYmUx5PTRdpzPYQomxioRkOKawzh8AGd3CdwM1X9Fzu6JOV3joQyO/Pdij
4XEHz6DeUEgtxeJ0Z4WHbDY2iCaSVaUkDId/hFuhhM1FBRLrz1U/VBYaavZ0MjDKTK0d0CJLPUsZ
rPBuOEQ/6+H9B9UK8NIVr4Zsf9pj/oEppAw0uqUM1bM/lXoqwkhbhmONUVVdRf4r5ppbdfgMfCuS
7ZSAA/TXozHPDDx6dFJg4mUmIbb4TNW3FBDUL6qxgQREOPgXsSaac8mPZ+FXM8IjmKFMOIztHULc
ekk2caxN1FhMtnLX67J8CdaX8BzXO9BSzOytgXgRA6fjV0GF+uNuGd9P50Udq1s+ggPDQTH/csQz
6joypAvtc8D3rhffpeYWim39VHGFn8cT/ORLZRK7+AICBW4tOXp6t0puNbRuceqp9WJ90h0zYQsv
iSu2QEHTTxJV+zOqxKDbz1HU7A3PtbZ1dueogkGSeQ3tXCpvQxvcjJxPqGROVHA97FkxZBxfTO84
e4Oa/GuIqmyeQBRTGs3OoQiOho5Iciekp68cKVFPEH1yeEePcnRfW8j3hdO0XWUZZTMtXLjixoYr
JiOY4VUnjbk0y0jCCiG7TwFvOSG2rADH4qUBpQ2zLq43l1KT42YhSkHAC5veAZZdlAV1/ClePtfH
t3GUyYO9Ta3Z9xldFnRW0x8e0F6Ho9Id8z4SJJlfdV6SZW31fVcOABDyKZfWMCfpA6vjrsTS7KWo
QNG9wLtpdAyEjsl1GJS/UfjmeM6HI0tTzjCfE+v5xfhr85XtMg8Kd7BtL6rhOSemqCJ1HdLUlh+Y
p0V7Wa3Mwyby4RdrtI6TG/9ub4ln+WH9GxvLnoD94xfwkb+v2+PdKnglkGwujT8yQ17OMEixQAlf
FBGt8Ppg8VoF3auOw3+B6usq66riIUx1EbgrtfnVQHyZRhzBLPSLalTH706ZTP7qW7EpvZrhJDtu
dHiPoWcIWHvCyagG593+AiEKJsOwJWJpo0banwF/BpwYkKZ5ETePi7vTUmGafwQ9limsAiIS8bAp
6tICNDIELE5PpUbzb+xY5/0ea363avH6Stn00lLY3rU3srKTiJrv4kFYkbxxW1TbuqLzHShk6v15
UZEyLwYpGAMX/SrxWn3dEomHWLxR0RpM5alLM5c2/bGucg3PaJwcXrmiu3uZob8HXR8PkiZ5NkgK
PeLriz+LGttjS9mIrKQk83vU/bBkHfPEV7PJHezuk6CtRDVTEN5tNN8Pr4MQYA2WBsrdHO5JNNoa
wzoD+jy7liOsvl9HmBI5JFy+P0R8EHC5CZtS47BMKyX48fH0KU9MyZmBCkuLo4T9N7z1YX9ayMKY
obKqMURVHhFDptL3x+6spE5KYQd5Il7/5fGXTieX9p+aPjYf4J3ncUjS2l6y1MDpywazoIWRK9rW
7ibKxSO+RmT7XJ4mbvDmCzY6TwKUjKR6MCm550cC0/fE2U+EQS7+7NiTDOlzFozqHw3kxFVFGP1R
PXsOZ/bRFoD5AG3nCniGBAk9M7T5nXopVuaDcoCa4Hb184L3Zqun0mt05Cgk/Wa9WnVFwSk/DjTl
AXzVzOcJ164BhM581iRuaeJe132ZDGAGEwsy2ukU9Cd/ncZS/6BqJqTaq0rOwG6PweF0x0TowlF5
rKZHh0aWiB3WJq+ZyccUG3wIszTlI5U3CD8XELwE/15HCr4XViU85DxrKLXHtVHvjwuaUjLs+fA2
JKKp95T90QaUgTqgGE38ZBMzeXwwceDyFkmlNnCXrvYTXAKPln4V28JQZrKKWutaqf/SMZcblQpc
MgPYoSWyDK+BvPojcTDBCLaq+CodrGbDlPlr8Sqr7CSYqWcQbwJMp4fK3kBg/O/Cvg10vZNDjk6a
oBeRn9j79V0+CZF2qotDaI8xzArjOdmbVLOxGGXoT1cxIMT5L6bqTYWGwnZL61A9qVTX029kgXg+
SKNivMAq/lWZEkGyhzTxWzOAvkx9hhfiDQOqGgAgu2Io+PvLoCAwYaMrQ38Bc8rVKQn/RvsovZCt
DcPN091eaTz/4ih3GNLJVMj6Vj1Wrtr7Cev68ITaGZYCqYuniB8fXBCfRjUGtmTdi05dhsJZFEDm
uM2FRjJqjCXh99WXatHd2UkIr691wEBDeS65NzdpMjgjm5ZGfQx8tGikcjIiG0thTAaWDk1iNZb9
56Wp9wGDMpEQ77ZsYdo/7YQUoz0zPDux5eK0kJxlEZe5yvN2L6gyrqqyyqjpoh8hu2Ju09v+UBJn
UkCQWnETcwsUdq++F8YG/T9jVJTxzkPEs9qjlRBVZDMkFxowT0I1pvmcK/aa6N28BGiXC45P4Jtk
J19T2IBkyUlAynidcf0HGu2jPjj1pDQo+r4DP2hGoNf4ctEa6yktDeLvCKHecEyL2diQ5rY0KWGl
H0Zhkrjq//yxGfoAT3L3sb80MZSxDhmbJ5MV/l5TLP9BnHJuwYNADhTuMlw7EHErMRIjiO4aslpb
UTCp0rmY2rgIUyIZrqHgv4OHojv3JHxWSL5GXA1/bC7tDEqHpAzb8UU2oDu8ShSygtub8GOTJpZB
VCziT23OV8PRtvYD7drXVdzkKSbCdTiB7SdU7UuJ7vxSjz1o/fPZ+zZUjiJP9X4QFwh+FHjQMrW0
Omx42ObY4QYUv1X8oUe5QsJy24gk1Q0DvQBqUmVxoOHV9t5TSRIIyH1hUWfCuotK1b6C6hrTx/Cy
GT01EgMhS8cVIRFhWvOVwj54SoNXRLatcpXp2tIQ1YyQ0+SLDjwniylVYjN8z9yYB+deMoR0BOQf
cXkBL9VrV225hc+3DfBQklz9OV1tDJQuVDXlwb+8dS3ck3/uPYdhzzL+szvtRak214w6XfICxdBY
cfV82nt+D2mQ+UveADvVeQ7S81yfuzjV+cAuPhYpIOlWPeP1Ns2tQ2W6NsquEK6jYvfNJ/2cJHqL
KgNOq9yOhc/NMdOAj9ST3xAU/FVvwAmT8qmnIYXdit0NJEVLKMHdh/OG0WWdhrgENGRExe7KBcqJ
+GEKc6Z53HCoz6dcliO8+bkz6YUdVnJa99g8o+go6mxoEBjuJChSqz5wlEEoYVi0uyFa1T+GANxw
fTHpJ818coC4JorBj30zX9JoQhqNrJB32jj62sT1T/K6GBpGoHzOYKIFigqsYBwRV2TRbVUuglu7
itOWiNq9JfdUDSDp5k3tUn6qF+N5DFyIIFfijbJmEcrDVr/O1Qhl4HT/LMODirz5DB5gNpF5FiyL
0nvJWTkJkeKScKIscYb2PkdPi9Nzdd4UmO0vsAd2+UXSRnti9uBHPb3ixxOvzedOHnupkJE9PgEl
gUlKb14UJnUrBZgVig36wqrjNS/Ji2WKkG/5lB2AcESNPJxs+YxwVwK6xe3y3XquGQRlAEgyzMud
30ZDMrv/twLyeSpeEjlGN0Ag4snsKIgja8obad3bRz0zF+0rz+RvCGfy4WmvCyzAHYm+r/yiqQQj
p9C+pM5ziGPU5HlqzlzL31KTK6FnDQFcSon3SG8g4AQsbs+4A4bzrvaFVFKPNhIPWJ2XDf0VS33p
Zt0ci1Uq0JmqjLw3rautLJFEF3j8ey8OiaJbniLVEVCjS9hdPjYLgxWum+K3uFEXdGo3/mM5oiI1
l0LKi0r4+gjRAgqU5O/VPjxr+ZhtcDkHdgrZfd3EeKELUrmXPS0uuROWN3X5KnHzbAta4vjHV9PM
NpZtWnDYZABQ1iyEAxPTnKdgOQ2jF3uDrUyfdKopj+No7LZEq4aYu55aqNDwXV2q8PGOmpZwvFrh
GAAjpALQNfkBrCQVQKOdbEtAT36RYJ2YXgbq/yU5qeXImPPc7Ijk5PtpE3MdR8DsT/wiC6VrlPn9
Nrp2jC9fwpyp2jFOJd2Yu/o7GfITavSIDd9x0DDhS5Mm1dAhSA/6DDJsFkN6tR5nYUgU3lbe0xTm
PJzRWZWo0vN2foMw3xVRmmkSkx+PisQ5f4o2xfAkRjDzD9BKOcDUGY5WToZfLb3zc+Hga77m6Lp2
gzN4DmfJQwMgoMd/TZYsJpA5/qDinkn7Qg/cxUiRF0hkiieIWPgMOr+toRzUg2zcwesTPZA3+wr3
FjTkvrAklYHGaKHSeuFQSMmTxPJ2yMQ4w0zgLW1DqxJrEIw0gZ4x7kKy2RjsfwNjs7QosOesPK+o
Gn4QqOgiP3H5wQsKNIu8g/bxgJlEyhdbQyR3LVCG2JT2SYm6aWm2M7U/6GtOmrl9EFbmiGsardx1
PXH7/7NUxTV4ACnmbSMLxoj1QZmE5DRu2NzaqLoeI0GjN2nda2Roewo4MUzQpn1F3pFtnl60Ztwd
oP1XkSeWt4LBWHfsieA6fHhu25LA7BVNyqpQqmDPacZYIvzLEd/Z3Hix914HJog0ZUCFasiGM014
RDXV6Er5gezOrnlrXWaHIxRKuiOkgzF3b3EimRdYcllbDHp+pWvUA6MSHdv+dDAQpgGGVMVucCFX
rmpSCvQiaiZ1+N0EeCnzVmmxvyFns/vwPLz3qq1FPxl4gEYSkwJ7fw6jjQ3yMxD0RKMkDS6yvjCQ
GOta89E2/u2URgqmBF+C1UOm8tYid6byxpWvhm+7RnlmrofhMj5YvHbE8zj5n8+N3JFef+Fl3sRb
Ae/80F2Z5SU1PJjJMDISp1Qo8pd/JmqZlwuBXlmAzMOAQjKqMynI8v8E4SoCHnmKSfWVUMbfyYzo
h0YK0vjkxQgvxb0FPXxbFO0ZtPJqpM9Ngz6Wwe+aeHIQhsKqTfvMDyZ2SSLKW1LOu3GukwmC+eYI
aRylkvnfq+sErbrMjp/3gp0jOSpgPtDASYMAWYQgg6Wpo84pLAwgo8SBaMK7vrx4T99iHDorji1H
JYMsAnpjvB1wrALEjM7xAYVPRkNqSYgUEJla4QADMSe1a+zxzmyYSVJjl7XMX49pd9KbckghxdAS
buCcczkZWl8O2T7RHW0SpdfXgOFRnQE2L5KuVNvuJqCaDHrh2lm8OwLr+quxPUt4KdHv5hNBmP57
UjTRU/BYjuu7XcBx2QbvVaKT6gfNP2PlP+WczQIAW0yZFPXdOtdpRWDBnbtvsbIrGjicxWHOeXem
wfDKWAqLsTlAejxDB8T5xNBy0GuX1y8tQ2Rvw9GNqP+SXPltXIWYxYVYjIKRwwXgJq3dAi7Yn7aK
1dzW+oS9X9JegX5WxDhOodnJjaKKkMDqWYSQE9NwYR7iGoXk9Kp8o5c3spgXksARZ3ykSxB5MvqZ
j1cMqhvuXpVOtsuHt0goqU/FMCGfxkty/DPwRt6t4ZcK7mzbAcmpUNLXAUNVj/+LEVsYEG+6zkZC
lTlBEw3hq/Fryj3EiY3ozPqn3z7GAjr2uDajqCSEMMniuS0APXUd6hdmkAae21cjPpa1PGhN3N0I
N3fsQzpVLgr+sisqxd4jjTaLX8eq0fWjd0mEm9+RAAvmRG24XJmBWR9DLdc8FqeKFSnqm73t1Idi
hSELXf6zDpTpRdFMq2l2JLF2OhjNZbjJVMKvKlirEwe0pFb4dTDYocufeGekP1XAN9dD2ILU9vqm
Z3M5ik8tg+t114DfC43vARZmNB+oCDz9sbMmn+wiW1FaFPxmUMqboNDcDkV9EZoTcAEDdkgf1SKK
d5Ap6wNzC31KXM5LUY5rTLh0XMk++zpW4vVnIuyu06Svh975nAUJ3xrxt7U5d5hOOKQhQurlaSl8
D8DkWiQifKcBpzLKARoEFkvctTUc8aCiLHzPDvqkCv4BoU+EfqOqutpzP3fhPn8UhB3dWPkclsX+
e22GOoO0WPQVwOsy8WbW7jRMhBZAbLAwXxY5X9BqMbx65p/Z2JuRKzqfYAIZEI2tbGGTYUT5+K+0
dRgrSlkH/kzTcZNOmcojXcLOeDWPSC7hH/Cr0VDdjVEuYitG4CdU0wvIfRoEHkKg6MH+iPTyTdas
bjHtGBF1z+bZc/KW6qIj4udJH85gM96zEWkSzBw+wksGlLrQLw1yxLzHZ8P5pk4vjBW87YoJaBo7
762tkuYoSMsipZHWKbbJSa4nv7vCmtwi3Z0QaMHPJFk/LB8pNkwR7K1QtpQDlWGv8P2lC+xNgaYf
wrIDBYvwfOibCnGUSQCPl4KK3U8NbJqprJzYkR4g3yPGX8yvnS8CpiI46PKHXmONFp5xzfPso4L0
3v2UMlzvAEjgxm60/kOOyOs0hTK3gwl+QfLrXIvO3OTj/0nEeEPYcG3zr2L16VMi6GWz9y44BJAI
lqD5HPtIkil8/YurjQDA7VIArxlUM0Yuxr+tC+KqBmcDok6WvFq9asMxXpFSnreEnabTWxk5QxSB
fNwZ+uRNmbTGWwH5G8vsBwRDgunwj67gNywBZGYWDnnB+N7YwnSoAAnWcJ1ANylCs/yWeRoFao7+
bKizkd7UKVyIGjMkE7mZgq5frIAz1WX1jcSPdaNH4wC564zrMQx8s31RZtK13oWLPTpA/VeV5KrV
vEq00ONm7BTwV811nGwMjRbKu9uma2fleg3NoKjZGegHCvRZM6fpmIPkyw7Ad2Lro9ww3F9apj5/
8O6x2SutpcdeyMJFN9jW94ucGwe/YUBhclXzfkGa+7CN4WB9SZUg9AZwhSx5s+2OmBvZaR3Wo4lu
uFY002A+NtAt51AT+J2Oz5A5Sq/3SLPlCYQcfWweowUTi58F6xNkYZweWmgOH4grZwHS4MsfvdEb
PmvPjX/gXA8SNWJMSHnaJgAEGNMmIxb16n45g4mZg5c6I9xVHvSc8xW3S11kPBY/1J5PAuq56yR3
eRIQW7h5k6oW3NwVsgpcDmyXmcbW3mkIGmeGaTr1YJ2GeS2Jn0ov4PzPGtVehgTGNHBr9LwOacE7
dSlWcOwbFNxyJt0Hc1yafh9itFYu5p9CuYGt9Uj/GCleGg3n4zTBVqR/5ZGaNwpqTa+CV2xOig/5
CKqmk4Wix8B9qT043eV1y9rVldLsDq3Up2zy9wfIjniXhykh76oA002Izs2peOgyFzCbKAur8H4F
MohcEO7Ha1UTu/mFfm5NL9sEwcGFcF12GYDVp/6wg+VwdYA5lcYeFiWtTTwgtGnP5TwbSn7LNHtf
b7IyXbN13/F5lmlsu/ZJZYIJlS3fuLzh/unYbfPGRWaQ2EXuFUr3QXsdy5f/q+MRcWGPF73ncgAr
q1lJFMBuKCKy+GC/ol5Y3IYEOPGnJ9STA6yd7i6xmwT2pum2d13wdEptUpIzyUam/6MoC+K8Ps2K
LxQE9hna69ncWOlW5g+Tj/LCeudc02UBqhEdycLI9kuyRPkS/SJyxYOlokBPdQdv6UxsJTmDr5g6
+/gw2bKGapCA2rrwGvv16smIIdeH4UY8fzOD5sBZe/HzS2tzWmhHCl8CZbX2tnMEmN/0yzsHehSt
jHki/qkhBc6qpLBXBqbbetgUqWHtKUADoodY4OeCn9L6m7EdEiEmpsiGRzUmN/B7CQ8NxV5Qlizr
as3VqWOXSKXZi2pE8lvboPcRBfKq9VTKE+ZsXpCZIMJyH8kbukmaLpQjO8E1Vi3Add9rBnYyMgEa
cpp3EgJQtQysh0seg5KcIeAIEcLB9JFssEjxH3aCXQUY5KMJS/aL/6huXW0LqIRHwnFyb7iYwgXn
4+3ujAzMRfO4M+2KmXv/4GQ2OjzgLq+o6Ajp/Rm6nWh7oUlG4ZL6HGxRClWf6dooBC1ayJN2aonK
3BZi74+fE8SNkm92JaKDAasbgs6kP5jrqFhYEGdtYqP6IMD9vTFiNKufuvt1RGqgReWHg13loZ/d
OUeoe2mfjQBAuo6vmQyQYDyUu9pLRiI+EgtGM0ZOCZtkgaWWX0HZofeobzGk7S6VOdTzNPd6hgnU
6TMCKuHkH0GVe/SlW+oULE5l+OBLjwsFoJEZ7TWu5bgM2/eqwW2CsNeNhENIYVfjHgxRc535fTy/
TGfYHkK4iZnW3DthAizxLBrh+Exdvc77RNGzM3UAVdSBZCXQxz8X5SaO9ril8jNpo8ScUE5dZipN
MMofj0i+x2LFY8nHXg5rrg28WVG+lzDo6D9achdiDnn4ilxI/xgxuopWrg7y5gsJlygVBAjBGbM8
L0F2oEPjOQ0SXXOnBqhgr8iyzyOY9vj8z5fQsQh5rhKLlqmV2klyH1SmsLaN+XUo99WOO7RweSI4
wcyPhY231BgJdNt9K0/hY0G9GXZHelzVi4h35h09MX8zQ8t1nVqA9KfKGU2r5nPoht0KxJsu9vb1
xg0/MGr0uyzcGRfFrySk4WgwAwyXHWywhPy+igUveBBOWLJ+sw9iWqbcm2hAqWloJkq23OgnLP0i
/67UwfZEwQGF2C2KdjVbnd4ER8Qzbf7UOAW0+xVgNeEWvt+FGI0FdDoCG84+a9gnzScNiVF8N3zx
CPtVYqyDaORvyVlZkH5xiUuTaQpxgkujao9WkEWGOQjiRXujTBe2ImsOGfT5knvIrGMCCdH3nOKA
w7fQQwEIKLGAlLVKcTXjg3ZwUZWBdpzpr2KcApl5mKTlUopY48NBfqiPf6q2z3/q9+V3zGUC3Q+q
+eH2wTCSmr08nE2zz1acVI7tZXEA0T7QkA2NybCmTcciViCHb1S9ECVHL/lUMOvvdKWrg7uIG2PM
y59+kyNNpqepABtLoAdB6JpD6CFZOh8Pg1dseUCnCmy8zgPNFhwa4mFXMSST/TXTSdXJsYtxP0lh
WIW7K8lxXZ/DAvacne0FLXLe85STYS8QYvS2ivsl135gstgONfAfPFzy77d6cbcqiBwEBNRMtFuw
wg+E1g8qWguMtTq0wZCSz/ByU2c5bse6sWkAHYlTcccCLSHCvS8Xwv9fJTgqWIAmyrcmgbzK6T4v
ZQPfrT/WrIhvEfw/VuJLo3veQ+BHpjQP8+3kCGQAOFakXZ6DIcC/PePxEL12N0/waIbSCamYHIOY
XFpI1/D6zC9E8/1hVvZteuVlAmkNimLGoMdwRAkGSgKRzzbid+oXF5n8+zDMwgMvm6CzmcTEY2bt
JluM9udMlaQEuU9aym3srHjyT/kbyVYCLu/ds5W2TB8vjn+mNbWFYwT6P+cBgh1s3jRltKUvnLPb
AhRRTeovnd2A+p3ttxPwzTNts9UjSwa8kHXzQG9X1GErzRE1iRGpKyuRZF8VTiAuN3oSN/2UCcZu
zIFAbGYzcyBnk730dnWQX66a+lZYScMK3IeP9x6RzU/BDgux5CuEM8GCTgREXHaKwvsYD1ckkB1o
CGKFq6kNyxKuE6IKm9I7G+wTxb/cb72BWSemtJyKPNrK6c6ZsQKTj2/1rqcfIdIWnbWAkEHVjrGn
/k1STwUzMFUYPt78/HqGBUqO3UqnVm2FYogl6ihSdPstpgx8C1jTSHjotUL1QLaTGPvE3P9BejJO
BQ3QIiyr8be3P7eYpIYujFJ/+06fKP7IYPWUQmAcHtolfn0swtjO5IuaCcif0xHjiscIOZkmh4Tb
LVii1xWdjNrb2j6hn7lXg7wFyWDbU155oJ9MA6l7F+UnLwRNKeVEidZ61E6QLzRykZ0KwsafNJx4
N5VkmkOyR3bSU4Ch8Qrl4kJPHf8PLckQgq0UtGgkxOXE12M7oXRTuVAH0f8/caSW0tk7DhHTECW8
YYRudzwFS89U0t2Obm93XG0/YJgmm9z0Q431RL/I1bHV9gxY3yftyx2v9SwurGbu70Mwqw7l3P/A
FIj/waL7WRj/M4yDoWLcedqljVVMSGxLV1CUxq4BcYXygLTR9qyj96fHqaOtCx2TeUIe2PbjUlpS
qUNbGVY3qMzKUCqUiv/rYheRsm65dfLc+h1XV0SYM5YKBaQd70F5t2bHFzFR1A0CyV3thA+uLHzE
YOTuf9ib2ifHcL5qieGqt8udywKOGxccLrT9ZL6yP4qjLuW+WiBHonPaVbTG8fA4QoUzgjba4iLb
dpfc+To1fjgbLQIlNRn3FPAn/G6QvtpztsEYmfXGgJ2MgyTSQTSJIsuyONAAASvC5yew3rDLRPFP
Fbugh7MaWVR46rGs0Ua4j1H6HC0L3Ofx5gOehOZhGTOUyFouXBM71Drv+e4ado6m+Om57xUUb3S2
Vqo3sPRkTz3EprALnBSSSu/xVFEiTaAV+YrmK5RnqBJlepp8Ldwe7Whngnlk0OxJfESOd4dlhP7o
6/MkcmdIau/5JaKLbwO7DMNjsiH2byl8YDb8m+ULnyowfgjZEdHjDbvv8PScU8a3ANO0w6gVoI5k
lyhdSJ74esb9BfDovZ/uUu2X9oC8oVYMHicfZ74HxhBNMwLJIGPjFuN8KwwBHNDrUpipn2cv2zh3
scZP5PUryZPTNYw1z5ndZEhwcIeeF15rFXt6n4WMxG/PK9ad/bJ8EQxtyoWFYeqAGSLVMEp376qa
uTZDH/RVkV7PMuYazSjpTg7+cWERHizraiyiUp4UVBzFgMcJaY7Fx/2EY3PDdEQE26w26FKves63
NUH9fqoONIH6kFWi75+sPzU4KJOg9ZiodaYAqjZPLNoXW4FiplmMcDQFzBaAkC8Adl+7GBCp5RVa
V65/9g5zo1xdY1JdFE2+mnO+8NL6n/UEL7VUQYxg5Ls0JxldH99B+FYY52TDQUleDQ1Iu/gj7FW5
75NKO72LhdPIgyiTf13ZR9L6iGV3iip9TxseHurxMyFcN8Nann2HHGj6N/R/DkWufWgiURZ4Y++y
/H320rYrY6b9oxzJjYoaO8grGKKDmSxN9yKByNPVx5ijvQiFOYQWpK+IAqZ8EiLwJKmMTZu42z2O
7AAY9wLfcS2iZRB/krvsgfmVuLtOwpUmkO1cR7vIxZVFIwEA+vGuYGBN37bA7xhM6yeMF6wErbUr
tHrX/Qt5h3/oIQddhvORC4Xhpjt38pNarycYH000W3cHvAGeoViv0yUErsxD5ikN+iWmFDdJe8UM
kujouFfUqAG0eskdUiWDymSAr0D5hpKzPwO4h33niRA8Z3ICuJ/cVD50q/Cz+iAtIyqvBLutv6mV
KNlobTFfTh2Gy9TaLv2Nxps0+R3vzWt2AMqj47Da+AMSHVIte4rzoYjn+7amOp9YUt9yUuY4bgqD
dvuBx8w5pjxoiEpGAtocZlJDCAz53E9Vuo30CsIufvuZIO4J7GNH7o11VdNs6bgwZR25g+c5+kbz
Z583LHmJu+ZlRG2fduLHU8QjdJWJTUf+8Y/o4iYKJOeMQ+NvEiTgaYt9GldAVLb4eGrrlrge6L3h
IpfDAecJoOoXZSmisQPAxOT4xF9SMeJMYPI7PmARggRrh26BUXlHYeuGbW9ETAsC0EcPjY/ebVvY
xmha492IWzNbFm4jVhP4PYKMO2wpThYBNNOeTB4aQh+VN+pvsY19th8yTFl0OVG8TCV6kraZP8/c
vrvdwrD0JxWBFpGnpUn9Q5cYSVGSysPM+tjHeC92kuiZbtfr9renUBYgqUqAHnTZwC0Awoyafoie
O88DpgkkH6cwa/dlYD2NtbHB6fRQF2+k8kynPmsr9wqRFgHPoS78okzxRUMYALHecNoA/cHUP8GR
GIxO6CW/vXRe1zysA4FMVfQNKPruqaBvwM2m2l/CdX6zAkRhR5TY53atI4BPJrEkd/ztis4d0Abb
V08SNOabTGuVbj79T3whWXLTYyTy1mLBSuzSvN1xxZZZ4fwD05pK3mjynmZfj9+EpCYdUzhDKA+q
vGGWUbJNlxQqJ0e5uGb6on7pWhBo8+CJHm8aSs2Ezac8j8WQRXTNFjuwY/CyqdiC0Iz0QtIQ+yFc
vMArHUw5pGyhoqc51GwF6pp66UfoQSgi4FI67cs7p5qwr9BVfyzwZd7Kv2oOUVelpqxTLpoyq8yO
PWakqGG2EwzRrs4qVPuW5SHZt0CaWY+dcwAjXRhBYFJlLwQh9mGNFWhNRP4QMcEr9wTs1Ra7Yk4d
mt6tAnkONAWIc5VGLS7UlK4bfC3KAxs5HAqN0H4O2MS0a1+ob6spLTAuIXqjl5TsY73Lw0gQVBrE
1Q+TarYhKQD8LyzjEaXgM/Evh/wnFOJLsExV9KuTtwtIF98RxVqJjNE2KIZ0WDD3wW4KH0y/N5PK
4jY+A3siE0jaHXfTxkWvvNC7CiV+bEf0Bw9qCPm6mWdDkXGl/jdtaTiQ3DjPFoq0ltAksAhRhpln
Atts9325Z21lL/7dhHDB2flDawyn1bRW5YPAxR2EdHn4IXdsypYc66dVM2bLRnG8bFVqqlnBtWvw
vR8GO4d+CL6td4F1lNnrt5yP2MVi/OFLdnnaJJRbqehUVNTEJA6cf7Ig4VyYym6QgMJKBaooKrOe
ljeGGqLvYSfKASS6nG+SxWIQWWd6ZEqB2gWrfSJFXMr+OomRivyot2a8bLXJ04FWwb8YUsnE7o+x
n120PEg+k1NriJ14ie0Uzqi+WpPwOF3nI2afkElMfZC0mcjtGI/CxmOyiZvXEJTLsiUCQ24vMdcw
0GJPkWAXMXcPvfZiuaYeZXPvdWm241w4MZUY2rvKPgR+jxrnz+3Tpprw5+x4hzZ74oS97xOG5Xbk
E1RZqeCOF9DeA5lQDjF9UoYgYChd+8BX2HMvjyTEa682pRvtE8E8/Tk64nPzOCwwTtihsRmd8IOa
YpCChwjc2rXePUF3QkPXDV2n21YJIH9TkbCH6Y1QopEQ3IZM76b6vn5nquyPniicNQGru1WpU1kk
2JHOzgWnKuKJSjBIMjoKWEMgdjO7S/C2wUWr7wJvKx85MTILfcPMuvlhbo9qNDOZaRf05GYL7MCW
X+TbGspQ7o1rjqTATCjgYu01TBL+QObTxDsEks5HZkHk0J97Ism3tCpbMP0Asljxr2ctSqPFr+k4
ZBnDh3qPnKYlZNaJHQ/lcSZiWc+MXNiFLXSZ9w/gELDlM2DbpNb8JU5YSzG3rrRFU3mXdJ9hAzgI
Z3t8L8RS/JoQrXzEh0Nj/2DuuvzFh55h/8BFPrhwjAuoB5qGNx4kdM5oYHGBU8DfUbWYAfTRBkZn
4FycFuY/4N+YFFQBP8tCDiNYX7VwirQr0O60O9cT4aK9anroRRAA93Tzy0VtAYaqQR2tKDr5Gi45
iHEn1QaF+eDlKnaiYK7RRK8rciUULhFRs7vghrlYeTQ+ar2iaHD5LD1kJFCk4ZUy0VS4VSIEyZx5
8aHJxL751QuTfU5zW4yZsi3f7nsUv/tZzCz1JjFPOw40GhBz46h5LJeji7Iatlqf5hNviFGoEhbZ
E3UA9g3/ZhSOStVL5Q66HRuBkyBxVoZEkTHfxhZsAqAwaKqSP4kROzkm0VVwjVcWAyBBR2rHL8r2
vVVswITCH8AzfqrltG4QuzFlamWBqC9FfN+xOydsTBYHTof4Lo+I12dnVGLtAc3AYVUeLp7SWJpB
lB6+VnX9jAEEwxl/x3/OZgLaSnbmZwUZo5X2Bw3eIsxizFC3EPO47nrsnfcIEzvkoCvmJ1wBEgU7
evsKVvE2YeVIpDKf6oRJuiBV9ebUofWVwpjjBQGMTpl+S1DajfBy3JeKdA7tmyqnqU38BgSSjjhI
zZy1bbf1zvaVrXOYFlTbXyOC4pdg+7Wlh/QOjtmfv5WMv9EON5jddgegfGy3n+4aaa/FgJIpLOGg
dSOdMbIkfi8a3kYB5lUdD7OyKeKDt50+97MmrVCOcFFLFzZEZMj3keJ/UHznADCdo7SvqgBbZp1+
n+WUwDSgJMzeiGj0Ya00gcipRhz2UTM4jGfuJCvhZERYcfveGlgwtmo2A47YMZqxC0JDJWdVElCE
iieGLM2SQAnYHAbpvk2hdwAmcFQBCrPy41POPEiW3Xv+/9XxoN1ywMnt6luXJplaX/Vg4CQZbaQl
Jz1s6AsP4xmKxqolS8gQzO83EzyULvAac07IhLtzgRwpILBwvQnHt9v6EghsFZbJu5tqnQ4j9DZV
MrQvgAIP9FV1FcMzd4+CjjtYOEiyx2hxHaAxRCIsTT1uIbm+dedjwYibsyD4/afoyKuhiGYYUlZ/
hoRKDxFPmpWBKFwbrHeCQowpMFDs0vc10u0ExEyVwgtMWMpuvAG+QkirObsIB3lPaKtgOOewJoZG
WyYBrfzk6BLybfEVTVPJ46iJME6+gcsY3a3cuJxGD0huumoYjgVqyuDPsxOqGfFunZ8/hKd1i/wi
4wxVGEjzqk0bkDElJKmajTJxf05ou87/cVCatCe29gBE8B3pUKjQFEZ8hYtQ8/k3c/obeKL5Qycj
B3qMtn96ql3ZE36q/+9Kk8TzE0/BF6onS29byiuvFGu/psKbutZkjRI6dXi6axai9BKVCsuSqKfB
3h2bZnL9mvtMewqC2RSu7PkqiIYxXD1wG5TMKWevLj8mjSa7FYFt8C8KLMrOgAnNNKpr5L+j0Sh7
oelDyHH1lzOYwSA0uQXQMzsnxaz3wJPkAd3MCajb8g9Mzdl9fF29DXITvTUlj6qzlAWkDBk0E5UQ
0E0H5IC2cdaZsjfkSmp40shEeJ6ob3rxOZwVJWV+NY92076ce47U8xikTKTUQFBCOedU9cUmcvLD
i40qIFT6sXkf93N53WKAk7zLOPh3MFh3zxoLiJIi8AyuGRv+41O6f7bhgOUwQl5VaNT892P/y7G0
WUQ1hXCGnf5VBxXjChATqpeCkWHC8Qr6b3o0SEDAGgP0mMmyq45UtF2eCdE+JLUsXHZQolXOH4yE
qDsDT3viVffpPHWfOGQY2S1YLnhKavtkzFYkvagcwwXzqimdP0scdvgU6YKWuHuqLQfwBTLHcYiK
fspEJxe6OrIlSCR8LPUBmlV67THRvp2NvEgrW3jKZIZV0FqTCP4G1kngsqfOs2o+z1bLd6xafvH3
KKYe1YFIU4qh+4b+UFSNAxBV0aWZWHEA3f5/Wpokm86fnHVdbggU0wLWbOBIrLliCloSGbEsPPbk
K3cTE4jr4bkwvgZmqOlmjQ7i6YujWRIVYP7DrkS8lYpiH7B3HbKUJMGf/O867qly2/pdl8nAlZbz
a0EXWPb8Cuzv3W7rQFTnHHXo5I68kETAt6NBeHO23zlL5OkUtiV/TOrVm2t7yDJwiHsvw9EqNrjz
BGQceQLaszMTe/bHYZujkvUeuoopXrVK1FZ5ySawZWZjQk+VpLzPwESr0I6d8V1TMVdF7HyE5KiD
MousdELkrIFXyiQ9gnIWb9nM7Ka+GUIxvIHo4dHUVxGriErg3smLLC4VBFxP0NSZqCf4V7RvGbV2
197eN4mobVZwnjiN4RDK+ksVixGY+ZzSJ3cf3Czmkiv9gEuQhloyx/ghFlYn6ba964C/ITnT5+Xf
Y7FM2n/pzgOektyUlTFCx55s8OBhEMzQs3FNac3hPQxERURBwWjwMUmGgIRl4fiVBwEBBdshY77D
fQnzf3BJTMqOVPxK5ubKPSm+ySBidYTFK0Ckd8kdDvFraQFUVTYNksT24OWOrkN+Cjd1CpXu1YlK
qqzg5hV5uONPRCRt1XDWNXDuUROM8kjinO7vZpUq+/jH/TxgOBoHRssP9qIvK/WwcPUSjjCqoCY3
a6VytuuITZau4dt6MVG5hxbS+ubWiw0wp6Ma5e3GyuISohRChWio2RKXeJU0Qge/1BBXYZVJmNDv
HeYfw/+1nFmo6u02WQWptLve8y3UW6EUbgHfMtnABxuX+/vg/JHNlqa021jlBvrnHpY2D+xfikev
8LnD/2qnT8irdstA9hx1UFdmEhqAmqgYS41PKkQ3QB9IHYRidvaNL3XX71aqpqjnZM75UjKEbwkQ
HVHrmv+cu5hkJW1rRZZxzbSgkhTvaLiAac/SRpjHR6/8AvqPh5e78N2JdeO6qm3CaQWh5z/levA0
Fvvx+PsPWiF+RtEyYLaRvzL8Gse6L2GqZqUmhANBwwdD2CcEIM4ovTqrs6XLuwzO5vBXMs6t2ew0
2SaEZC+tnfKTZwdep670NDibfjvL8gNKzgCMT4wDxVlqBl11H8O5QdzMfbrx9YVdHjTWswFbRbRG
7HRNvb+gWrY7sFn5BRtGgfFV/4Ih69xQOmuDtytCkfT19y2XFTkajCvLuv13+7zGKBlE03QgwTVx
7wTnnjWJc2cKeSxj7/I03Qw6NOhuWjZxkaywJ8Rt1msfOJPoKI/7J2sWc5GLKfkdspAoyHazIAGH
8BYci1h9QrFEmNe83LRSi9IGMnppq9HmhCGS2A7S2TODj6rx/qm29HHvqd1ANXVxq9cn6H48GhbH
avf2GI4JmhfzRq5MzX+rPlbBNLqANn8zVPFFQbSvlBZ8A679pc5KABrIHrQBdScK0dc4riTN0U1U
VoxRGCn4bd2DP6dIbL/IeCYGqU8YSBh/clegh8C7sgcglOsOhFIZgcV9imwlf+b5KgEFwsf1WYls
EjjydxKuNRL3hHgzlParsbXvtkrlzaDUDcR5m1uO6Q00xTnPrgNgxk88un4sGMsI57ZgenFR2c4l
HRAnwFUVEjfJGMbrFYU8DC9Sa6RDR0KxF0dHz2fH5jJjiMNpdmvX/I77j0HRDcdpxRio5YK/VSDc
Nc01e9pehxhCkb5+4VrZDBRnFs4n9I9gQe50Cv16Q1pbZxewIrtzEfS7bYxZXn0wxbleffHUaPTE
vvCN+2KNMTotezUBWtoeO2ra5pBqvW392A3fa6BpcWXnp0Ju/P3NatKcipcMgwmmY17580/pDYp1
QxfEiDrcT7y+4a21R6e9841QX4n8YZ9p2hr3DMUY8ZELYcpAZwqkAl8jkktejtDsMNZpaFWr1dZn
Du6okUK5WGUU4cfJvqnj8ulf0C9ybbFwiYP6zb+3SHrvE6jAVnGsKB7z4vqOOLyIMGtbUAGepS/v
LBMB8jU+ReLqem1YoZ5fddsnbHZMrMDaLxFCIqExFOfWEzfyMA9JtsWWehByMXrryAV6he1KpX5j
aqeWqMdEzEeWxFiW+0u/LwzkF4yvVfc9ThYbgoMlEXVuzZIIgU3cdz4H4SORbL2x9bqduayVzRDG
WIUjMRKTE013LO9qu5y5SPHdjSBp/+7oBWMwj5peUXxZoG3hLrUvucSlNz5/nquXtoJsH37Hz2yP
I6/BacW4X10NV0ET5WuL9P6EldyAZK67YBpHE8LV2JtgkD2LF6nCI205GHdl/fAWXSxabsqNlbCF
7XE47UkIQLiSIhZttq/TO5wE4BaHkOfeA332qYJRLcAekS6BAwaj02leiSZRqqaJw1uNdyTw/ems
vlZRPW+OuHqQRTs/fOgoQuddf9BfcRwyUnc8piB++/d22XZlUVKEKtnFd5sfW15CvV0JNvG5XnAY
VQ3J4EUA1Jz235T5WCIEBRr58R8gyL572pxu82Pk1Sw0t6sMLxqFI/g2rvGuu3194cOr3yJH2BGg
VRgcNQmT3Q3LzY+RqEjtDFerJmQtPmd6bz38vC76Dl6zkHxJe9aVXpr6Pjej0f9Xr529OYPE2POy
xdLdV8vTEODHXEmiDxpLDO6Bp7HpT1VtOtkPVwcac5P52BFFwiboTl4JBX/4cOaaFW7pj2a2jlCd
3QeOesfVewY7Yy7jy4yvocMBoXVC7Z6wiuopmP9qkvUZLH0dDoo/7orfymDk1CjgarkfCC9Jlg/y
e1EcLZi56WDYkDWmmtuKYNc48s3v2XpAgUuArRzqoGQFtTy69uMzbZOVRWdwb2DndfNfWfn3/RZp
p6tCXjpX/kHf1RwgqrcdIMPFNL95KzJ11mH/YxJxGYc3VLYHOKKCXcHijmHlMNn/8rWzT5dhLbHN
8bHu3ejmz3eD6plqydRKES6Z0nA9dBEX7Aj9MEQTB87ZVqyLxBe98izk48P0ZO82WGQMDX0gXM2U
gO+BHG0CnD3CKXjD/+PNnrd+hgDUep5wTPbS28zFc8RhyhkSyh2btNEeCn3mltn7UXyKpT67W0yU
JugCjcyuElglcj0eAq5SjlYcy87g032m6P3gAEEbKH6DymNZ31UohacNzPX3/Y38XkzK01SjfZhV
H6C9q0UJYbob9rbVw+M71WHZN28in7P+rJz5pB2D+4AW3kiq/PUoZQBDFK9O7RbUKXVCJxO9jpOx
mh4AcsVRR+no5JtLbissnkTkd03LYghvwy9M5jlwo5J0cocZAxggxB0Bqw3lu0bTdfNN5mhsRzmD
bQB5Up1J/GMZ9xS6q7qEQoZxGdCYuH+YWjicGD05AO/TjEheTLDnduuefyh1DCl6ZCEDml47ufdQ
/n9wpuweDRRF41jSelGPgVGQIG9NA8ugamxx5b3ewSPnFsQCn8IKYtWJLIZ8EvFrl0N62CFzPMPy
7PprYCAOpM+gU002dF/q4N9gwyZqaMx9VfIqQgdB0A+aLN22KA6/Cr6rGmD1e4pClFcdaKRT8FES
tSbFY79J+OEpPDqPyDqbwKNyV89+rBoOwQbEokosw6jX92QHz0N+iX58LdLCykls4mLz354f4bEM
pOYvzrzsgfW4KawCgYMBVMwRdTyS09kItz3K1ttvbHOGDV1FjIy1XHFP61QN1JnrYx7li3HyFOvT
4zO4eRL6/O8JbTYwNUojJSWl8htx/1OuqNjrzQmu5HTVTEuvrUhm54aYpcH6X89MRxiD+w+bjctZ
ZJn4j+ejTf4BMMNAhR3XyREMl+GWc50QW2EQ9mT1cueN7HZX2OtSOc2Pn2BxCESgPq8GDGfyu3CD
cD89VUJTCT5OaOuUZ8jB2WJuvJJ/6lwhjxhTQ6B93HOLM3zUaUdp6L9uijTVh1nRmFYFI65stJVB
c4mpODmaAtUKAx6CkV9KuBzf/wd8tW4PdWJmw9lsqsIlMhJIzLJFYSiUI/42ofxqk2ZzDOq1H9iq
DswCMlQfidU201usMmY2V1bi0cMtErvPZgm+BD928VZpIYeHScLIFlfbEecxxAy3MVw21VWuT0Pi
+P9luJDdKZBHoyxxHOKxBsTNUAQW9+2oO47EWBsKSbRVZyBnA8hAGLaV2S5dcgNfl5dAfhXbxUo8
2HVPGNzvo/xwLXlGhJ778u6C2X4NkR0TL+oq6ottWSv0CCAIbbQSMaHbfugDC8Re0PKGzOPQRn0R
Ub/5MGvvaBXNt934+mwi4qrJZalcrRsjpr6dge/oYIMLrOVa6GvsxWqsyWwlCoB+mPc00OP/X/AI
KgRztKWwTPO1NGuXOOJAZaoFX6r76TSyDwYXATrnyVIWrmKeNAU+hjLP6jofMxsU8Xc6lSxxICwe
PXNKZET//t+wYdGQjyfmylqXAzB83AhJyf/mlVcJak2t2kD7SyI7oYz8WMIMAITG7AfFFTCnzocq
L6VHryDbFTHW/1jL6G4o2o3mqvgDNs20E2PoqR+ZEIyUmdLhhP6XVnMyNjxD8Fnh5YCnQKh4DCgP
nqVudrIU08BMa3FEOt6vRiN3VsZPCJZAV+kJcRsy9MiF5b883N9Foz85T1LOehSnxD/HCE8g5rwE
yi2k/DkiJUmVKe/7nszZbBrkyyaPgStxzYcdVsW+YWCmDnRACUNZxHRzBuUkeL9+WR48WlGKmu1M
w2cc6V5E/kbwo5LVBlmsdUucmgNCoq/R0ffNmxrQcA6X03UM5LiY8L6JsY3RhjHas6rhsBQX8CfF
iaX5OzXWn3FOMzFqLV4oTF2EA8owXxoMJFqY3ff75IDaMU4x4Kq9x9cFOqYQ5xAJnA4NWym73aAr
z7l7uaO4FZgAjk+U3mbbkbB/MP1DusarAExQYNmpKdnJgrEDDomz8+CtocM3UcmbjTtFVDuZlmO3
jFltxKlWDaxElbC/C3iLumWruQ6sVlee7R+BzvQxsaQKuhwPr9/rJ339fQ2LX7jgWsXkX3JDIf/H
4+7Z285rtozw/jElJ74SbmAZr7OfWJlkkxEoLOJkbKo3DWVqNKA94UGicWUdzbk0UTFLC4AoFX3C
ZQMW1uXYZ2duuL5r1ATycGHuOgj7EgwAzuzQqOeniDgIDQgsMDkrUwGQ/RupGrBU+9ndGUhnRPZa
xX/qCqVR11u8FRWhhpiGlTa4cSFBo4SOFaRch6aE6ETOqhCZ0SGLUF28i3N86aHiRH7X+8fxbwSM
Nei29VjF3izp0qzKb5kYiF4RmJoDeaSZFyIVy47ulJIXYiMlGqB47jC2q/KgYRNrz9SEYnLl1Jxb
3kr1aC0hIQf7GJlUg+JJ8LAzO6pNDnClEOCPjGAbicTxZ2NGkRWJEZ2b/+jsA+Pr5M0NcTJDkg9Q
nIJEFasZuu9p4Zteobxx9A5bNlnAEPqCdCt+Gw/jOwnm8IlPibgVXLPYtd8x6S+65ieJZlfOVmhR
kGZqCNM5Ekab7syouJZoHLu+6OB3XTgEV9Y/3TYhF03lD+f6zg/KsHHt3QTkrC8FCDuANByzJ1aV
eZrdR0wMvoIjbwfAaF7q7y4+j8+4Kx9loXJahPU5gOcFdwNW/UX318tGXGfugP8GH4N4P8o5mwPl
p98kUm8jMSSz/kstRGqENTEq31nmuGIV/+vsbmuijEpqStb5jXC0t0IePtIUQP1SAus1qAUP4lxU
uyRApWxwHD2Dv7SA/Uf9ItVt5AZGgmITYy6xAuHsCk0bAgJK4IcLeL6U9ffavQ54QzyMsUzeny9s
Qg9frhB1168o9xlBObIi0ZG+uDdg6LN8QcCK36xGUgmnR2BgWUw4eFZ8oQRXddujtlDjFJpZWVIW
26iBZ+IvFNu4H7zOJIUXN8T2buglAnFqRgu+BUkrqPyvNBLdRCFRMaipUdfV9l5EvrFTul6sCQg+
HSkx3X1KqSAcELhRCq1HjOBQYapjjC7UpoYIc4q0oKr+o7Zn17pmGYrTQTmi8GOdZsQjd6TuGPE6
6etSGdGPpy8KtA5S3QpyjZR586Vfuu2rBWGnapUAQWQX3fn5IAwnlm2eyQkHLgyaxvgU6NsPsljT
90ezUmPTb4Bx65Um62figMtnVLzq3k0wy/KORbtjtRQNjp8HnzS+VPrTZglNEuD6rrk7j7KwuuKH
sHDlv44Mpi3gu0pavrO9Z4EFHXDp501Dfqy8+yng92n1IxX7GKLoYxaludgXOIiItpyjq8hW7YNB
TZCtOVXl5QilASwLavuwbHrkdGO/HotowliViCbxEUEAwxFlBMil2Un0p0jTzmx6D3J0EsoV2zOQ
VWVbtY3R0h+8c8CL/1l3KQgLXF2QWXrt3EHfkPKpgYFo8pSFCz9Dl2YhrR47LXLs4G+mFRA7HG8X
lDrhJSBMF3Bu4LzGJh4i6BhXL5cvHtTjKd2nXENgMohEVY/MbfUueHBdGE0FDipZqCO1FwyQ+uu+
FH248nRbQptzJXh8SbwTa/m7GrOvcqyIyyZKHFNpNb06dRXjZeoYCxBL3yPqPzURNHAeZlYC0T1K
wGJMxXhxPn3hLkxSF1/St94eatulsGwkddmr5L6GqWFFvehAyLstXaEW4eMYZs1sGReDzvozshLy
ZJVy8XYqE0mxfZgLmMZKGJw5WkjB+04N5f7NEnTqCU7ZnhBjRs9fTUkPXz5w7NXwFaw9BtzLyDRV
d0T45gJHLp3cR/JtQkeOllG62NxYpY9E+b0FxOP586H9DhzvQzTwjSEtWoHSUF4hDeBo/kmJ/06v
q3icPFTy2GanKypUtxc4g2rLP5E12unmNS+NfuojD37F+zTs5Kym2GJ9jUW83j/Z4Bd+QS6Z2dFz
0SyaN6QU6T3tu68ajLwjr0Fm2AMn+bdoDUw5Mnulht4/v/ewQxmlJstPxhAuiLHEMQT3M5j6Rkyr
m3YV5yzu7aSK2YM5quIp2pQ7gR/1M3mzXxvTPOarIgg4i0gF0fV8MtF+Sljq/iMFQDPQ9BKU9JEz
qHiD1KCdIPBI/iKpMWOfpkanJaM+YkiwL9SjT/SxsHecTwmgcqJSSQkGL6K9evGkXoRypUK7CYGU
/WGIRIPoQXXgnwoRqFdMWGVLFVY+Rkc4dJeNtUkEa29qySMcXSBRYTBy+YVuzoG05dHiUlt5qTn9
ih0iHjYveNGm3XBKhncl+XNRIskCZb4XEzAix1Lm3H9MwIeTcKSNIODEqJpY2dA28GiHiLhrCqJU
7z1WTG8/+QFwz+OmBkDJfgExnfQ7rHjPQSMqxB+h4lpqjdLQiTsPQOu+7RN4CP5XnNBoHEpU7rhH
6ja9VKnnE3mkN7jeC0kDQSDVSuJL+oj2PK7bD65QWDcnqyBudTY3jZXyXa9mKtdxa7qYlqVp/U+s
O6KcoYZu+fI2MR/Al1y50XqOsqGKdDDni87Mie7bVaRl4a5ACvDFXueTkNrDvo8wKJhf/iG6CxdK
7iwFDLLIFWT9T1RfM6fWWqOWNYkUwQMDe2un2Sqq0ydiL+Llvw8tkjO5vWXQ5HKrR+5gaOPWcelF
bAHzBk58tde2l75VJufakaqSOn6HQ81uhhRvRHgH4+hxqxB3cGVQIoszI14gqMgGV8AjjXb7faEM
CGmNP86w/BbL1iqd/4Mu4avTVRmo629pSS7mmL9uw12XBPQKZZAMhZyCLsNXjDIl32XpY+m38NSS
vgqwGsShtEOrfVGUaOUe9BGxa87vGHN3k+iYQeozkT1vtFS4ViJ6XO3+kRogkWlZ6O62pMRJj4Tk
5CeviMmGeZ6V1QUL51orTtRyYc2oU7WzoT1ueGY++IT+sNwLVfw3BjKDly900HBL/Jaq8NcMDCX3
p5uh5vKgXDebWTxK2U+Xr7nzgxQtv7xF3P3PAwd1IyQ/EHc07mrVTHBs9h9uJ18RuGnygILIKzvs
fd9QpY4A/NLbDe3wPjltaIIfv2SDemQneeskm5mHkOX2aBnXw5bnO4FmJJxsrz4TexdbPj1iJY/5
HdmLJmSFjgX6VfYw2Kly/5eJgfF2LEuYj/rW1HgJIZBlfJd5hcDWgWVIh4MZ2TVr2a2iGxTF9kb/
+m4gD4FOEAy2J0VZ3GPLXe4w18Mt/TsDU3+UQl1jkeGKs9hzLK1R1x8l3xJU1gt5FIsSZB8RIPrV
wxGNULXw5187AI9e7A9R+IW8/2AGJ8V6XYcrveb+iZwD8luOsRHE1Yi+SwWCVIpxGrJEhY1m/DwQ
p3fzxYqHIjB6PzWsGuvsN+Xq7kzN/lfB1QO1YSG+STek3fy/MG47haKQovz4ot5N7XWkvQX6cbYL
PvcmKaTRNT7GxIcmWv4nklwo9zh15ldEkVOGxlx0QYaiBHNB4uXGt2+Ki/DVWDQABNtZzlC/Cual
Ii2cbSfl0lrxY99u6xHgzYgouZxj5mZanZT4VI7R4QMq+06UWcXB1WRANvmcytMVc8zq5goR1xlv
H/y+TwoA+QdgeT7FvsuGDUMN1UAbHF+2wn0tLcXN6bbwAA31PW+EYCsmXbAK3LcKIQH2nY7ynVM0
Xtu/SgRAg7RrpPobJg9+pORtuxea+ZY0J/fSj3MJjt9QB/iqWMlt68CdMG0v3gLrz0TaV14iqQ7S
KjBg5iB7qX6HHJ9gB032fzOmpuXc7KksXHjU4tGHdcy4Zsq5zmeUcucq4/pMtDyHXnw+3x3LRVPA
mQyLbEzkKyQlwa0KcKMW9rt6T/w1jn+CYloW0TIpykM72haw+sbEzZecjZRBKRaAw9b0XaropTn6
BU6gOIGKGKBo70C9GlvEaQZti8iN6LvhlRkkB4mqk+HlKR6NcxkEDAtnUXMILTDYjSZKLU586M7d
lTTC3eXpBD626mCl6yeehgx1A/2Odqya100nwEshRULKeVeY1D7y0r0xoK9llLn5zxP9cX2yLSmH
RgkJUDL5TB2BOpjMOHjsWve/jhcrOhRmQHX7GyicNbxac2P/Ri73L5v8iGVgmtmB5ix/j/udLbVv
ho/M+yKACWO3dMJEIsw9G4PZrcB9mjTok8E3DsaI6xIrsZkA7cy74KtthWITj4KIH80cFWsZDTNt
KHhmXkA0MOYTIYHEtdYB1avhupgYIx0KlftSvHP5TSurczI5P8lC9hw3ZXrMNnkWQ/pQ+xVhm28S
v8QDqwym1sXuLntPzLanwuE/meWLG6zWM3I907gGqiQCcjJlZMwyQYb1ba0etPz6smwVD7oKa/bE
JmjR0xS4dRcLyc9t5ivV52YLqCMppHRFtLe5CXLmQ1SkjpOB/6NIR3/X4UsRxyQtpC+19zTLC1LR
7dFWi12/mI+1uvYuXJMRO/OFV18M6QMC2usKess0l37GLZ47TAZOQ9v52bIVTstQ6Kk1Y3xaHJAx
pkAdg2W9WZAvpYqnkxIJRZAvBFtG4wylKUbrSD49vTKuLWVJTT4mCXKx/7j8RTDu16Yp/kmJm0Yh
egLrbYZjt25HmRqRizQM7FWmg11WiRBa7ixM272IniziiosOqebKQA1NlExbJz2WZqOcVWUP2ruz
KrWKCqPO7NEDsUNG7JJju1B8EjGJrVTVDtWclUfgiJqjBZ+TnpquDR5goH2jEKLVSGCJ61PzVDNK
IIGFpcBU4F9HBfao140wPnQWJgEsmSFVKWe8yYAEB1CZOt2xZeauLt2Z4s5iTim6/ixb6fyqunA/
M+a7hwGjQxnI9MHjfAxHVbaf33x8nKVDrIQHSzGLM1MlYXWbeSDX+lEIQ0Jb82ABxAKNDnWjW4up
VxnuGAdczE4+v7NmuDoBcYdv/LJpTAO1vpiaKpTNBOd6nHR8z2YWsug01psbS6OLLydtMOQF9f6Z
89MYMJAOQJheOqrrsXu/kUhvvkUzWFrlJNJ5lyZ3QGoOlUolBrrU5n9UiI3KVx2XDwRF8xWEe34q
3Ae5PCnGJDgZw7GfgvCRYwp4ZLt7STC06bOnI6C1yoVpHRvElfTys7y1IQFbAjOvmVvaovatRM8/
JXaca453YbSWqeI5b1lO0hk/w9Ut1PheytR40TjtpHvLojWY8jHW5RAR428FtKDpZyDF5FAzpoCr
iS/cGOoNxibjK845W2xjHjBffABSLZbDFaX94Cs2Ae/WA0hIz+Z3YEwtn6UDbMnklA9LwJXHbQFD
9fYylzpdXWlmOzQ87pyg/nOSqPBb0LzvAviJP9blECZcZLJGRI7P+iE1jeIRHpZisJgY9fL5uj9I
jwTzQNVd3cdpHrJbVev9I30pE8v98k+250lBouA98vPpu9zqiOavpTPfIMTAEIE27L37dq8ekI00
5guQz8YAtKfrh+D9zw8N5WX1ajGLPU2KIEEY0zsGYC3Wwe4uINnA1kHGCf95YjeIV2VtU/Lpifyn
mOJbvrlBRQpmA/ScpB6kgZmp5qf4W7x/6tuiyuEMmBEd90uxgHB7fQABqbdOeKpVtq2bZzrOWUw6
04ZZ5qxOmft8XAq78wuJT4LKDwnv8KaPz1fwX8Nj2ynhjM2HgHWdL+QWnB0BHBZXRFEkLLU81GKE
HZigQVgy5EUwr2nnVp/EGmb/SIIvPo8UO7UTz0725/PBROl1J1pI/pnnn+6WxOwSAtwu7wkc9S7l
X6N914IDZAczf4JhyA/ajGoZqOoHvjXJX1lxSnLJy6VcVABAo0FQyxj5ur+Zaw3zuWLsBG8VRBgH
Cke4OgD2kauIWz9mDiN9bKcTuyU0cvxMJ0nS6PsWnAsrynIvGBCFiHaOUBpSy/E46HCs8/NQvOKv
SQVSoE7Au/TyF2gaFQuKmyMReL2CIoiS/OS94zy51Yk6mTCWtH02QXXPwshtiP2Caxo200USZwKU
NoyqzgROhk+/dd0iHe6JmarEEi/Sfr7GNhfz3ItCraKqPRip8qNCJ3AZ244wv11qAbSBXUgfbVCx
MliqnCGAB8sw+lRfRfmalq/BI/8rGSaVH66E1NctL6Kr3WV508f0yvZtfU+Q3aB0uSMhJg1Qt6XF
yln4bt+fgDoN13nPIxYUGjSLDW5aiaYABNEVTuqJhldfJSp6HX8DKzaAz/9LBdkR0giVxHZwMsJX
P2OHQbCzasdgE2WB1OVIx11qxEfav9dGcmIai2LPIreBUNh5xd4cmgCYc5AbzbzW1+2twrMUwauS
NjmCX0o9Bdf4TsRvKJoJ2hTr10HyJyT/Hx1csvfRImj+hq2xJZiPt67U3FVwBp5hV1jY81VHVca6
W4WNCvgMHCbIMDTTSgQliwx2AU3gYWg3RTZhIex35ZSo2qNpoayhOfFQ8YpyEsi7AP5oHSK52pXe
m+w1XzR6OanvGYpyBfgXBPK07zryJxIegkWLzdCMuYv2Mkilp/l6J1f4eGCTl7E8QRySMkH6xkWL
WcXv67UvAFVyKjctXbBaPvaxANEB6AAM7a+o7STC03JzrDny6EVcr5BeiPKHAAiPXgqCDRjxbJeR
W4E0FP5XTax56740ydNgnAeiePTEogcmd2wJy92TtTBNs2+fCUJh6VLKMrJ3SgUAHwSb4XZ4s6YN
vzW4VIM2Wyn/W+z4kgEoBxmj1J8el7nu0Y7mr1I2194K4IwBQKXHAUC16XFqx7EK2vBylt1X9nAQ
X/qfcS8JAoq/LYGFil4UqELOGbl69vMrcaqQ395x+CRHJCg3DERiV1CkYgylegHdJRA0gK89pq8/
q03YvcFYPThMFL5Wb07t+bw2uOhr9wEkIf64/LUIm+rPAmgr4tr9ZkCSusaitPV3MFZIzpZY7Mds
hhcGcvw4tDoOrMrLUPNYTXvzLbkH5UQ/QqYPZUtm8lyDy5Bq7yv4TR8gEzT4pskFGB6RmH4J/DjH
nMRnxcs5IHOCiBxrtFLFUr+aAxbA2NPCpR3bvGCotzUY4p3AhhgKJ4N3o2XzOxuBi6GM2vrpkcJG
T3Oilt6K0XmoDL6j4ocm0bWgfahXPRVRZ8VXrCejItU+m+HlSSC3jinmgQE69BtwcjbajxVt7Q8g
AnPkTP8RGBJ1LB8nTwzHrgAyMStmpqWE7ZMMruWqvqGZVMI4KPg9oFFceFe+wUjpLyaFigUon4k3
7foZVZ+JCA4VK6iHUUdS19h1B1qOcBixvmK9+UZUDZr2QbKHulllZlL0KFswH2R1M/Jv5jDhWVU9
N2WyBUQkRZm5VQQER2X2P7W9tAPsPEw4ng8TkO51kdjxcIyR+B5kWFeoFGp+voVO/OA1GYuiMaBE
tWS/0Vo4m5Aq3mSGuWioivt8ckZL7gDaQNGGFhKRPE+aHxPAy2738yJp88vEdQVMvoTFxp6OkcjO
6kEiQhcWzHNGYFwdEt6AJqd6ioXTdlKZkIvEe5BUplz86Qrr3gviCIbtUZ5zkfZb4qFVxbyJZ7h/
HIiElO1QuyujRapdKX4u2TRIpMt+9XZH/FuXxU/KQZk3t9oeqrghzWtNgJRIaE6iG9EgkcQqkSXr
RWRFpm8nW3AmJRn0J0dk0pEl78NyRYTPC7jmySew/39oxrI2O7uVFnrv7Pqr2zgekYHOaOdLHXnn
CCqDA1mAlYb16q9Vo5MB+CD6Nc3SJnZybSiM/oV5J8UWLdnra73pb4PJQLy+GYy+Q9G5YD2ZM2e2
LxEzEg13hjOP1uit4Q0gRo+ipq7B8DmgAU834QAY9rm42DGUI+Xbg6gVIgAUFLfcEfAVQwGj+kwJ
qe5NPKcdLd/BXPi2kkt2Obx3n1FVRNBLn2KFHAAdpybs3xQQi7HccKhKGAAlgizOQ0frPldTgKoC
aSq5SmoYJgvkmoU5rdCbajSHQ6IVJD8xPH2xfpIFc5ExV6qz5B/do5Udr6z9y6OVq/nUpOnjOMAN
0cWhPYE7Qe54b5DdewS+CF+9YGkkEmG6L74ey7BJIklGvgjVYL0AwJkZ5nM5gqSO5Y7tOcv/YXl9
G7KlmHwEt5sl/NGl6SurfxxBKS4/5+1/Na/dpRdDmt0ApyjXSUaZTMUOYFulM/V1YwblyaaL9+9b
lA2zVG/SsJUpFmXl0bKVH+L2ZWNbmnWlkYerVj77HemjKaDf3cdbzCyD8s+XePwhLNNI3BdVkFfD
PqR3A4+b7QeZ7G9OQrTBWZKCjTIhCpQ9kVAvVNJlEFPgK0mFDE/8cqZicfDLPmpsF+nK0RC6x0rH
VFMVVBc5MjS35PeSp917SwwuPqOAPLIu0sIMoeBdihZdEm6JLF/LhDBBQI+RSihkiqRqZfj2nEB3
qNqz9bgih7l9CMcUtIUOrGGHmCcD/YSYnj8jMPcnABbtqX5WSwa321yJOXqsfDdYrQipUGDP3UeN
njimNUsShw9GTFnNd0hspvvozFniJZzC7ZdhcvrnTBPWJ+ulyP6Gft+hFxPcfN9j5ctDLZwO0rVg
Q6Lr7S/uURjyIpEwvui8nmEHT1RGm446rBvoMZGEGPbwQLmE4rquMvV7RGm0EBUpN7/IN5qFhW6R
t2TV3THvyd6OfM7eZRZJD0ZFS2myCnEUPOHmKdT1xXWInHg63wdHQo5H/5+18pUhaZ/tz38iNtHc
5nF1HWP1+gIP+7Aq08eyHL80V+6H/7PIu7bqvv/N5VlHmCrATQWFQvpji3IVPky+HNB9vEDnnnyy
IW7t5gaiyeG6y6Bz9vw9UJ30sLWQ4t6QGqAd30Nly2RIw5kov0Zk3h7Dq05HHCObVrAIJhxAJZYz
NjnlOASM/VV56/ZzhhzxYvPI5oORrkrralpcgPyVtv/rSTlIE9HZD90x7bJ8Lfl5swjs6Cng7947
bEtt3OUi4iO4h6XVP8EwwQC1wn7xlV8ki9BH6MYbR4j/Yfz9eqAWz+rKzfeRaDHmAtmiGd/2JYIv
AYGoBXDHQkheVzhqzmrgAkgUNwDwg6tqYvV84cVcZDcBMYlo/X9Udv8DqJjl9gZq8Ecg3di/9X4Z
phGXV1QYPrsGktuafyQXb+SjqxHQRUnmTIe8N1Wj0PRmIo4MoEPic0Ad5C+U1l4qRj2AwRk9wcjR
dewBg9vK21t3gI6h71tZZfjh5kBPGuASPxZc/Yo6H2rQ3ZcDFsLHdlSy+AS3mT7KFUoUFDug+hv8
4CdKB8Tg8cnI8v58WKUzxW/gvxAvFxV0cx03uejp7lRUISvAdh1lilJpL8INCli/d37UYwga2MPo
G/GkeTd6BDOUmdoyN/7yXIVJuFv7zWnzvdbbvwUCK+Bymn56eu7K82U/OueJgrsrgdrTVbVIeNye
p1dylvOuCfQ+wgksGgeNa5LfYuer0lBqRK5QQk6Uc83mELJn3t84okgmM0u+kx3Hrtakiepv7ksT
bQhf2UmAV6nC+XAHyO3coo250VxRkFjm39TQgJxortd0HiHtCe5ceyCxX82QWrDzZvfA74M7sNZC
ZZidVIKLkMjIAskjFDF+hhAg22gVMuJ82YrStztwWS2+6bCjE5IwDEvW3eIrhSyy2T43MFz2ALr4
ZVTx0OLP5EbGKdirc9rY8xq8xgpu68wKE4YA6gXbYf1HOnFBB5pjFf1q+Anor59EP05rQ04MzqQM
mcWqW7Lo2KEQ+emMBP9x4lpll3eSc3iPGJybrc+zRRRLVnKhoQ7eC4XIZuEQJmFwP7E7BBHsp7sa
AZzjUKia+6h8nDrY1bGt5UZmpW+evC9NQZaqEY0umyypHEZAf16XftYqdP8hyESUAxxWay6y19Mr
Gwp4UxZtVbelc13AcoZVlegqD9+uxgPXt8xiPVDFRVhvVn+SpddFq4epNr1/BsWp8dqbzAsHR7FU
GiRoBf4oVvikFzh5lxWPmxjaEtUXiVJq9r7PcR6rUiN+bLpQvjtEXVlkoIEE2qFdUySU5Xuq1gV3
iccbFnNm+C07y0XiwjvwTIp3lvezED8kcJSM0PGI7HIPyZF1U74qM5yfmTB8iqGY2ACChhRYcIHz
dZJAwy9bcYCvzat8nX1UA6Nmpp87D83RAfaBPWWtM2Jkl4AuB7teNvmU4nNm/YrDAlsTW4KlnITF
nNbWpS6Vzna+FUgaOr/9y06xt5WJqBgavHwEexj6qLD0ZPvgvVM9AxYNHG7WRiFh2M6ZDZVeIYN4
53tmqFTlkg/f63MkBY2YGJLKmAcVBfCBN3cxWpMHDgwR0v3Y/nX0zF1zduvvuBRv9HueNcc3yk/u
Fea08qypH04mNJdTirqW5xld9t9UP4ActQCKTBQsxxrhPGEBFFOLFXh++d3UT4gY8Tey+TBBvikQ
ENTgbskke7D+nAfnE8bTpE4++byJUlOuz0YJYW3dYaorbHG4Ir/GX+YuSSAlOEYjYcm11VP9NGqK
G4ZzRh0D98UsE4uDf84oVmrVQ0MhAxtb4cTJHaznGpMd38tnW5UgQkQMel9iFKGV9aJXKTdO+9T6
YpILgu9TgjuUlnanHhu9g4JG8agUtz75b42WZ/HpiNHf6iZq2VxODFYIRsbN7JgLKDJYb2j4W8L9
cUx5I07typ2m1hqSl6rYxo0UR7x1awgtTfAfaP+CBwmTFG0o7we27aBo/G7s/EJezTyW5Va4NI8y
pGjjL43J1P03/7CfARsF9z0bFBXOqumHAaIImLk8zpKCn0alWq+U7xfxblCWsMsUD2jJFBVtZ3Z/
TJezioUCNFOyLpITdxeCrrsRUtkzqRd1H3JzfqMBTcb2vca8HiAAP9ZWUIWhXk6IMMAkDGN2RDTU
kgytxQpiEUbXJTdzIUbHqwtc4LsPWRwkdaCO4F8Bxv2pARVQNt9NTwRrI9JohRrQwYHVSGHZz9cc
gkIlz4wfR1r1E9FQXH4BPoNieNo9wHezwNjsQsDlTdw2KRiJi0PVZ832thZmo4sdJUWcgbVPG/Z2
zDeFEDlblbruocw94XpoCol/q5t3qXhT17cSgcmwyC5LsILqke2gEPAdCPI3XOHoqPdXJPmc4jCl
dVcV1XvXcJIPJC46zMwg0I2NtDOnRbiZCvLjuTfH4M9EUt2PYHJqaTh2nqpI57bxx32HMZWHCheg
0DucYXiAIDui/+bfKhKyPyf24zC/0fIMlrEoGdPBHO3Kr8v6ehOr5IoAvEqrNkt0b4sM6ytuu8s4
OxadM+rfvkmVWxOTdimjPqAAB+gdM0844gpr3Um4VfQa29PMmEtlJngISMkgTqDf4gdDkRgw9Ut8
w8duSh6cZhW0SEYYMAKGnz6MmThUJ4I8dahX4knfXPsMW5jt3bgNRHN8YSKiQgWEV2EoWb0tuSQk
yJT9Jz2vCV90e+IkIPkFCXULQtlW/tCf+worlSGwdjqQa5v5dBLNFPXU7A7AkPVV/FqxaxRCKAzk
CmH8QrJ6GhBRttfUHALHVAB693lrWDnl54JH0WgU8ch1yg3rmQRHoPduMHri/43chbeTDL/4EDwJ
nAWauEmOPSLdP0eqbDwJ0hEokqx4YBWwFO27RN5P9DfUz0mfcKrUCBjy7HttJuZejjdJw3iUdy/R
lSrf+fhXDpcGSa3UPA2Hp5FC0ABc6X1lz63MGeaYW4QP5sBVDgfsefRQFz/i/Gtc2KLljvCeBcTY
933hRxCXH2uPDOW8hMBAMsKBpEoW2P2drqMyNoSGX/nM3rmLtHWxEwQ/6mpOsW7KgNE8PFNY2iic
5txgEM/vmEkHQjhAZYPOyIJ5xF0Wm1ZN8i/ZVAS7yqIIfVtOF6X0sv15LmCjnM25QDN6/Iz/24uZ
nb9965JNldk91yG123z8DB4gxIc1SAfZzrcYRDcJNHGpLqSwy9oLxhfnrrMdrVMGB6sqx6sMbmB0
2GRyxsQx0G6dpgmWEQyu2xjLBzNONyMsBmQvTfKE8kbtetp6wqvAFep0h9YQfcJDrAvsIL0bMmtz
DroMfSdQ6lwWIKBvW7FQHyjaG0Z35iDG6L+QFWte0EkJeSJaCoCW8J0FFMgUJxVH2VPJ5CcBiUvA
HGYjbN1GdyA23tkHazjbsNCVv5rHUisN5ijlYJZFvtOEAsHED2c7ZuQSgcZX/Zh6iAdxPLkel5o7
ZGj95ytX+byiAntwuxxEXy/vzh4OKwwDcF9B0srRLZSLxDDLgksVs7TtZGiIljWDdgTgwbU0tf0a
xer41gh4hdFqP+d1YSs2YbnhG2PIuoRv+HiGwZ4PsIFW/6U9T1wEazOny9jsRyD1O6V1s8Fj2/6n
+wV6Wsfw1O7Mu0VKy9r5HM42vMQ52fUszIXwceZITXxPE5pdKF9ka9DucR2gRBuet4sjytbubZ6t
7JAeuHnN2FmzAdiiRtYhbGe89504uJCxpo1GT4AIolSvW1DutyJ4UpTKfSbXQ53t9ztpyKlRY4UX
TmA7h5fr5hf87y5njONThcz8D0Aa9LEE34cGyPUjfY+EWfLxpHtRudaZLj/zbh4crCGMIoSbNMbz
Pv9bbYAQPAn1i6JZVSzNt5GNb18qmbO6s4Z3kKB/TpQSSMukg2Usi65NwHP1x+y9sb4cGWsImEcj
Xn3mQs/t4I3gDY72nn2EszyPU3ohkZjak51bIdkofwcNoxoFv/N+oO3twRHmYEoTVMXwI77Z3aie
S2wpUD9JcVVLMwZjaLxlPf+JY/gnFO8JqDriUy/Hw9g+aK5khdiC+BtqLGUbSkq1WRL+e5NJhT5N
jELAW77PBUzo0BDyKa0dzphmkrwvu/G9aYfR3sgHXkNEqBntS9zMV59h0/pI6/oEpW4rgFjdrA2m
9oB1q0puQwDIGXrUETBTfmZHJylCNECy6Fb39HUCqBWSjaXebjiUKgOOHNq5tnTzJdDrXpsVr1WC
w/g6r8M3idAsUS/8AsMoRpQrvZPTt1AEN+OCzFJr/+HcfEKb0KhMoxxFTF3byv06VqE3OdL9IL6m
ZilbkXsXMJGdPLLO9//O+wOX+4uLTIJcR7niu0p8IiaOA36N86ozD/2PqkoL1zUunYRqd++/TFq4
2I+ruAAK6Ba2z3zdH2r5tqoeLT6+6XhhpOjpdrR1vJxuS9L2+SXzKjF/ydvfGaboRFG0jlUD7Usc
dOmUetrkC8k2/tKzvuJfrA9YK7K+X/1Qs/XrH0FPrnEW9RG/KQOHwAbNelLZXWWQRc+4wqEe+xxo
c0gmMEcVk8hafL+0Eaxcm+tB/+ueK/RjoY85Ze+A9pnAj7LS3FeRiihvAhGeiQHCx4/Fwjivglxw
V+2L4ntGOdX64LvGQ21FMyypqFimTsqCdGLE72YFxpfhrnWwtAYqoz+IM2I7Ykxkq64v2YMNc7Ha
D0VxhIu1A8kF0FaxV+gbnHjUySJVI2JoO72z/DRNxF4zt257/QTYdmiyU+w+H2XymIrW/eyHKzKD
Fc8hmTUxgOQDxGcfHnpaErhu+X4iY6VENz+NhKOT5rdPmxBpukL6e0pCtbAQmC7UPimYk6KEqF2L
SAn5ARMBSENkeVrWSQk3TV0AwjG6AXMZKtydqKFaAsU6OqnDoNoXOuoyV0VJ0g42+KJiuQzjdFcX
854dRLqp/5tZSosU8OwU4afB3yl4VLpjk2dvIr3d7vKIGtKqz1LKqltsM2Omg13Oq8H9nyZQJ2bj
xikGmwh+UwU86KkFSyjA/F/tZ8tcDw1IlBA8mMi4Io8oJof8LekhrE90YD7Hjuc6aIOfpQzEdPPk
VvZle/DqMlqowHJaCrqf9GRDGampqNjIykv302pQnTQIIW9twzCebOnMEuDQsUdBarCO7Utdw6Up
C/e3zmPK/ML1Y6cLdkErPIEI15v31QG0IgOxuBMhObdCvZ8Vx+PkAYomZOO3hzgBS18Da9VNimHu
XnMbpIc9OkQ0tomJq+EjW+hp1nvFo6oPgvcPWQjpl8lglYHNV8EVZ4yRmFtftQLuE0JLdNCkZSOq
O4exOoAUpgpXPJ1pChw3ZJuHKm8Vfm5KN7j1TVqA2PjnfPR8Ey1ie8rmYRt3eEBnuD4cCLkOGuvP
zt/31iw5glXTUbOkRDH32aPjUJ34Mu58mh1RJ2v4QqDK9hEXbJGZncyCBjoo14A9YhkFWD/gJfMX
KpxG7C0/MIGOR9nskpLU+kBep1X6iaJbP3X44HAO5bjO+SD20lFG8ZhhdtFwTM1OBzu3JRbgdGXq
1eJdzD74VG93cRX7iQ6TEGYoe8v3a1E6P+8nIgROcTbm1qgEAAe7kRc0YOnvHglfqipuLKt8N/2R
JX4Z6r+wdfJN90tDg8E80KDtHsLITmZliU6MqQTwWUVHIrBG3/MCr5kzL+CXgmxQovU9nPAt1/jt
bMcDy02Rx8CTf/h4H1gDFTuL6ccf7Hq3rd1Zqu+tuHSjexfkRR/mnHI24a3QSRJU5MranKkZEOMK
VnoU3YtB8P/n05RxzK6t2n3f/Cavpjw9O0yirG0vwT5USAteZrnedSpm9oULi9yzaOmEzPar9xkO
lVlTHjUGQ4f/eLuWWt1Ga+RWtunB44X2J9qBBxo8yKdilqg5Fozwk5c8Y5BUS1dc2IhLFmMgEH/K
oc4Vm8NLG8bc/z7StTWK0kbQcNOMLuUXlCyGd3PAeRRovbM+1F0MCKMQaJ08rmFCuXI/+zRtxcBj
9jhS/rs/QDSmXPWGqLt42/kiIYS8kObgsirlLlUYEsYHmm0ECFeW5inll3XJWKEIct/gEJbP11e5
PLkfkvU2eQPuhiNgVuc87Hvl5tkcjIL+Mn5UE7vKtrVp/oQxLZ1Kbr6wtVJcD3GnFwuN+b2PiKxg
HB8fQjd7/hg20pXkxOe2yWg2L33c55M9C7x7yv8LjwyLxy6pD7EBrEIvtIASjGwes8nyIcvQof8R
Yca8CvaQ+I8R4w22g5Jw0FSicWAkJLw+Nmqo3yyMRzK3PU6ovnqsDaR54RsSkdzx367jrax17aeg
ZWkdA3sSzbSCmNByrNEY0kOHm7tVRPF+bc499C6G0TMJSDxO+jZFBJ/ru1j8atUGDZ72PN9/SVox
q9fNj+6UN9t1lT1PF9optFSC9ZpOweiQEkkXazXaGzGhL18cwH3lUrTFskdHtdvSLguv5jvbRN3d
gp0jZYBrrtIfgIxgMYZbJSPDrPuvwQPV/ZYUURF9ZjbVGP66SoW7Z+TnNaJcx/gl6nYDzkBlmkpf
FVSYmiszTU1uV646ducVvATNzhFOzs/yv8JWPuK3oAziuKrRrFCDqjhiLI68ESFi7Yx09/C6oAV/
y0iTZPT8KvD36pa59KTwHk8RC1zLNNOPcjDy+vHzQjc105tMS40PPDUg1WsFesLo6o5JQDsEAmFP
cHCUksmjT9GI3yFCuIy67r3ZqqYe4mtTk7itIOykJcYggmMq768QjglLidQfEHCrrXaiyIi5C2Xr
J9vEF+i7llHSdRT/nDXBvh5tH1redwAh4rs3aUonOgDHz9gS1maGdHV3m/CTs9SQwf86IRLJFx8u
whob0rukDFElVFV0W/Hf9GxKHh8a55C10w6eph1CLUhbxyI80bC09hbHFplv6rg5eTxOK0WDGSxW
sx/1I9sD9+q4HeoJ6VhcgeTvpYocs0qDmOXQAXHP2Kems1LFAdjChZLCkmzjxKJoVncvICJTonOI
X667gtrFYNkEGA/FarOtWQYAag+zE7zWyrCwrbfb/cTofa23FRFVNcufvqarPPN4+L4SL1TJmgYS
jKpp8n4FOMM+DB6X0wF0u5MoW/2L9UdswQBZxuvcHVcwhfvJF/MJd2QNzUTK8RXGewKBEH5aUTAX
je0ui0t/cx2Jv+x2xc70mc1+auBbkNpLXJx+oRn+CE+Ex7zUNgP6dWyQB61rTmU6t8pCIg59unJS
VLgUioZSis2iVlWanU5WYRpyC8HV32h/VmN7IJXJYsSxbjPwEBAjbGu4rsUQ5j3ZGEhUTXrCVCky
w3ghNoBWjOeN1mN/B+5I38AHytQ0sBHQ/px87kF2CX2OkSgiXzX+XACVhyoCZSlsrN/32c80YnPd
L2cT0EOaBGoFcsF8orUSuCcYK0OTkLc0UlcKjoNVwOg0kKSfg8M8nSZ49vqrt77PgqWSjnX7uMOV
T+hYWlplg5HLMjC5GdDhIMB4li0y0V3TrMhIsOUqKCJEKj3jnxk7yf9BnhNrWSF8UOnYNP4rVgBe
qavf7gf9SJ3Q/43qHW7D6DkyDKBX/y2826EBMc8LNT0Yh4liKU9Dfv5CmjnByysL/TTJGACiI90n
jJEGFSk4rvg6+OVu0nkNMC0cGlFILq2lw7gF65PLVnpfPV8G1/RXj2mb7+s5kDMLWtqo3zkvMB7+
apMkx2A0/bhf7lts90pI3hH4FUXgMk+vyeWRfu6ZbbPwsUCi41NBqqmKd7PsnKbALeCBtMOcx4LN
RDseJyJBoeyVtwH7kWtCGfXuWp/4fQY1DIutGAZuuCbEKHyLnBrcDLZc7zEVhQVTCeYeG1CBR8yl
huh92DDlS58CYmqdqi0+olRvLE6Oha4E8yHosEzbRtBaer8qIUhm+3NzX8fhc9LGxasrVDQzbHIx
p4iUNjyJNl3Pyvxx4nkV8Ysl+g7uY4SnNVbbXmidFz/dS/QCLVVU8QawMu2Gcb/tkSGuIGVt103p
0BVLvG4hrCpn+2x5g4VnHK3c4UA3kWNLv7GheA8gA6JNuL4Fp1j6TEMQ3TE9R38mIFb+O9JJ7oOX
K61+d2hHJAy0GYPKRXFea/nx9VCp6OEL6WzP5a1lGVoPyCfPR5fMudYi4Nnpf88z9ySJE890OIUp
jEnDXhFtoDfN0spCGbYJTCBs+x+WCaGmTY8KaC/ZXau1JV1V672cKwVlGrXzOH2qeejhaSL3E2Kv
T3In/jyHUPpVFQesjeUbp9ljVdRB8jpnCsFJ/ofzGzPkieIn2mrd1nYOdLilWWgKI4fFQ+3CMRok
bOGucBOBz5RhBHE1HijJJbm71rZakECr5x87Yv2YS4bPlT5b6KMGYG80n44+QBn9C9L/1yLtb6HI
p4L7NKPBO2i+x7pjCAnlIVqcMDH9YLP7x5Kx0knD3IhcMJcVrbP1dqaH8JcBmd0+UDKnLGRNZhpH
BchTzcdqOkQq7O/b7hLic/SMY6zxiMT7/7Fo7LnkTCZWmzDASG/ianwt98XQEkLsPm1IJBgogysd
O+p5Dfl59hbQ5MgDaKSf+VWI/Wrkigc19YV6G5yqA1tv8WWhcThqfV1sXg16P7et7b/G69iodwk0
VWo5h89BuQBeE02aFLhUZP4OzD7aPOrSgw9G+XMFePM+ILqGDlGH42uhMkWfJky3uDJpcSkEg29Z
RSsrxMOWvvaiUQik69YP+JfGur4l7kpoothiRCw80vdo22jMfSENo+SeF7TBl5Gb/9DlaB0byEdg
U6KCF5QvJleWL3htJ2ZWNDY779IyWGoDFnxLoVT/h7eRRzavGHefGViEsueq6HjYn/hLbYNDK+X+
kmiUI3UV7UJDIbAx/LEKj+dB8RrY9Jcu1UfKUWr17fcH9Dm9Z5q74d5xL7+9hjTTjxTIDkmTC6PY
epWTdiWT09e5E7NMzswlp28s3XhQ2GNaXfreA/Pk3SpRO595lFz514K4L7Um/Oo4ygr1M23tLbo4
xSuFDX133ZaW4ygXmP2T+1pDTZBIMO0p+vXlQYfkf0ILfl0iN6kzU61Mj7BQiD/cV4c6kArlZlw2
wfzwkFoSlTQJIzqcehHNZr3RcaZARRIA/z4pZw1UHVa80Px1iBcFLbAnlzedsYOyB/oOzMeE86uZ
+QrFssU/tKA1n5ANsAE4dMm+oA32DWY+t9q0//DcP6qH4xq3WaY8fvPkCiwntnz9EiPec/rYywyJ
UVGKtWOjfQxIJxV1dcW8qPEs8oXeT/UtrtpNATUaBeJKDzFrmVW3vYsmCldY8NhMJuzpXNAE+YPT
jRoZVp9wWsKxpayOM1H9XgQ6JkEeEN+KCooP6Kynbjanc4WHtpfxNUwwDXfI+CwQmKilvPPzTFO1
HuXbUe6rZEqFHFyqA/+vXoSAbaXS75O5gb5XOvB924Lb4OezjNGHOnxs4gHl04ouVUHye/f05TS9
WppzUPkqfkMflbNhpt00j7qN9GB/GCau0t68iRavGYbFBXrow7WuFxq0SLFGbJ4nP4nVfZoVB3Wj
6ftbrMHJzd81iWCC67szmBGduNroqYqPKk1SGHUCJXcMivfAsauxA6wMPp6Ak2f8n0WY+D/k9abh
+SZ7pkpii0q6LWf3KF712UxEUW5BU2jGLbmsn6yOt2nt2vWtjjdvlLVjyxZLMkDSbJ2ql9GR4m0m
mk+wnRKmgz5t+oKh0/jvoXYWxSsW/Q2OIeMTJoaW3JCm+T25PcRap8+ewpT0w7X+2JIQWvnjWn2F
Q93Hk2rTd3/aVXaDk+aHO3uVJlkxi/TB17AMxlG82kq6SKp0/1EDkiCn28Z/dMpq5Ijjst2E+s6S
U2yqwQ8OaXZ0IfT2Kp7Kx/rdKr54nItRtIeDKq6MmxGpjfZm09acMbjn0IEtHZvV/ly/lbtGx/a1
b8Tvi9pgilHFywzK5exJnRsQuerbSm14Z7JKkxnebaHQ0OFtkS41A1zknNoCuvMds9sZYwkO2Jxt
6Atc0rd24CRDp3+3CA2T2n6KA5hDWCm0hrO4qqDRKDWThkrAFYQm/ClAkPMniBOMSGlU77OTEai5
Ia317ZVc/i/oZd/WPzViiHV2q7554Q1rUeW4ekwglWi2D94aTnQgeF7GJlY4PN1zG7YuTsBOiEdp
IUbS+rcL0xcicREAnG86fkRwDW54mv2gN7NOdCOijfP1GNMg6cM9AWRIz+a0sIK+fIzbXWOY12zm
BsCY7XVrNjaNLDHfAaPYeybsKnadtyoU3HEP8NY1u2/oefrvUPR2fcOva+AV9Pg3phntV0A+bw0O
WZ6Y3nXEHDEAXntF/UmA2ao6jTA5bprhRCGp04f9owaxuxOhcbaKUQkPKW9qqXQppBf/NlllNpn1
tdaSeZnHkwPDQVuO5evps9qNVlEqHjn4nqpxs8sXLwGmpxOpcEOdlbTPUagCxYn+30bONZzB4cTe
IgiP88a8OnouNeJkkjVd2OTW7wqblPy1ll5h4zfr28s0NH1UXiJBB8E0l7KuvoJsR6DD0kUsKYpT
h2RHZzdWXwWCPpU87bp2bNfLu3TIzSA/gOR/p//DbOYBO+zuF7IKZRiSiQ4lViha8nK3w0/52rli
z9RkK7jL8tbtG65VNZyXCTq8OTeBHqauRlO+xk93yGmXjWUMIIGfXJfqq3/23ea6Ar/SFiuWS34t
boOwBfMZhy7aKnQaFVva/skEv/e/Ev6OBYHrL7yDauz/oP3gI2jYfssi3d3j3V7EICDo7wmg4egS
aplGR2mceHqFqcvqWKQ1RFhggEjn7VBLC2Cp5HLstCv3t2O6W1gRTmUEoCw/j+vDmHM2q4UN9Isl
i49zL3kEjkWcS+NrhwtyJJ7e8YLcOSrnSGalDctR3vkVAIgkGaiyl99rsnkz7lAnzGOU4Wjla9Nw
zDWwmJrWyoCd/mXJSymUODBQ8w5Cnu2oxBJBky+fpMR5dL+pOG3+PuLDxQDvAQQfty1PnC2fW077
zyxNtqxt7qsg/3A0VUQmFgiYK5Ewo4qLad2lGPqUOkRm8uEBCHghmwd1pE/VExmWU5zJIesp+48b
bmESQc+outLcsaT+ZF62VFWm67SpFMiWmOm97yCmqnIz1/gx+dAIr29e2ojL6G95GVzcSLHwpzeG
3yeXNORqVN5Tv2ed5dI/bFcedVhmSW+L6ojkQmns7MTapdEVLw/YMpcwRm0KAULpaRKIWui4iLDn
yP7r65nlUJH4Xk3E6qjR1bBP8jAFI+ElUWfJ0mgtpAXDBdQ7fp4oApc0OhKT5krkUQvJg2SobexT
A1PZyBTZPEv/No7phdoYElZCDhUWmHp7EToZP9AtRi85HrU0G9ovhLqwH8wg8NnndHDzgFqzkXE1
1O4NpASC8B+quZujaVIgu0mk6Z/h4k5wc7vnAVxnhr+vuVicqCMX9HgyCJhDUZjBr3UfaHN7KAPQ
zrgNGHvnHWKqALI21jM3dOJCWoOxonHRKKeFSkC0FMIboVjQOI//UXPjg90RljuV13PWJgC1+kOQ
Mn3wCJhpPgdml0QLvTOGjdfgyiJCJlWHdnhCR+5vSxg8NX2VKnfBvtGdTbXdrHObjqtK+uSCm7pi
oHjIxLOyvt9b0nOXGA5XBNhkGF3WZQw/fO3ig1HdoRHOPYeslWVSoRMF4t3MNNuqBKDirdrUg8kU
j2igD1HHvXSFezBO6v4LqkFC3kznS0EnMU3r/thNDGVnDud3LY5Sjbl6IPWfFHvkSaTVT3KkvOT8
0A4u+tPSrPlKeySFn0Q6Rl0LE9aCWf0YUUCpMjZP9GtA3aCcshGL7gcTqgcyR5JIU/J+cnd/TiKf
D6pRSVrUfme0eQBQmp/33oHS5SHqZGCiVvp0sqULEJVdjQJT59nuEV7E2zi3C5C3Flmo+LOgl9gh
UKolrCro3lEtCmKUbJh22L7JN6ybL9vIg8yz9kHs4e7pxRrVa3NPUxoHNfGWo7lGrGVBMcDzOLvU
vBvli9ShatwW1aiLI7HyHcY1gGxSMwlZyv3MEm0oCwpNZAHqG3jcJa9ilFou7kUD5HKX51zonddk
gBEEMH1DLeqByhrjCcnsYaG2x5CNqvUo9Paz6YmE3qnt+gzt4cW4oMRfmD66T/kVRIU+pqKgrs3L
CbGdrDbsgzHIFdgOrnUG21nmnPQNhoCdqAzPnIj2rcwnj7q1ryPslksQ9mU91PVwmbmT440tRaxw
l4sZKbt6WRaLVjeHqk0HIKc0Smqnv1foMbLa9jxL2S8+BFA0tBWijYKANX/qOeq4Se2JnOPOofFQ
pU2FB5lH508ksmcUCGRSC25YDzRNJJ0pBIQhwS9E7uyNzkuNWY1Xl2GVZ4rPlf3yF4dW6n4b+Vum
cTFfxG8EqdSot1KljlVEIza8Vu1HTktBWLD8lMgMpxVvelSo0tGBrG+DTqtCRVmIUKot+2sWOACx
t1byxtLEt8NsFExMu0x58rq1GN4hj7ebX2iGH7pNWUnc9tFE1WrnvlWaqVk8qZOksWyYcHXHEiog
83DOZv+xk5eVhFiQsJ7ODtmJ3L5W3syOILFFwCFSaw6bWIhBHoG09hDcZdW1ikICpe0ehOGy0fyp
RmDa8V3SUIXLE8l5rnO1dP1no+Fl4xCUpOaJvFGkcQlmnoRO5ipSEpD31CmGFs+lFniSXvky7yN1
/EerhzPnYpLvR8HJg1T4139GAG27zcSXXjTz4kZSewHrC2aNRd8Tmt8RnORli239zCAI8d04PZYU
6GDX0ldi3dwEv8SlEdxb7rNMOaxF0dGN4V7Z0ski5ACoeP7iBWOpJfwlZAMS7PHyBFPsF4bG1blU
ihnN6e5s8eBRSRq1WXL8Ppv4bsx+AypetBPofP//86pZoDf8szCDW7tzS9/mOkJBRvL80XsrQHT4
I5aZrZrYVigdVp/GfB9A2D4FINjlJ/KMJWRJyvJDdQB1HYu/b/9th7+L9m+vLTscm4UjS+azpkLy
HyWE4Iydn/1TGxPoIhNbsZJBdxeomvO/bpBUPHp8MBSesOi9+b4nkiX044tHgMOMnjTavoek8K/+
bjpNrrKDl6qvC3r6gGkE2/Q/rpAnY3yx2/6mtDqjDJQTmFPJDiY0GT1JqVep1NWuNJ3e7Yo7v40W
zpXi9uIvosyIdt9i4LLDVb3+1svwLmm/gHeM7F6aRNrV4PcahQ8TQurIyW+HTMxESM/BMARxP7Mb
iN0gWQNB4zf2LI8oKE38gdM5w11q5egqxZPgx3EFz+Ic7N9rgRO5NLEXMXZnE4uE82qdTEIWaGHg
xpBajh9f9p0BmImua9Q1s4ACZhxamknxBOwkq6DkIHhJgU21yCBiVTBGHaowc5awTzWKENqEtPl7
OwdslPeGjnP+qEULln7VvvVOZmLVXp8lLGlRQIqzNurlg6LTdRmKOiZztLXOefy+KX1ytddNTTif
L1DlUTdbd639bYpc24SaI2KbAcitcPUXFaE9Le+Tk8xpWbiaowBmJ3UROCA57dwniQLTV0voKuBd
lxL4SsUDSEpDQncCPuPJ3gJMMw2v6T5Os4dCwOnVAVhPzVIWAUhMcyffeAGBloG16WjZRu0WdaEQ
9cBTPhGVMug1r9Jg2T+LTsAu9SnekWgCH1EJz4LjB1TG7lkEFspsf+w37ZSZLwE27bcrDzOCgN0k
giL3ulFRCqRot63ZWem6/DsZZUlgonijH6iIex/WEPPcryVQdJjK7V5QzW6p+X+Q9mopcUTeFwE5
Dgo7qdbNkmo8j2/E34lzZl0D+z3abR18hYeYjv58iCNVV1qzu3beWDiYckx7Tox+6ywY/4jI43AA
/OiOPDdnuq4B3LLM7Y/DwYaTswVRLz7OQyaFRliTjvB5FdhwsUVc63EylM0/4lofhFywFquaZK5J
BQuh5lYX+HtJel/zRMKA5m3fAexasnP3r44ff9ZIbdsjwPw/KVn/vDp8BVjxcJec7RIoV7IxLhc1
DWLW35o6jX3oGyRoJPc0jo7KkyHLq3C7IR5G1sQTLGjTJ7j6xIvVU48fZXYQOb7fY/UDgpmHXBNK
/xak5XLzOXRM+4w/uxfxTqpc9nD+41eROzA7WticdwAx2G9OanSUPHo7+jd+ZE7eW0v13Cy4Q39n
yoHfZyPd5hhdwL2cnJ+VVrScpZTft+PlsW+SJBmfHqjEO5oVvp5pysaFPqVgK5vfSWUgJr+oPFcn
Gy1qSZ83a4l7bR1LUXBPPHBuF8k19BHbDFPoBPVtRaKcEFxtv66E8fITNlfkVZlO4Oi9VcKfEr33
pGUtIt/nRfQfSu5bLCGktk1hzqRA1MfmTyCpO52swJJP16ME3XbjZcwkOsCG9syANbkzHy3rgVfH
4JBD+MAMNhPIYyR3KEHyRzEpsIrF+qO0/7NBl7vJY3mOp8sTC6WA+3DvTPcZxKmCfantqHQyBjE7
T87dPTI6K2SyDF88Eao94Qg4oeQpffHTAkY4YEn4/Z/xdskf8neq4NTCaoV+bk4lyRwZlUFFY9ls
nxtSf6sDDMKejHK4yl7IGY/RhaEUUy7vwR4+u/CwxbKIPNz+The1/yxhi+QT80ppB6KPSrzVB4qX
Ntmtcno1luqSbfMV1jwxwto8owkFqCJDUjUhlm/X4Z08ilCG7ZULNxJmhSxGWCO/M0N+RE7+ORFU
f4B26sE5A19Tubt5ANGHy4Ul6MBSSuSg7tdvigt0lEPtPpV36sU4brSEY2VjK1U3CjaMeA/QIGUN
agCXkCjjExvp9WKlcfZwc97+OsmgzWTXjbDfrNQJjUwknGagR2S6zN/vvZj+T4OVgZjqBrtmpDP3
CnzVKrSA+3d5PtdUp9b6IvBN85OdhPv8reSW+VrxzsgQI773CVc1EAD2SX+KXfqI0t2V6QKe2pbH
exTQzzdPUq1UfMtnzWgYYzPNu6admiRPuAxNP0yafCbsrvCinF4v1osTFUXz25yOPbLTGC8tYS47
nr9WLB2JjJ1YZc4zThoOvHRrOXyLRqZhBGtTuqYWKrhO8nznsNnzj8ud/lJsfRX8zA0cx/4d2k3z
AUA54WhuPLXSgjvrPKUcJnzj69c4Hu/Z0TUvLsG1Uh+eGSYOX9b8gWHj5G4ThXGr4Wg258wsMWSC
ropxsg5KDLS4S5hL2JxDGLgXbnIO+CXzaG2OlAc0YgjMaeCvecfFwiUFk4zvUi7egx58kNJwy1Y5
fngJ4gm1Yf4oujuStSdJn4j/65ToThCFQ08sSnsrz1nmZVIsNQoHAgu2ubVhsUR8GQiCoHuj8Rmh
TrU3FwQ9/U32nBYRN+KChxzEF3yqAAU675P1EKwNT8G0L3nHxTnqMdJA0fyoHcErUj5KVkZsneBI
yioY1c+6z8ClCBbzm6Jc1HcOTvaaX1BcURaWDL6wQg5av127KkfySGPZCwEqOKqKjNfE0B3KBG8/
O0H9iMma6YczkaAf2KRBBpMjYsvolMbBkMGmtnfGdQD/OTkDBFaop3/eg3sTBc7InMlAsg/2tgBd
AZs2Y49vRpfnOGt8yCs0oAS6E2Ckb12ECt66cU0H8j1Q1ndSo/h6kAjCT0YZO5GgujE4rgHMEpSE
Iwjq/LVRQsYDq5fplislcNAVxUcP4zxH2CkGveCKDWaLg/u7kxzmCbACninETopUPKKMMTSRFlT8
XZUNiVrisfaeXjolfvi4yMgRkw76OHwInNNoAeWU/wPOPs81I2mZbQmZT3fcxQe8IdjgoJ/TmoAA
pH3t0NHURPnrmlR21Y8F4F7RyX6pvCUACEHeoyKRBZ46CvDmJWaMdXXtg1WagPztKnaZECVMe+1Z
x1dxa6olo1axMrrRtnpclGNFZoEszRsWQ1VjeDSbe9LspwydaLqQbYUQIGysUdE2KTD0bkRa44P9
GGLkVZRnQLS53+QpEzXj4whwhQtWQzDN/leuEMGDFkDwy2OGmgthSMy3nCUFv08ICzuPsSe3zc2c
oojKpsR53cOz5n5QgvBsdJT8hjyX52IFyvA9e3jVZN4ckI3qS+fUoK1QdS3iRSu2xzDJhK9cKHAb
inFkfBNwHezya7JXxbh6d0yGB98lH39rknHyZYN0FuE419rnT5o98/UCVyw6DZINveiWRyr3KRb9
6fqFZqLAB14yxPxI30seyyO/yiaJEM6gxoe6X9p6wx9YtAOnLDyb+/nfTLwFQkOIFtUg9RxxwhuF
dNhsmMCQTHwB8gx+3hMVk7k2rS9zDF9Zr1S/hm0y8lDJmAVRkNK+Kc8tdIQcTWLF52IBpNtcclr5
CxW/NPvUfnWI8InnX4jZeWpE8LHHeTSklK9IcnCqiYNuBiVAxtxz2gvYR+LF+jSJAlyWRIpu6dZh
xrJZcl+gDkyEaJqc1SzsmDdldXeTHryTUj5WdRCtDeqai6JQgLEMDK95OHsnwNSGDXCzctLlOp1J
g8r7omAg48vtsncoDgoqOizuk8shiF1l8g8rgzU0OjagdkDn99QE5C/TE+aCIcbZTOfzWe93m30v
PWhcv4oUOEnkf3tvB4lX8hgjpOMLBWXFzr+EiH1vIaLU8v9FAHfeOKFAaRTFU/vXvsg8pCMUI/9x
bX0U47IUoL2v/eNhcKlWyM36L9JrIiEpcjJA0W47ZET43D2kO1zk4PEJMGyEAlOwOMsioDpw6gp/
zPLTJFH9gEUx+nM73ZFwSjGEdk+yAn2cWr5QLaSvYAYAdqhQvFfMyOH/Q+9+7KEbZSd2bVsL8NFh
ajkiwUJcLoNUwGI7WDjCWTH0BaKSNMfXntMkF8Sc225obl3hbDgl4uKdV9/JuMEj3qw19ii17RdS
4wBhxiLLsESgL/xAnWPRNuCZ0xRODVpdmMEm9ePJxp/JGX+Ok6ILqb5JPVuZgIzSzrT7e3wJL5qy
22hVWDDo9Ip1aV7hJk4r+fkZZPSEL7RSkJXuNA/oT5qHPywqHjeAwoEdRFC2x84YfA63omVvwDmm
spXt8yLJOwAx+q9NnAa5uhbkUurajOFvhBYOj3KFN6Rj7L3a7kQwONBSLoh21nCEUqcECyqIOZ5V
tsEkDo+xNHrZeA3u7ifRvmObzD1M1bAAM3LwfDWf/PCKNw24vN7j91Xqo6ToEx6g2+rOtfPCSGdC
SY3wHYwP6eySOvaTV+iFi2ErSo2JHuP+Oa9ancSj8i5k/lxJjzZSrcI+R59u+ZNawIbxy8miJbES
RrAFZC6yBfl/CDNlBnYZilLiYc4UtX5bxFqS3z+VvLaT81YD8WIOY+DRYSP9WzGkKAIVplTn8PI3
1eJgC3rpWWrPSRu2LQgZ6DUqdvNiW6yk/hjfwGOhNCKLCtw17jde3Ryv4eaadI5zA8JpTxB+02dU
yXENokiUzfCVFgV8TflyzqXgUfS8Iu0wb7L213CA2euqGF6UqkoWbjkxw6c1gxsMTYUKZ/qv2C1c
biEQrQqDldS2C+GL43AEC5x/0ZUKnJKsnjvel9R1D44VDq+2rqW7Uc9KPYXZPZc1e4iD+kF1JgSH
XYNK6pSljT6fE+GyFd8nQ7ZKh3lCOTEZa4eT2RY/PtQx3Dh7D3CNBAsrmFsDRRbhZc+Q0wqeRai/
DsxJrRVQAr+vCIVRkJHQp2ew6UWqnOXANONZ0r2VddrG3jwAuqV1wsLOvXbOs6W1z0dhRhDPUNR7
/OUNXooopx3KyefGVDLSQFPRHlmZLEXjEhBHs2ZQ+puKrQ3Wd/csD3xHUpTS50sySrvfEO3GkO7G
JOz73zsbPGNkclszsV3q5hHqgkI1OoSjX/gZ6ye3+4bo8jK7FGJcAMU/h7u3biRldgM3gCl9341s
kIoF90xUfJGl07bJGf0AJN8pUdEYW5HVaLO+V9lvYxn/GuQsiqVrXxq/rj0RC6wsRh7NJZ+qpho4
0BY7gT8Apfu23ep3maMfHyOjMiq0ey7FYtOhAcSMhDYNlKnK9I8OkZT4y+rERIk1mbWlt/TXLhRE
DVV4tBc+8nrSUUZeU4m9M5RNh2EGFJSNKo1+VNKZRyZGLiphPvI7/RxqAQqcxEvtIuyJUJCf8vib
KJNR4vNBVaQykEaMYX9LwB9hKHCYGspioNBFMV+VVaFU5IIpjcGj3rWCCjRdqRqApTxtOVdYDklH
GP+SNNNadA+h3T9ln3Ioj22pFbPz6HsuD77P/G9nFq+InrbmD9Qeguym5hAEUEsIoXbC1i72MUkr
XsCitaaAdh7PhUw2/0W6tr54bTwp10iuxH/6Dy20fTpYklpspESUUoKtFA5L4ekBjcq0G6bg0wFT
9Z0ASs8XMIAgFqOVxIIjD3v1Ym7O4dIR5AyzRW7v7cSx/froHonAVUl5KxjW0/M3b3Sjn3hQQjyd
4d96ftnhElYwUTmTjglK6O6zzViUtyBAZNpA9nL8qjw+svddKJ1AKBbMDPZtlVZNnKs1WuLip6gj
gM9gJlMpNgA97IOIHAP7GBtJ1tYDik8RcrKqo/fxDY4DacOUMTsl41BH7tAHeMZwHxNSGSjYxNK2
QjVeXKPdxzNjwSQE1FjEU7oNqoqlJyVCZpn0w0QVeKRkvaAiGttkib1jZNJa+dnuNomnRDg9YBin
jTR9euPuyekHddYiLqNM+xay6KuBC1TVsDQm+V20Bagm5saYOIVHizv931fz3QAnZSEt0mVWtPza
Ez+PbJWg/qi1EU9p607XV+ojt+AsBt0OEJTsUotuf50nCa2W1R7zdJF+qv9M+2s6slG0lUirUaRV
M1J/swBsvivZWTAh0GmnOB8Y7AjYkWFhfZ743I6fDvLc1zk0f1HTb8j2on6pbpSvkZz7PNNKjyAr
APhTOSN0gvBfjPOqe72wmiSiblTDRQZh6YEL+FsOhlGXTrMouLdxmfbpP0Gc+3BIf8EgKCC3aJ1j
lk3zOKjPGyfcQ+BiCRHzcTIgHi+MNvDyu5f9MsDGUjYzKUD3M91R4XWrnh7IiVlkmGtecd4TsKLe
OZXuxO3kEOSmePGx744PGggh51S6NT+O58GQkHqQ98A8UCJMt85BlQEVdBIb05MlaiLMfUAdtwHh
M5a7R4WheS4pBO3+1e/MxwebUc3p+j5m2c0JasywvOEGtEpAHiOVSEx6yBIhwN7HFxzcvSc01JN+
lXFbOmyQ6PgQbbD2O/KhKuSLlStsAoEl6MaNuM56PBNmcLprP273/GOuLl84Y4hKwfc2QNgKRD75
6UvYbVbagOgZ5PfjC4b5+GID4Ee7EHwvg1ZUxV5DMemfRLjhuIEtl3XfYp7ZuI3GluzXFfke6fqv
//ifZmDxdV/q9IPmIiio75lmRvGHV8ZzL+F1n7ee4qIXtAGrLJWDVhjNkf/1R5fRSWF3FUDqT6zW
oBRWi6INtK9q51QD1jE+5uRIG9WlVHrfaLdU1clC8kBWwMk+9M1/UnlPgMwRq0H2VX2qifcGdQfq
999PCYI4LohF/A/rWyakUlnH6oASXQK2AelJzwSd6OuZwAptSHMY+0SytAxencUzMutOe05UZgRC
ekNZf6S5afRvb8NeDxmycAhQGxvVk6R7PAFqTA1y0EApn7Kry8yqYPPQw97dmBAknaHoEfOu6ahN
ZDeMaCsbQxlVoGa1g5jOULAT1WzXcgwAk8zH6tcwbJh3xxZnrRpQyWQCZO0det0M3WW5NAw8bqpX
DIMsgXyPT0fHRe+fnppuojZnb1ScrC6/oLq8Zk0Bo3IsbqTb39CkEEEnqKG3Fc0OSpA7FhoF9FG+
O3rMOSRlCBxlJupCookguFGZvSRKFxvMBwVux07m7qNux2LeC42rB/LKyxpVC8VhPZYBl5Kq1anL
rPoHBnmrFrFiptUEmR2QjjQDmakz18wZPvQFw2JZuH5hHa15D3SyFAM5yQMAB1JUY8HXuuUvjXp9
JQJIDTDjdYcCMEyuV4gycT9LyBcVeD9JG01pbYM1IxQbdY6s7inyrcd1a326MDecEaa2r5MaoL3G
EYMNkSlv8MS+MUWSVlgSm8YMfEBpJ/Cp5GIqprUSSRZqCIqOALzHswasDDau6m3PCWdhEQzAmhDb
h52K5ShddkDVRbe+n1bAZfUKDhtenLdfkuaobzkKY0TvZSf5B7x4VkvcbLxPhsegq+5sa1dRLUJk
OXpPgH63nKch4aXqNlyhpWduZGQqPPtgpMIaWdwmNcsUMKRwklaMqP4QDK0ZzEvfdDsEuk2NaqMx
MhMrWf3500O0vaq5uxW4jXc+6UgIHlXXtRnlIv61nNjpdzT9vyuLAGmKb/pF993iEKq+mqkHYseA
nKKWQt9TRbgrW5EzEVEEUV9lhHFCROyaxsL6KQZ2z7LI1BqdorI24Z2E60+gBOsKni7oJlZZ3o0y
TChoVDm6wpGnryeZSz/V9hLSDDmMKIkkFbPThAiXc1ZKdD52YIj12RbcC7yIwzIpOARB8LhirF8U
KKuj6nN6OnkobdEsHK/4XKM0AQ7JC7X+ddxhm7Nv7XETjBVpRkkBtB2knm3BTiHF7EZLNb5zDkbi
L/85vywm989GnUTPcOlkmvV2W4wuAomK3trasU3I2qh25CgUsDsolIb3yJHRjrUwVSx3GHHjBVv7
5Me2uf8k9ezo8sSEsYtaHWGS9k67MK7m7muDvB8SlS90FlDudb2Ug9VcVVhqxQUe//i4Q3/pBwxt
68XekSV3NkW2QjB3rENn6NxXz9TIRzYP0OX9MIR3d0hF6fJiU7/PTRgyXZGZVJfpJvkSV9veVOuX
8FDx4IrIXaBUflZkiU5HiGZBFYUyzYUFfh9HavnwXP0Rbqf5s26UOYv5AiBwkUq4YNNeqdPtDUR7
0CjPejDE3cByWfkSV/K+p6ZTSyZYAOM7spN+lt2+EsK4S5GX9q73VmgbKegQ5kl1infA+EMH68JZ
8CXApxbIOI6cNsx/i7bf/GaF3lpAVXF1aq3Gn/ldaKJM4qG+dSFSsEoSvu4pt3DBoWML/03BVzGb
C+OMrudF+48PZ3fYsu7IHyMDerm6oFyQ84KA5/LMAqmjGDJbboUBJJy7klRJM51kRgX1szV/BCjm
N8xDEBsqujabNnqcgMnru6ZO0lVZ0k1+fKnudTJx/I8c/nylKgeke+bdOQVXZ3xWvd30u8SBm7hN
4nTPC3V0cmLM74ZOhMR8nxgRgm2T2q1WMU8MykFNlQHV3GCbQnvhjHSflE5AT3VWGm/M9Pc9geOg
pOaAWj7lXo5h2lDmvjVJSBfUyBzaLeqe0a7w8fl6RNt1AbJbIQ0KwlWS8WpgzYpSFwFhT3Mbp8Dm
x4iAeVGNGsTgFmW+dw+QzZu3Fimz/NpUxKbCi5DG/uA10bIvs8UbxByPZ1mPkXUchxGgCSXmgQP0
773zqNkJEnbMnHjuad96Z5A2rj0CoavA/VyGroHubvCZkpIdEol17SmaZttsVuZhIgSEr8/enmzp
ErjMQWn/aEoDEfd0iRuJkDiaq5jAWZDbIyCUdMnITH/Ap8ZUfbYFKJkNS3MFZmUpII3Ho0wwNTLD
YPgDCleIOcWUaexqfJiCyMUPuwx5+ojsHmwRjEU998H/KQbVz73w83s94VmGSRK8Nwm7qSf6V6jr
Mcm8oR/hWczOyc9Ye12C3G/XBijCZVfD3y9KMsX/sc8gNE8Lx/9LTHCGO8SHmv5iDvwRxpuO4MVd
kHQct8pjqlPF6E5fll/baAUAgG+CTsVPiiwBSGR+pWlPnxOKfWjGTsefsx7Xi9V+31xjRl/wCMn+
rzVTFJ7lpPYgKllun4JlC9HSgsgIxL9AmO6LlnhATsmaAHgVpFepqD5Wor9shvKW7AyCpuguhpOp
BCczYDPZfSVhJmVqxoe4/tbiZ6NsHW1aH+UVv+DG1vut34qcjS8rTXt3CAA5GHf145ekDtVno+96
cLwkXgUhmLYUJX/5AqVGriTVL8Gz2IfnKsY+/pAfFgBblU7f0YNwD0ofSUjp5kNLiX6Kgurgcg7J
+mbY0QmX+ubaqDNQ8MRpxzwv4JXJ3WEto0ejDNDrxwBO5zA0t7Q3akzjltHbLh//BQkczXtOU/3e
h/JpHaAjrismYraGz7AYA6Ke01VnXlgBdshvaHnJo2SBU0OVw6bslspyqk1ZlXHAR73yb5dxceoU
+g7sYDzVeWizqbIMW1MfNxqJE14dv23Udh7IGn0AuMGN9Rp/qyExVPIEe+0sBLCrx65Mfq6027iD
uI28ZmUyH4MKDJPqxRch9uwTYRCYl34aIERTwgIZGhsMM5BRep48jjeIyCxUwu44wcHqZ4gzMJUU
/AB2rvBa8tSXf5qnS/w2Z4SQF3DRa+QZQfuuqu5d5sJY/zOU+euuFtO4hvlGczcU/RGuNamBHejM
BuMjbZcnYCjWXvpamxdBUZ1kV65ZrasNduOg8Qqjr2wQE+wqCCs4TkqecMCxKwnTdrjyURrp7jJQ
Lnvqbt7y4/yEW0CgqMQRf57jaMktMx+9nihctRqE4dNuIK6RcDKuFdvT5WhAy6SUS03nMK6DUbpM
x0Yp3L35rt+iySfTDIYxmNMnpzvZDN4E5kAAVbt3vUohKpcGy8nb2BajZmGzk3mQ1qqNYhMmUYHr
aTRJCPov1RGlxVFo0RPYNmlsXEfjkKm2PfklVq09WmFqlNPd9MKReTWc5P1IDV9AvH3GD8nrbm0P
4+coGRZJp4Mu4SgLtObMkUb49cDk8SMm6iCA/arjebfDw+cDVEZIFcpvX8iEqv5Fh3TCjbxPgjuH
mEZA+u3erozSyUbtkdMK9RszH6QgRTHn/so1Q0rq1vvc5xqlxtPqsTnn3yQLIQECKLuoxO6orCQz
t7wHXufGLeDlIbvRkmT+hJvYowrna/bkOrL5J7LE+rw4ikJyVafLswsMHsKBly8xOZ4ykSf0wI9l
dUA1wDUDMIINe9xvB2PCcJPOS44p1rbSjzDrkpeItANhjzGRjRFEGxGn8FIapInIbDOJCBre0FxT
O/ImQhePU8AcmbyO/TVYvGRT2orZ5iQtdnaCHPdRaRDxGPZJMFttCb9ZVG4mLeC7LFYVHcRDtoX7
LKhnC1LIVH8P6Vm0acZ6q6hKxVWNr60M3kzNmZ4znPYml/TeL491I6S2uxLEodeRBbfrZbStYOnC
BobTo6PZNzaUNvW0nMorLlZUCZGFV4RYKi6eYK8IAtwaxveF7upuWuTr1fjL5BAyuYJxHiWMq823
ffe40nhmKJnWc5EcWFHvibHnMiFIHdcNr8GKPi+HBN9jaAuRsvUUgGfJnkkPza8P40cajlFTem+K
v8z1LdpbTUcmwTGqGcHFcdmjBpINk3rS3TROIEzbpFhXMedQVImSvGfTb1nHtKRRvzkZ8wVMGKIp
uMO6cyxFOD9gABwIIH4BYjaHC4ihx+pXQloXqRA7XCr9kXRrB/6Q6bZBd8z90U3PkmBay+LxkPvj
xSU3tDqaaJeBXFJEifmzaxZAO8LQjG/Y0VXVp09OLlw5bJGtbN0q6tTzX9GZRZk9UBYPOQeEFPDT
8Us9SuTw7aNY3uB20X0JcEgXnbt6vsDsycwkI926tXSysva2rbpHaNZV9+HQqX+p9jM053y0VoNU
aAsj7ulFh9ue2odzcrktFISRUIbHGyb0jZrvHkgYDaY3NzEntB4URMONC1PBvWlwv4up3eZN6f3V
r5LX7UH1NUO0n3hr7mNfOFZxJNxq9kumA128TvaDI7jzJs7grBOO9zsc8muTLHlPx0Sha+aT8QW4
AL4gzd8ShG3TEgt/R3puur9W6977xAuCgusOeACqndXrDzCgkFCgJGEetNE3zuXdZ/9WVm140aze
ENILB+97WSaACnAmdWYNOXOW9gsC86LBp+db0Wv/qBGoQ0Yg1HpvFp5MXZubdJqZ+b+15roAcwO9
2xT0ppQkLtD+JPNdSF1t9fQIZ2nYSz9DdGsjM3H7KHjEGl6nxUkFaOzhrhES8YxBGjd1DoHmbpMv
Y7l3IB4MeENodY9zYNlze8dEb4dQwlm0IasBqSbXJvHzJOd52e8mtm8/Zezd/UXO9+smdHWbbzmt
gmPJWJEnbHmBZkihe6Nd8Omm1MFUEx1heI4YGkeh16IOxLEeiztQztMTPs2bfobkzQg4rl1uocLL
/gVMlccIkWz64bHo6+q93Nu7le1oyCv4FXO7Fkf+joiKoeuqZrL+A2ZgdJw8LxCWkAlaWZ99dyb8
NZXCd+ZmiyQYLgk3YyNOsZxR7jgxbf3IAobVnZfebWu7V/U2IBJw+81JoF8WCAABbalcSP8G3di4
pR5fNDViDq2qK5aH38BYz5se+wkEAWcRPung8m8gfav5nSbRcluJRscWm+A2TUwS1Vekix9wP2U3
nDOvjAvMAGe3+TmE1t1A093VKxyeBDuJ23IE7uxDle0K8goHG3aMgi+dlU1U8UjQmx3Q9X5oBXl3
whzE4ypko8MBrxL6vNv+f4VE2gxGapw2AG5zSggVL7g5ITv/Y63gMy6bTNHS+TD9QHcrk+jN5vow
yGvawpEJwVFkGwOFi9jgXsazPI2WYhOqlcswRXR8dx3ecvQygYkhbjcPYknij2ZwsHPyYAtmK+qW
f1JFvxjnEDc8NJv4+ZK8/lgIQXkcY35iuLjzDqB/BADh0RJ+zqtYuLAUUDMrbp3gTc3wVEaoqf9a
OwYHL4y8lj1G1KPgR5g0gYbTIz865vHwNoNsiWdrFy21YJKexz9j7kbPBdFBV9+a7wlje18uoats
s7Av6MsdQ16rIDR3j5KPA2ONU0I9YiwcQvOeTnIIoWq7C6TDuZu/UuJ2JrUbB+DufT6FIGYA0mGr
nPC5DbNLD1fHLYBciZ0rhSVnAN11AMO3a7pG4kFY58791TC4jV1256CpzbOh9DiliPQSqGQKiAIS
rokmj+XyCf83Z5DyOFpSBqH+HB7tttu8rMIvKMDWMGTSw179blcHaAw6A8Qp490Cn1FvRCwINy0x
/+L/KDPKKFySXbEk7acn8Cm6xDX8OX22how/BO8nARDiwzsisIt3FJwQ9Ot+CxhN80IsFC0cGAGa
oTuLcwxqpEymbQgtMQyEb6GlzKX0upc/Wq5wCpVBjVtxRC7qNfuhOzeMwNtB0bWhDfFZI+dBPW9s
Ax3rOqogCo6OjmuorWnQq1oTHfDExDku8bYETP9mhR13/SqO+N+F/5FXEjJ/Nu2OlsoG6HpTgR/P
LyRGTcF6commA4kyq8oEWvINqRI3OrL3Vb79g444E4+12wJOFBp5uvZMkCxdS278KQULkrc+pI85
CU96BjtQUpCFfVeLIhHIUVKcdfyzVhMh7chd8wR7vopPWWGLsHhbo4H27wXNaLskftlhcDAvkyU0
pv7idHBsfnEFTUjxxIWwutna/4azesSM0nIKXY6qBp8zD1tpaQfFyXzUy5XaseEVQ/ao7Qx8akoa
MZmVx86wTO0yIpZhwbznNulAq8rqFMy1kvLRZ/T9hFr4gJRlBuBJvYxl6aYr4qYySk2bMJKuNJ7z
TrOiixJfw9yHRtcrBt3SZx8LMOhryRs7HcRTG+weYU39/8moEg7VzO3TqU1svF6zxWdj4FdDUNNs
NX04mLTYS1L8jcgl9yHOdSzRHP2Bq9sX1375fAgQvH9dq3kbsJ4tvxABrYoFBcsXs2z23P2j47J9
u7mxJIu6M8AqUyyEGmcUqMjyghUmE7I5kazDU4ljx4XY6pkzpLN4HwsyP3KryljofQD3LsDir8HW
vJYfHjJUpSLSjy99r/TmLebi2NkWt3NT28OYpXsihl5+utYfbjXcoLLyzGYo8hphrRjxnmLLTruQ
ooIgLNDIRnKp9r0x0mXcSijwgt6kNiyeAUQgpJiP/ZBXD0yGsveSK3RIteUT1ckQ28yl0PrGTD1V
sdmxCegdztoimNb2LjfGecy3VQN+Bf2X4/mqA/cocYu/dw2+LkShZXUdbG0BpUlDH274OyWmZRuq
Qrowq3SK+dNDRhSdmez3r5DPaxPSVbyyi2CA9XAvkpmX76s9Kk105MuoHgVbPDEgfSemNrcOoCMI
4QtnTA843Y2GyQ0ZFlBc0IE3mQezDHFBpvlLDojnZxoXLaSHMcUDrVsFTDHjcT17hjEkvF/cgfJJ
aQKtimum0gi+NOtvPvF+JtG8Q+TCWGIXnixCPLn8RX6eAiQ+KpYoKBWLP/WypC/kswkVMUrozade
O0Xgk16dTiRSOxZ5X9g4y3LCzePFY0UQ1FggrjG2qOidA9eFjH3cOA2+3xMTWSVpJFXUzVFliYZm
yYkadIDGQ1URjihdxuNd46d+2rnInyGdclFvfwVSaLjGrxyUEoBjABm4ao3+hMWd+ZhpliORHvqG
cxzd2XYB9uOHXGOJZynS09fAZMDyK3VwCiXysvadc9W0p+Iktyh7y6o/KbKCubgTERGg8ScbfDm+
0E2NTUqUmUCgwxs+dLf7TDXJbJcG9cJN5satiRVriHNLnejXP7rbJ2sgo56YCIjgVERo355xRDMy
4tNFAIrK3A7q/U59MMNGmBWstJOiGm8jyvXg3fHti3QcjSv9YyvZM8ocpnHsFQgvdXQCsy61pkqt
emZAy6coukEG5Q2PNjlWcn0NkN6Tt3O/T7YfTpMVNyE/GCT5mzKoFyly2od6eRnohepFKmdnh6QL
P0j3z7aoOXNnuDh0/ZoDC906BWIake3H4PxJcNivsSNqFLtSjjWkr/Nh5YO694EyhM1B797Bbao0
Mio/bQSBkcZh6YYVBIL6uo89Xf/ZycPZO+m1VQy8KrZVljEf7bQkEeb71ANWVkg2/NJ2f12rZcVc
kYMlCUnzRru+CzJpyh5ey2/5+L11bdEdp6NqA3TGtZwvXnsjtrWP4LxmIvBxNIuDWZEdKohxmdJc
lzvpXsFiRR3yQeUbhzw880Ej00zilwfwu+WoZ4wvpPbrbSDPxtxqypovQeK9fG4uCtmf0NwrDyTi
I/fIu3QcYlvodY5QMYkHs41cLZL6yeJk6lkvk39LnUWxgD0ADIOrpKxi9CBjgw6NCykV0QnM30UH
dVGBpRBQ93VVfWmaNDw7IFOAZ4yq36756UqPEf8iypAaJAEMAKiMgcdGhdWVGY/w1ddWfSOXaiMS
MmsXhpJBjWj92MmvoxohYEVfZ1abDoICOEYCMWkS+1QdVl6Ml3qZJtAHKi0XSTfDfKSC9gq0SMhN
dz3P2H97qwUq6Ve0CfrUAy8qnUAE7hwTjL/VJFLtZvjbLSoFWeoHAMvbchWu2aLIcr1LThSNQTq/
1MmnywJWWP1bUEQggKSkldJCfYZMxE8cinOeQwyiKQ9iaQBBz7geV99bCs4lGmKZLZ9itVOCI05g
Tx1OvEGCNcBGTRSsmRPEcoCJEM7wg8ZiCa2lFaNtI8QrTbwMxmC8p1f+Xg0nh1HqVjquq2jym85F
8IsMwR8OQQABU/gID+8SpklQN8muWu72Ll5S6NfdUv0VZXG+mn2wQ36kqcaSJFTFnsFT0Enfmxp2
JFhCLoojHlfQrrv3LOrQ9KEGvC8riaLib15YHm6oYiXVFgL6zlWe8UyOczxRkIPMI+iKFSZLciiD
6g1aKCxPK/bXvXj0BZUH/BAUlHJZBZ05RQGuEip5lIQY3UhGoiIXtp2UdDZdaVf70fFBkHB4Cxd4
3I5xx4ri+UHgg/yHiR+pJ/K+A4XBYdRjFvEngpSlxCVXzTl5eoDOHA+o9c9CPMzAex1RevjyH6bc
xfWB38uZ3X/IMxmZIzey73x52d8ev9xta607JH03+btmo+xGOYMLHqu8UuhvvLloZMJluWXsP4I0
85TVE3jF5uJT9UL3GIs6t+V9ozur4xsqTg0YjEoY3TST8RBRPMJRTYH+3BPy5Viz1CLiLnd8b2e2
AmtHBQHsX/HTbVK7v2vCyXeYmzZer/YHDxWZCb4NOfnR998gMfzqOQJ4qGt3j/uXy53n1vcrEo1h
FluxXnOPFDeaO3EryHeiBPi8XldEowSo5GtZqwJVsMy5VoCyXNzp73WNMYLNuTY8M8lASI0Mr2ZG
u3d+bPiW5hDwll/GqF9IFP+XcrPcBJaEWQ86ob7EaQ+CyTs3+cakd3Oa8PGcCByfBZ/cCDTutHI6
nno108KmKw6NfKXETpXGtDGahrsdLrnyegEhc+m6RoXCRSmwNKCAxfkoGh2bQpq9TodopTW9anU5
OLQcTIiZDiNWzeuaidTzvDK4DdzWl6faq/Mm23Pvo4nXdQhkoj9fO5h1GeHjPsUekJ8dzJVve+jI
F2A29W8j5Vv+OppnX19e7/Eu6A7jvlDItJ4BdIcgm36L2/3n2eLtPLlQDMZlxobPuJTeCWGZGPiv
XHRT28CnvfzhA1I5iOAV7jqSC3EH31V2mPZBRih9wU+MUIV+eTjSh4tCzeO7hBswsx2YxfN1QjGA
W/OQweHI2S963Fk9RGpKhz6QfDkbNLu//IKMMmjlsMS21Y0IF3phBIrUb4JCKy5/6iyoQKwWUih3
4Kj22jznJH+idrGYmBxzVe4vBLwuqSxG27Ue1BiTXFsmr4IDVnSs4s6yejxmtKoftDtg0ohFgxFL
4MMtZLHYCxSecWvhTUn9UfUKcQH7OAYeSvxBbvoTAQvr8WYNkGbe+y3qmC+QAsrZnrPb6Lli17Br
vfmAkiYw9e6u+/UxL3AdJz4jWbcVniq4cKpPuCsar3U+11Y2hWC5SfcehgsyaR24CctsiXw/bRn4
IFW7u0p6Q01qA50PmWCq7NVGVcnfGkuDh+zUSLjmH0llWdrX/JmGfSH+LXqbtfGCUIsqBHBJ4gLL
gF/+mgkAsU49hm6Ibm3In+Eso8tfIAjAQJPVFb/bSXCZhuskgPtXlTjEaAx2vKdbVScDTMoH01z/
E72k92WFIKno/iG5iqzL2Db3EVDw9zlo9vjixLzmbu+lmmit7TuzlOVDJzMoiZBs+0spDa4tjQnP
G5AeEOqjEqFMSLGT0CtiZZ/Crp9nnDkI7EbH5ItveYYeM9jAPODwNwW9SqXDRuzJtwJruoTw8OCB
nZ0pid5bbXSVOAZyQM6lZszJZvgPtXPMoZLFNvhGs6lm5SILQXR3IgL0I1cW7gJKpOjzBxSLwJEj
0iaM2gEI2clq2eWsGxqbJ82DwCKBXPA7QhfZU2CmZloNDfYFvXu2BRllZqOqAmchV7O1StCyuhi5
a1JBEYp+5NJJQS2xRxKPV18YcpP0kvXOAm4D2xtGHSc+Dk55A6aQ+Wd4FxFs6spIlu4TwD3J2HXA
zltIrv288ea01fh5f8BmYT1r+VQTYNe0ZmGG+iksiEs5QpnJG9kMQv5U/rj6qMsxO9WUYePogB6Z
flS3gM5fKX2SvEjWXDfVIzvZ0koleeqwYSTiMlbp1nzmeeUvI7fMGx0muh0oGT6Tp/t0yt+KBbZ/
1RpWAnRQc/igqOp/rRDc2FRtE2cW2qx9rDr5pKx450fTMDZZjKb8VBG1Q3FlAkq+V8Y6HYsyUjia
zHnayEFimGGbZtPmupR1DryQOXJ1AOrHO+Iz9Q/jFWycABFhe4bF4yZPBF98IBMJUr+dffkv28hh
dwvMdqsT3HDZicZfGkB2xutXje3Z+zBWcEKeE65fIWLOI5ZNXJfWlh2F72YL6tTsFQBSdOXAgn/W
IGgvztKkfxBXL2ssPxAtkPXN/sN5iZhBW/cupz5iu65N68mSsSELfEOTv+/q7dJQYiEnOdfh/w3S
dz41c97755cQmlFgXgY2XUMlLeZOzSr1TfBJJ4JVae3Od7LUwXpLFvSBPcXzSW6XrgE3dvGjVMWt
Sf+N01UtLvvFb7p8mxCaWxJ/on+75CPvsW/t7rG/iA981i8ljW3wJ2h53qOtmGi4C49JaC7bEDT0
mljFDLdTjxfEbpe2p9zp4bsppx4/oVaZwCdUn3wdIVUGLyq0FbElZ/Ah5LrsnmsOhqWOsz8cjmiF
h0J7R2jNrPw8MS0r5MjQw8MQlffjjqGkn2Us76B48Etu34+TghsKxsZdEXYYqwnweHYx/X/ws/wl
DV0lCD0IroW/+wbPtb3skoMnU2gJvfRmyNUXiwmhJMxcSClRvtq7nciML2W7wk1tMbgnkLpLmkqT
a5vmvoN6W3V6mOY++eLenMlMDXqwlulqU2604Xl2/OptTSaAFWNXVxCfQ40ie20b3bNfA14ey/D6
8IQO7HfUjCN1PQMXDm1yLDfrU3C79HKpLXJeGNVftCwPWFF6FAq61ramjsBz3rZD1BTCo5o7EaQl
9sPeAIhssPwxs48F4ajT4gy3SgsztLsAuxdoR/sNJxD+FBLdV+8gXXCQxY7u6rTtd18W7RtgTUen
L4AwZhBVa9xg/elth/x62nL6gt667PSyOgaNw7iNceaz8ZTb565ngMdP1XEUhGNb5UElYSx8958a
Jn63t86xmIP9ms2beSV3A7Q4ARSFILUyHV1rZr04TCgspIJjyjFhuc4qg/A5mVqaeHRQtRMjwVGY
KjBDRLTvn7PH5wD1Vmf1DwqRPlsaPuSrVZKFuR3FN2pS72FHttIDrWfKzu2K2gTpAwaOGOGI7jug
aL9i2/JJfmL/IqcnAwGK6Nuq3ZOBusDsjG1yy6BZJiU6YPiTXOpkUOeLvrSwPdmbP/Gg9Qq+jBWH
OFlcEKbRM5U4NJTjZydRvD3LmuhU/3MvxuZqlL5wTXVXPAPL9uWQiFnm7McBElPoJRup+jKAjySa
KvnmCc8BWXIYw7nk2CmY4Y5X7C70nr1VacipKCKD3JfHnmLh0LiDeVmx2WnnRMRQU2swqqu9OK/Y
l55mwAoGCvA7Bd0YM68e3QIOSxJMPl6NjGtf20lDHWTdzS9dmU1phI0u5D2WMs4XnzEyFyzDy3BO
fpPKjb7xJB8qOWBo/QwZOSIfS2G/r+Xn6u7yvshhAWiMt3Bzk/PYRBTNtc3bvfhvhBZJm5TgLJdV
OUfWE4fzBNG0S2O7FrPbRTR4IG8mdcGKXRa4g0P9OE+oXH/sdMGXzOAG96I11x1z6Db6G/4xB3PH
2QCj4bCE9p2Bh20xj3UgmRxhSWHh+RKtHOI7TMxJUDNC3pShvwEmHOVsCV/1f0NBBneTVvq7o5nh
reHILUeKvohdjb+50hcCQYh95l/Pb72fonmt4n65amwqMaL88kzu/5ZYAwX5EyMojRm54PypdsZp
ZuxEoE1Bfh/L1Z0DiuT0myqDVPxaXIqBQlcamGZ+uX1uhwW1+QOgZvxilEByEjzFk2uTfmB8AIlh
/7q/Dj8VTOYfEnrwEKaH+yFQ58fc/bv2N5IO4VFbVHu7kwea1ym2IGxQSXFu0uTnTe1ageWhK3W+
LYW5LirdLjJP/nDPMx+Js24+T1WjDKdapngGsEhdZX9s+XeNLMA6d7BfXNCN2aPEqyc32/av3U8B
X0+j/6h7qYsIWPXizmqi6txPAINJSMtLZU7+T/oh4WABkPQ3y68loFjHuY63Y/QSR7j23ZzJHT6O
ursnyTjVbjecCNuqViOZSmFIAIV84+IWnxmnmVDLlXXcfFXKWH0op0SV8KxN+eDQz9hkdlFL22tP
9nlvfNJxN1tj8rilQMTTdNyUXafijjEc+KxobybO9fODVVZMx/WAwF1linkrYnkF1OKcxO5LZ8m4
+BvlSBEbcwaU9GRW+8hv9Wc19UMENQ1mu/8yr/eQrf8qivv8EsQeMW7n8qTGAXjCTRhoFcgt8qmT
AVbV+3mWmDvZnesfOYJUfcVOsKupBtnLD9lZPdhJXMsp3WMWwLuz6R01V3CXu0vsQ5NG827IDK1F
3NS7kER+AupyOrmDmbMGrfmAWqhw8aE9UDlTVuSmgYwpydYYsW+o0kUUhx9pffvgl7zbslvMLSD4
nAKqUtqvACVOXX0x4aAxcz5LYsQkKv00yfed0lbzZa2bO8BK9Tj6SoSJMm2vDj3BAyVGPi329tQn
tQJWHP7jBxGPvH8VqO7VfxRMJYlgzJEFtAeGu1ZXx9T8uAi1CawmOCQHxbG4Kw6PLoxUvXsMXcOd
3Al5FipAp1s5drI3II/cU0/52UNKmgv+c37Og2PHgw4Ux9Q4elptHcTGRh4V1+2h2Wav7i1mh1qr
g1uOT1kA/BT7b9sSo04+vKikM3+Q0sS/993lracexTUgFWbAYigqdUrNkHbp9De0PGkbZo3i9RyN
Rp0ZinJ6ZyvGRehLR2xKWBpxMRISiiy5xESd1wqyxreXh2QchTfTAwh/pARCLt5OyvJNn+AW0f7L
eXsk0BKvh6AfPuBXIHAfei6kJ8fd+Ao5xmRNrEgOMfgqUKsbDAeLjPPJSzGTRRp9kyFj885xcITL
RRpauMjOkrDuNOnsBkyAvMc8Q7vP4x8BcFECxIk6JHclHpexhpajFt9Sj+ycMBxyBmmjmwl2QFMA
hC7pM7QBW5j9HB5vIDqxCbF3HT/skkyhct5UX7gPyd7YIWSgVMuBWRqNdP2OC2DAPkLdMYg5zx4C
aW6RFs4rvsaeuAlDQbTZVgHf/8Yo/a1P+Pz8k+uLJ5q8K/DWJ8RCumOASgcOJ3hmagWo+L8hHfgq
D52eiYSiJm1CJ4SnmAkajCYJlGuoLks1T5/dTWftqDTpA26qy99MLhTwPcQAtWMZyvDVD8Q+up0h
f2ROEdaAldg1+0ZjYiXroOJ6mDo7WuWU0/psKg9kPX007mbxdPvMPZM8f6IS7ygZFp0iRbYJv5YS
84v/K1rrFZwR7DYHnBiFtxszqFHEKU9myP0sI3fge9Ru7LyUUkXNww3xy3Kos7xWgT4hiUFTHVoW
zRljJk8NxnzAwW3zMmPoDqboCc+MYg2fy1BsNsVUceUlcHS+bQ7Wt/RP4dyITzKCNgI53rlxuuBc
QlzipvYHOfC5iSIRvsvmwZfv2RB+3ebd4wRrLkteK6vGzKg2VIstaYQu/PkAcSKfn7dfhOqnsWzB
m4rBOxRhlKOSnGs4+j1JIrOnrj0upVZaEqRhcM/4E40+8WGjMKV01kXg2Kk6Y9mOq8LmsnDc3PBo
xO49PHkhkE/tpe0OMu4YjLvB9J+cm8u91STfPZfy8WVKJ2TburJowO1Ah68a6PaFYeWHzbTltzBo
iVG0qocrmZtZfh9UfsmgAnmItdRTMnY3z1d4JR1YWVTgVMPuldOUiOWYhev//Lw93yKj+VPocgA1
H6KVrsHtBvt1S3oLpdBgLZg1y5mxpQfb5J1kDU59B1JtHiokV1NwPwxFE2mWeFohqQ6cFGJqy5vt
jxd0MUUWZ+1dbJ4+MI9/9lu8tA3zxunGsVFlDSmm6yrLXw7oQBP8ZKNJwYIVIzKhXnAyw/L4JbFU
J3s7T+10OgPreFUMKP/UEoa59mPMG9+XdkvHpxnhEEKJgTq8f1f63H/bkL3DkoTAuj0hVLuljO6v
92l8TM0kMiUCNLDasth6jAI8d5L+YPkYyUrEXxc2pF5GwGyID4JGVd8kdeY7x36kHc+MveZzbvdS
38APGnLlEoIT3tnbQCvvRA95zg+ADpJCva4rqvLxPDF9td6XXzugtF2kmRy+kRj6IX3PKH2xiaFV
I8f5kAqPYS/wpYEy/UPJpmL1kALKrwIXJ5td8I14Gw7/BI3Wm3AOP9bo/+UWGirVVjia1VbWUqQs
sgOZ7KUvUhhVlmBRYFaX8mufF8tBa/qd3qJTMVcCN4AxGYYoT2CcTR6mjBHwwARwOi+HR2MZBLY/
ZtSZg8CRTy3wu0NCP5QCKk4h2+riTQRKAxR6pUobnYkqZYjWyxSTf6Lh6UevaAmhzHsv3UJ9ukYc
xbvLi0u8nUDNSvnp01/bWaPI5SyhgZu/CQtNulnGIGVPBz/Ys+3hzLBKYwSFuSCQpStIzr4fXtRr
WZhbHGVvLN7igWfLawGreytlRYCSQavo9IkdLVwSO1VcVx54dIQnpVvO/FJqU2T0ogMcWoNs/5VF
rYy1ByVJIrtswmxMvU8K7ybR7wUvJJXqh/SL9VyEx+FxRRiAWCyN5z5iQ4eGAl7qAVhI663IcmAP
5L/Z2UGUiJUGEB0zvbnWumrv9XaOpD/XReqc0jdJU+ljM6iinMn8x4DySPU4VNneq7QCwV9vRPXK
MpGBkEeQj0xjn25FvUeAI7mh2tAPVjgA+hoLUPs8bhp0OzmtIKsjj8feVon23u6A7CO7srEEboxO
QLjHZbyphe/Za053+03pQ26S8elI2zcLEk71ZQ9GOgydNDV9gx6EhgHMCxjjYEMpxyoiLREXbx9I
WcZs5U5ZFuMtz475vTgJCVtL6e3GoKdPY2brEMLNjMa5gIXOqVCwINCTj+h1FTCZlRzFiLqhg39S
INU1TJmdawFSTFrOlEqgdWs+CPWGX4Aw5RXmus0THHfbFzQht9/GkKiaMlgcC/EP7fde5glQexV0
+2+CBEXQvw8l6vrJo5LxGMrghfeZARN6sCyiU+WLfEHk7GyO0hJYUyETl9UYXHfvtIom4wWUqMev
1OuN03WjxB1RQRvwNwl0TiVYD91lwseuW0kRbPZ2d3wP7CM2DHqUZPnm2GJD3B43w+qLsKyeCnmk
Sa3gEGcDxTnXOYlm5ibqENz9W4IkaDgknRusRjY5+0ba52aoLHxJpxPnZDr9sonNf0GYK5lLQbon
PYibDqgOnCYTJ2qra7ofipTUzLvvCU78tL9l4f3CrV/1p58NSCIciW2v1sWDTW6LB22hT/IPrzzS
560sLEboJCRADB1grjGgvmGksclMbaMqyu4bdeb9tFcog0hOvM0b1p7ZaS5Gt6in/ypi+ifwkLpy
VUrUnC+PFbR15lfCQ3cWwM+TIQuGiCE3CMvxEOcEfXe9ngEkBbcp3CGyBuZcY/AM+wFYmdyh3qR8
utelkaGiRzOVMBTq2oI04AF2MSHmFGuZw1ZWqjt90PdU1kfYIYzDzcB/2ksd+nFompSZMYvGs1/Y
Hh1tLGQeEDzJ3VDYzZaEOr/pqgfdONjWVVn30t3khXZQfI9INTjzQ2A442Sgy9KtLf2glc1mvgb7
sSLTdo0CtmoLOGsO9UDmyZ7RRuQ40zRaHgd1dXgqUoQeevzeHTFjcSDe7BRW7Eici2jjDAJJq1X/
dimq+xPiijk1WuTE9SeI+lIbCx4T0C8vM2wXHj9mahj2J5uvONvILjiYS4Ig0DeFfExgE125Kz79
N4AAwVqqH+11o3WhSyh6wQel9/FDJeRxa802kzb9WnXdZam850Mmxe7qNmOGFNj63y/3HuMStstf
T5ZFHWXn2BMJCroATpMiPJlq+XeUIc4oYFYXdF1OU07FJdu1PdjMnlTn2F6NHoQHZQSWB7FhE/TT
293gKooeRiMe07SQl39kQnCq5M5I2J5iVE40zc+Ge3uga18Z3ICBlghhQ67isR24bQzhfLQTB1LZ
+EFjKBjPD7L0TNxA52RDl7iLeXOVtH7TLLu5HoTWOG1JnLsRAkHLUmeocMi8FkbYs0fGl6SA/okF
niqKYNn8drOoSVBXuYuq+ZBgCoH2++2O+M+qzZ5HaPP6gFWNU0OTqQ5kGK59tLewtLdwPQPkxusZ
teCJ5/RsGBiLfebAnntwJlKyI7I8L3EqR4cY7cYZlOlOiuUjnuc61AEhsnFMHIUDCoHCSR2oPeIA
TuJ6MwDXAW/kMFKGHhnM8u4aQpuhXBS2z2EN0XcJsx9vq1Uks1twc04sMoJfoRhRmqj8dVDYIPaw
6Y0A+0vXCMazKY6fwbnXCNfDcsQ7SO2h1y5HZuUqdPtJGQdzEv69f1cieJBeKbgX077QBg3iQfz0
EYq1JNIZsCdVP8j0NibdIQ3v9Gl4yqqw0+9WxtgDj92YqvozPr1dz0+0dXIMEEl86jwiqVtPj718
i8tsDHVFKPVsR5D03yywB2fs59+HHf0I2K48O+vUOMFHYIkATmYu+3E0VyKdKNAThkXuAXUgz1Es
aBrSZvDiXr0nZUn/xT/P19l9ta2r/gEBYxpKxAtXkQmZmr/ur6uti8+Xri663E4k05k42mYeqwgu
V3FUpRnqMdbDDmJWMvKIBYwvQaVH0KLk0tbfkKJbSC/7SRZuQS+affL8SCGK8d/cYOeN6HLH/99T
ZQ0H1d4ggBeyAjUXXOD6qrSG1K09bB9mWuggNSjuaDfxzlMPiRDN8dwPS/qlRQhEmlhNiq87L0jc
GAAOFy8dNa/9XGLhzffeXLag8gx9lV8Yx2L79kmTu0EI4vjyFgrDYBqTpzVdYv/GgkbBBd9H8OBX
SfOVr+zzUtQrJvSoNuJ5AVnEH86/o8ouZlAcKlx9SmoG9muzR20nG7cKl3mKSVqT7S1833dbB94X
sVtG/FBbLm4TVR/RqUYuB9QF3ZJRcYYJZtijr18RRhOhhkQGXfS5D1xBdNuajY1A+eRPZO0ip6TO
bWdarzofntQg4SBLrUR0QCSjubBvKWnKmfLHA9U0a1IVZ0gOwfncuTITomt7pKzhABzPJ44Bi9Mn
czGaaCzzQsjZx62pa7v51bUni4rzBwviUrWAlaHxy2sHHFOxgXAgYORT++LbsezwLRU4zv7j2t+Z
fPsdxmdiUbTnlyIZOcCTD1Y2Kiq+zMtg8ztezrdxrbv01m6QyOSFf6RQI/OGqn+MbvPebU/LdFh/
6W+0fWOhv1tLL4VVuN/lVqzJOhL4TdXDe/rrrVYftUsxesGtIC88Tm9BEKvX/uEQy8Xr60fRy4/K
Neo0d+5SAyqCAPFw1E8E+j8hcKpBvql1KCP1UxlzfGkMDPnow9nGJsrKRfOvmIYwc5yJziRXboKI
IP8/A+P0xbWVoIycpaZWi3Nrxd729oDa2qy6N1u/XW5bodAaBRPlISd6SA7QNP2dIuqDn/nhaU28
yy5exmhvhA7UJtfBPTcvFmYc92IWQ5yF6Gc4kf2Luf0jJvDgzfCWChS//ECatygYmb9gE6qbw5MF
NJ5d52f+/0f/8gpm0C//m0g/1GNh3jP+45t2FnoQ8tNgvAQ3YWTwW0UqFBIfkiAF9PZ7BGrTyTz6
iz7oSfKjnN9mY9trMdbhs4vwfKdhvDR3VL7MrnUql4y+wtTLY/yRv58PZjiBrNHYEbnoJhYZr3b2
OxIeUtxCnegEPt5je6TqNMvR8kc4moRMP6pYkeQTGGuGB5GQ4PZr3iHNMfbUEbtYH0vZQQvxFZFN
gQjZGOL234NuG97UM2wWUdqPk1LVr4aXJe1TDpH+zCF9AcTlS03dyjwN7i3bpZ9LQJAq06Hhaszt
YLYubodA7/f1iPer4NzcG2zy+WcjeKoS5aExrZECVhiuHOANpKC25f1Z9xb89sJb8xjZAZ683wsn
4nUdP9rZU7wg8B8au+u3xYxdnEq6IFjtMAZSRyFJHaOiv7r9+vUCOxOisz6JIOAMnBTyO3EWhQL9
zIQOoBl4iP/mMFBLaQpqRCEyUP7mJI0xSvGLI3tBoJ/WUKk7TBnhW9Gfvzmo0d8+BAqF1+m9AP6i
Ip66gqsXRVu8Kii0It+dyuIMNIPdBGuDDxmIU8RVYhqdUl0uESThvajp4TijE+Dyawm8QBj78UlN
4tmd48sCM+D2ZN3oFeUn6xVeio0sfas5yJ/eg59lZLrWWHoWdV78CHIEwVCjKRU5/S5cNaaHBPDa
fNd9XqVXP9ZLB0dXebT4NXeMFEktz03Gf1SrmW2c3+gSQKMdFNWrt2j2W91ex2wyFCQbCwaGkMBZ
Xi4RVfJHtUl+3xvRts2VlQ5fJXywnQmbBS9m9bJYU8Bx73nRDhHZS4W3s0onygxCqWXTQFWKMq43
b52KG1r5bLnlBLC1XKNGmJ6JAP06CD/B5p4OFWd4UPAE0d+4bghyCQZYdPkYpRGyuQZkJ+6H2Qj7
D4obM1cuZz3PF53ouKmyHf5S6tL7saasEDQE1Iu4lCP1fgz6H25JWmipVosXRkq9Y54gIdyfTuyx
gn9LZvLyr17bMa4Vl3zuTGsh3IzRj2qMSOLVwTvbuyLr1fKbQr9q3Rtb79OHyZWRG+EOjXsLpydz
yoyOzGDgicwS5nd7ey0qkfcjGZxtvtq3SPgdWMCWlIypLoXd2gcFtAM890aUy0m0LWOdh7Ily4S8
K/dlzGYRlmc+2tPweh9+j6So9mLZxp9AC1gQ8E8o8uN/K+2zSeYsvVtCC/KsNBAy3W4FPJpqvaf7
xbrfc85XGBo21RKcd9tjKD1uZNBKMcJTS6oyTXxEzBFPMQ4dhvZpDA/B9ljZ113gpiB0tkdJ9LX1
jHZ0b6PCL/Dfz8QVa4GIbEDzgXHHcmx/s6pqqG0uQf9Hh5knnpdEX5UtzKKtu2sit2ozKUSaT2aS
v8OPr7PGBRLcXgcvYUPZGsZr7BjPgzndDRuu0QRC4xDP/C7GeljGYyl/feiBFRnZK21Ry9vznEnM
fIlOIyVEjPds/zdGM9Vkxc8GaIf3BsKmFThuBC/+CUeygv7M9RBGGgsCnLc173ApvZM7fPsubGeu
lv/XDskW21fEu2GCFSmbzuk8HYiCKzIoD6O/Azl53z8eC1SBJvsMPeWGJPxg11lRDYec8GVOjLfs
u6NOISytp/cjXFS6MutPaFPrLX4YyzeLyyl7E7NvL4A/0j++nr5Vv0YPdSnHpWpxTC/VWH4Wa7Sd
xT3tMlrdaUsHt1SoEw6Z7dBhf+wPTU/mmKciuvtYkyXcQKZuFTx/vLqZreh0Guun9MphQNl/pDxa
9qy3BnEhkm1SkSjCUbGZMsI+uTbroYq/WcAyaO6S8O1q9yCkFHWjJOd3gJOX2LC02S73m6znBsAK
4tqQAZFM+A3E74PTzMkvxW+2xwbCpjc2wPrpJbRwTAb+3aCb5N6X5sWuWK+dVekmfUnITVHBNlcI
SC5DFqA4Hfd6CTyuzYYuNBLEks7o4NxuPC/RdLpX47ueT8efg7hzSsoQNqww3C9oUv+zGo/po+bR
3a0I5ZuA390My1DsJR2ExuQadvoIb0B/kFWYaTAC0c+Rgsq4P6vT5vZoonG7QEK0e7BbP1zRZDUq
18dq2eLO3wNlhNFDvsBburWJFFTdl8nHYwNR0J9oG8NLm+iOei73Uioc8xDyYgQB8je4/IQ1le3K
AaukSfSNLrlzl0wurRXBAvk5axSxlysrFWbRYB9u5V+Dn5nGLt6wqMJaPQ1F/rDNLEv7Z/ZLZTa6
TdNcTVvJ/hZ0Kmr7KsuBjo7i+9WkaQ4+hfNsuT7+7EMkwFl2A5uQd5gEz7YVIfbixwEcUI6LMrNs
QtjfEi1rdzigJ7G8OPioGDh+m8VxHNqvmmIsW38kHo/bgB8oHMeoUWPrA49mf2Qt7x5ScfpbNlRH
UeN7sDlfpXRY+SSQ0ew0cLbDAyScpncklg0Kw2x/Fwvz5PBZkXKBbAhuzvnyrVZW/1AxkkKItaFC
PtpooELc6g3ZXWSBcAif5ZK/x1yJmmTjmAjDmxv5nINjuKpXAr8kApjOatH1qkVrSp3fN/luDb16
CR2JuKB2Pz9PUNcRxN10yKv7EkFa0vjm02x0nUdhv7Vf8KgFOUL38Gajv7pQ6EzPIa6CW8EYIrQU
8b4L0qDhIfRIbYf1C8kW6wmgrVlvlGXLsTp/clE6IGQULbMp1ueb9oYzfui5rdJbrG1ao8I4Yd/8
Pge66QanQc64agX4CfE0DGzZt3qHvK6mTMPK+fgzOywNnexfA0dna7IF6cM/jhXKFXRWyzgHGhky
ybD2nohgABK8iwdZ77NXTfgug7p2rgamvCcFfWLQuc5WctybaOsrl1lNKJI2u8mf3ihMAtagxOKt
lKnn3wuDcbSAotrkpBVwAAOhYLFBu3L2ry5KdafiWva0oW8EZ0uCrYirZstX6Ox4tloRWIdawpve
jWQuhD73A4x2SgI3OiE3ijy8G0aLWi0lY4MoASw/yAU4oFkV6XwbBwDY0W49TEtX8zudpzT2d+rO
A24VqCnE6jy0TbapfHkxCgtDGjqvMsjTIUilr4F8V4xuLVhqBduTLAIJS2m27kE7Xvlqw3XjkHDp
nQGBltRU1vGY9O/tqkshPJiY8zIDs72HVCEAnKEkPsjWDSOGiHjnu1A4NiReUWOYo7w9H727jdHZ
/SxJ2lNmw8SGAyPmxhlAKoVrPG6A5Ba0usa5Ww67pMxxeGJTeFcJ6jVgoKSknI/zz9l7pWFrffgk
7gF1SIZyO9MgC25/5sdQ9pYxASlbvk2MscbrSlFxSkkyPckkrUmw2nyI/HYe5iUufI5flaSzBHSz
5hezU9vnvxCA8Q5io79wnuItS7/Z1V6sfVVOiurxwoauCmDmiCfmduDgSrMMbWuaGyB785r2qy5N
vPmlk0NkUqPmVEhUbOSlJOGzHzHpMc3YWK86uwyfSnr2mlZsLycWvA9O7preiOXQ+HPl1zCHAk/4
NRWkP6ZjqIMNPp9SRHHsMN8Wwzw/Q1JBm3/gdz+7fKQVgSiq0TNZ38Ijmh95Rmtv3kGD+t0PjlC9
EevE41Lgp/Zbz3Xj/XMl+TnLTfqaJGdVu2AnQwfP0DR8IRowNLrXM60kmZ2vhUOxvOeglwuOk+lM
jkoXwEe2ZSWLBj2nKEdvXNYMcTPEiapFuKJrYXqktZaWr2QJY4EBLceqhM2lvTJ3PqoMr452fQ74
cmLREotgV9qNfuUQ8CIPqIrPZR7zs4Lb4Kd4TttO9RIOFsw91C/nzrvpwmLe/zpzq9kmsxeJanxZ
c/XSB9rw+dg3NbMVxaYU2kxf/77CsNhZIA3SX1oKGbDIVIMeb+PbxIPRZazu2KNd6dRP0S52g10l
DOvt4pSd0bbRh99pHkAOv0HV7nr/dIKP/ofG6MhJXOLeRIxcgs5skG3rIRayZaikyzNa1wDXeq1V
5qHOd0q7ZmvE66CfkT+dEl9kRfV/NJmi2ArBxRDl1FYE96hc8sAYWwgiedL5F8E0yFkNdCqXmIRU
L6HivNW4SMwcN0PglnkODB5/AE+2/2f/jm5tToQNlPJxgBV2L6iQfR5CpnIpBXPFbQXy+VgzLbol
nrkQh8JsE0eckKnzQghrR2BTnEvMJaI4ShpGdNIv8n3DOAn39RlnI1habZxCuh6Q+Zvh4xBioiV9
yq8uxRuDSdI2EKKs/UuYcaGyhklaiGZeJRtDk6UCzXuj02mBrrn2gmMEeDQ9qpB1+U//wZDdvvpt
CeK5bIF88v2fTvhFWv3062Rqxny/FjWhR0FDVWmyppcldI2v0p9L+T9fw1gPAJ88yaGPCQG2YP7V
7ZIFzqk/NUIJTgIR8/Upqog0dwLt2eUEXOnfgh/Xyn/2M/SeMYgXozlsCqMwQPjSackBo+uBF7M8
mZVIV/tJ68fxaCQ0GcZ26Xq2eIyG4fP/ttHQ9QgqDvmRAlwGPr4gWxUgxXKNIelh4b6hGn6+WHcC
VLVr7zNjAaZ0sUeM7GeKdAfQi/wJtSd5fBMTyiHL+4FFB3itjxUK34VLNi16KiyTjgwNYnE46dmU
yf/+pcKUF/vzRfBT6DGycqvIni8MQodnuRL1dp7VXlhOC9BaKG2ub97qITUIuxT1rYmf4OHZEKs/
6dBWkYlBVvydmUzbScJdXQpyMcRenv60/kStdHs78ceMy70u009H1N66+5utzAZqSjRbAxe40juQ
MH87prr1K+XVOKaQQqPLUlwuFl0QMX9coe+bZNR5xMkqZjFV1dwcywzLTkE+TIqp5NLcCbTa/hqC
xEVxS3/dkK0uGHdmoy0fDV54D+4hGvMfZ05CmS+myb0TD1zeWIW9ClqN0V/3DpUGzoQz5B5cdR/u
CcTW5pk2EJCS219VULvsOIa2QaYYiiDMNawFaqV9EOdZU5yiUykQNjtHR/VGxLsW93bZ85YEgY1m
t6BiNReCxm+YHNsBlveZ6o04ops5B45G2Sn9TJ4XQe5SbMbRbdE/iuIwivw8tM4FzMDcVkvwcjvB
86pBwFfVn7bkAV9uKjqrtiBgnmUIpdTCxzdDwdiXxAfEYD3DPTi8r5dMeBHOEePASKoythL4+S0d
EO91VBCy6j6BoOIIyPmC1tNlaPQrmqjFVBBj0dxjY9eWcr/oEHnd1GuFTjxKecbxSiEuhkaPe1Iw
JHTkoS7RdAPQVbn05kPJDwPHFB4ZqsM8iD3Y+sgZXikTCKoISL0Ifksou2yAj94svtYNbmFsUTFF
A15QR7d4UKZwKtDll8rYw9MX6Q099gUTPiBjOrV6hs7VclAuE5V1Vs8YTZquCrpyIpbzkc62G3ZK
xzAcoyvTd+zzRIz7qlx+FIzoMc1RfrPre7l+YB74Tc65F+UH5e9RNSXi42HrM0MBqbgsOkyNOoPl
HWHQspu90H8K9wyUckPKpycQqAVXgTpkmeLQ8uwLZwZG/N1/KvHrj3Kuz58c9reC9SSRXXHprdUt
N8hcoAUcG3axqShlOYBCvrJMKMIfe+vcZEex72A8Jug3mKYq/ElmgX9ySCW43V5PaINsteVRLk4Z
bovE75XuUbFTLOnJUpyBsoydTU72S9jn3PTZccbH3qFhavURcZyPXJP+yNUOiHGC2/AFayRDveYd
1uumRXBYtf5kffJiZsZUMM95cGyMZNYthG6fTald6Vc1gPDSsS1Vxs3FVmguVupcQQt4OiV4GyvS
AMnDbJBgyb4UqsdNPfFqkdfG/bbzfwNr7Kd6Yln8Rhnge6ENZOuP1lwBIfwB8XgnGa9EEg9mePcO
6a/rlWxGt2G4hgOEzAvU6s6jElROh2JKR8R1p7wXcN4VgoHbK5rzJLqQjbZtXoY0gbr9hiYiVBrA
4LEoSLVEIl87oPA79SgMYFx+i2vWsO/C/mtgpsU1CtsKkNjyRAUMO+q6ROQXECQu60/ysKhn0lAF
eevb8bRWBzaH1C2fhu2TzqcK/V09DT8RLrhRGYBH0PInhWBvrasNAxic22fE2WYNcFOvyvDyCiV0
WndvSirjYNJVx2GY8+X4OVvbl7JE5FwboNhqzDXpbRSdhmHWNRpeKSvj5iobl/5lWe5LVOUO3W6U
D706vtmZl4Rw28sha6ocjcn4OqzxwbK98fyEmDLAmVD1P0j6S6bjGrYlq2Ru37+c4TbJJt3zWpQE
D3em8ai0jFpC/WBzakzw/KRsiPnqJYdQG2k4M2tfenq1pOy+MO4LNXwz4GvTRu0Tk9ubZxsxb0KE
B6z6OlOZJU4VqY4eHnaj4t9cAuolGgQE4+5G36T594B+g5BSvZFwitwG0Cqj+F+wg1n4/kJwyPJH
HS29zz/0zSiIz0FaT2iqUsY4otaetsTTfhML7bzDZWt3tbHlF/+aPHAf6gocYnCNjmeZYombOiVi
fM2lQcF3GGUZy/QEg37tKVdgzog5UW80uEY2i19zs0wp9aW5T2ks0NTgpskTLUFUgaFevpdNkM68
h9nbsiC9T9S7tBzsIJgyybXXy5q2i/JbfgRt7RzNUqKpMCocA1b4seRI+Q19ANY7A7OHcICkTci/
NRzunAr9qF4Jzjcfu8rBa+HRbgPJTTeDWJMJdbZlGz73vJt+O2nS6z406XlxN4/IwNJeUDwpOj8m
HRT40/wxk19edl0IOvzjaFe0zkGg+QRdwEInJ9BMgxm+8+AkZ+8FeCfTdvrSVp1kbyD0fR0iMQr5
oGrYgR0Xsxv0zJJ8IG7xsedHE0Z8X47QGJXz3ChESyM+Hiezd5E/US7jKvFyOOBJ2CcHThZbKkfP
gvTHPJtRWp1kbOunLI1PaycqS89fA4sXd+G/7utSJ3kXoE2eOXVsQoWwPrT75teEeaqlfjUSI7Q2
FNYq4RdkbmcpzZbUY3DSjowfFZU+lqtZtZtwgO1rzGP8BlEyhA+2Uqot7PX47/iod3hfmtrU5Tpj
2jlRCXPI4PI0aM87nJDPkvc2k1zD0gLh6R/UnpryVqRGhij1goaxpAKJ6FirdGxp3dBm3kjVNXOt
pOCdmC1UTJeE47UBGPWQF8NNhxp2FZN3FpObrwAxhIzprJfUVuFBoUSAiikok1WnR9xyDEEXPir8
QNZbbm2LffDo/pxaoHdjfNpfblPE1k+BhUdGzZ4mtRXYNJxcAVBEm75YiSyoPfilVmy6RNGNSjaV
3GKhVZCZrU2TqfJFKc1xEJ1XFKDUpI6harqiJ8P7E2s+Y1FBw6Qau7rJnTpiwyq0BAXIOEekIM58
c/ZBgfEAsFI6SWX6qMqW5mPPky2BocLlheKE81ogTHbKxHZzeCjnJcfQl/rwpdzsDdeuy1P0TQtT
XqeP3fWBUsG3Ve4PlN72voQeNzXWJT2R3t5dLH2XSPxnPrd6UyLw3jo92i3WVJKzVqblSc84bgME
GI3ubJ486r3KvWjf8qLL/7vQUQTePKIXo/Kkf2+4bSKgkmJFGhlywgqZpMIwJ4KtJ5MZ0NZgLVWw
FkXPGzPMfUpwLnvr1P9WW+R+twd+nTlJIwVLBoNVqqng7QGn8Uztm1br5a1Hwal8oKGtDScQlwf5
tzGUSzMd6dovJgTlX7ZpJXczOGc59+S7VtrDNSWCQ68Enilbu0Xn27AMgEuZwYUVCOj8m0C97cGJ
l06bNd5dYljbACnRDdqjWJgBm+8kOBWj0RC3tr3XRb42fOOfbudGFBpVYCRUKTpAvjHtJshFX2Uk
WkvcoZlYbc+3HL0+4RT7oY0dLD8c8j4LkeA6sdaKGCeSmma5np/ixtU12S0RrSkp910RtEUXc/8I
TvsV25pqhUsOFGBZitJZCsGwLnh7hM3zb3RlJw8dRRzWU7SWh0zH9Rmwhk5C+RIG+5Nt6IqXHaWg
JOfqcEZBSXUUAJFkiP3R6jAd9TH7rjdnXZtUvDrcZwYnkC6UsPuR8pumJWsKBtefdcoArZ8a3y+K
uT0jIZyGIM2omMOp3QgQKJ3qf1BbP21EojvLrpl/JIKqKAY+lQlfWmvp+86RBDUq1yV4EtFI/c+u
rTMUuzpdrOz55bTRAonFoRJlmCZpD0ZUWeeZJO1F6HCbzORdfRjYGsvWhI8Z39J68Z4Ht2ylAkyD
qF+3ISpIRGhIwxUzw76GJ/9ScrpbiNjAQkAAxzr7aQYk5b5jDTMArJJbUniD0oMklHDXtvri+09J
0xkcv+qJkCoWjz0C6uqAJSKTP6u8k3s3KqHKvuQt0GKrubW/Iaa3O8ezH9SN3eEDlJomc2MuEYGU
eL3IjVeTlxfP1W+jIRi2kLPaWfKDCBQmm134lQiRqgyJ4Z/rbZ5cYuHhHOY78PhmCpcP6M/SYmob
Tr/ByYj/nwYqqAig5W/1pIBe1P/pz2bvYUDFTykf5iiRKeisy/O5OqNKopqHFf5YXrVcqYcWGFMi
UJaLjVFM1VwfV3c7Fbj1ze4irkT+SIX15zGxeq+cU43nR+Xp89VOPijdfwtX4hSkrkqFOyJgnDFR
fKEGglV1f//i2GcZdFXrDv4eq1/uAaL8MdurhkGKiOTgp0ZiptHikXcsBm7rugpEYOQK7THlT91f
fJKqbyJmEcolRFJ9KXKXwLMM5ev5lDMkmmQNtnAg6dsqN0V/3bmGwmIozKOcVsUsBmMFGqqD+AYc
XIH2daUpGwfNAxybVwTRpu3xwZhwNVon1zG/AonhCFtak3OgjWr0rjFWmulXKvTKrn6t93pDVTWg
af6FBgjOichApsQq7sXAa6/jFa95QOs68LR32YDhOTDszJn9LL5pPej0WinAKZEoo17gEUNJfr5a
Y53DZxOUQSadIZ2rEZg5wcXjhyNEFBk90iDQwKHbC+c0oKjT11Yc+JBiCv4Cgp6/+x6f3ncixGRb
Ggb/fIIqPv9dwclzsDAI6Zs9BqvGupCrdc40fzGmhUjlqlBV7ptAGgLKKSVawk47oz4AyhNF6uP7
z1OdkSKdMvVJzJqdyZS0dXxFwphL6klvSRwL9QjRDGw3D/+9eoD7XLi/eePKPpaiBKyNQmM60sAF
Hvl0MZUJFJi1mOpybTbeV0bP45HD9nWwGVNV4ve26PcUBOcZmfdKOSM8nZTsqb1EGB6KeGqkXNHQ
YN0JrMuwUIJEi1TxY8f+69nfvpHdiCrRke81ZnexiKClFTytOGrEG53PdUarRMynNVRJQhhfqw1L
VRdTPIbnWJGtko11zXkp0AsmqMKUWhaAJwh+SZt3rswJaVLH591/ze+v2/IzdT+oANXl6XTrKINM
9aWPY6s3/c+bHdJLBZUUsTxXhzOCDkHQa6rNGEBlwwEbrgBC+why38yjwYprPGLuY7l48vuQrQxp
MWw1Vo9tV39W4HPsK+B48LHpZmGwwzn9aIneLzABNyCznWv03D/+UfeMQnAWwh6lj7FzkERzSaTC
UO8IPmgyeCMJ/07n8BxYjpdsjCwlnBCp1SGBgjaEumbTO05qOKNEE1yOE9VvGtJQ468ub7fygWI5
nIJtw5gzblIApQrmFXvybRhTnAlosaXbUlZP9oRVmS2VE3YCgnZ0lVAbIg6ZwYCC3i3dnXeSxlaH
p53mDRtnF+VXotCaXHxHzTHM+E+u52LGyOyr28etPI+HZKycl/G0mRL/mitlgmTUTBDHt22JvDqS
SSfOPNKAce7QP6ZFFcVkq9hwEWJIiWyxryGHactLStVf2BVuGMNJsk4CGA4rp3jUGEuG74a4PN5X
2JsSeFjOAhgOhLUNkt45EwBCP2sMX7E9iVGkm98/UYtxICFrBeJ5ta/MYFYVf10t9GBXhnzlnVRQ
VLgN9IYiyrAeX7lfjwCCXO65n3P5P03VF2rBxdpBbTTrM1hkLBBzit8i34bHk1cH/Is585NLjX/f
ozEgM8DQJhOeOt+IFl1nc3epgLIJkOR4U6lrvl09OL1X73ptMuOzuADRsiFkSofvGm7EBGEBayaw
mg80UXmS8YQFn/CGefPVct0Q+XLTl4hYS24Z4Xcga861K0NkP5z0oFNxeCCxXyok9OzvspUlVIzJ
OcKdFIMN2f3N2rX5fj+5INPmCH97y02LNLXx+0m7XdKsf9v1vQnUxAGywzBR0tkTICU+IXaqsDKl
gfbH9wtCjOVs0rSxfODkf+x56BBo5ZaKNyFWfuDQEWAfGVwjz6wSXwvcShxYUgBMp6N+kHrd1fw6
mzJBBhWI1sd0SQVnKMYbHrUytSMBr+x9kjIozBiryHta0bCnkXHlQSiJErNQG6zmEVPXV1+im3kj
JDKbfZonmpzE5q91Z9Oa+eOyhsRnj+nTYmxiDDzW9Ah6Rg/WiBJKfMMcPsRUrQmrVxO73pUvariF
dMs1I7sJfp1YgmuS8HlKdSggxW6ViVU/9/uenAQwyVLESpgOsS0cA8yqpWcU2iAbHMJh5ei9IOqo
EuItNYXuMqabJf2OvXkwAgadmnnP52x99d8ueNt+4ag6gNJY2gCfiZaAW3n3D72ElUZxF3H6Mtp9
v45ivcHbLYrlMSxcJVzzNU5qZinIoXF1om7qe7IL52xejhktvVg3hEzKYPlUCindtGhToVnv3Z60
hGqXKHTll1dyE7aU59n7leigla5MVjyYSUKmp2bXvRLKnSWJphq7Ov62adK94f/8i/3PcooTvMGH
JmbtjUX0+hT+hVoQBxYcet3C8pM44dv6AUSBaLc4Gim3QWcasCVzR/2VaeTlqemOe3NRfrYjjQGa
KTLTyMrSaRNK0Z2odefBaVthVxHHtU7Rc0zOIezEJyWPnmf7UeodgtT8uSXIcpRX1skxbpCjllVw
85o5GOLV2GWBCea5F+MF3q0HwSdZWl2iombClOKgHg+dlKWGN0WMMDdWcunno325OMe9U67Ku3qL
cMRWxcysc/shTrNEpygX8wSY1bIp+WVSwoUco3Bzo646e+D2x+8FodbEGc1vk6BGk1h5YkI+tgA0
rD3SOKm2aWKppxT9RNtf2VPrGidfnbWhraNzQ2sf9z6sbXbqA1+CiWSwbtfxeclBXrapt1a85SjN
epcDEi2sxYe7JQJu78PPDgzC3iHonJ7NtUVbOveaPEgZfpqPtRzVPNflX4SvG7hBZATl2wYYuxeM
/ZlIYqqlDlZfeOGRSMATAxgVubpw+BghSSceN8+6rIUE+0a2z6xfxh62L7O28voXEHfumtsQrALz
E4XtSrtWADUhSxKJuebuOBpZtjGwh33afc3hLICbHfzkQ1NGFfJSHyAt95rREBeFiV9bilnIlEk9
F8nui/7Ae08NUCmGpBOVBTazrHo0lnSsuR5N4LT8y4tKxmyddEvbtQthYYdUtfj8KG4ZJYn2JbFQ
WoloQv38wtgzEWpl2bDiVPmKZ2N79F+AtoKBLphAQrQVheLgEsYhZAsmkOYCFay8lFL7Dzt66C8e
5bT5K7Y/sJ7Y4RvSITCznY60eDBKLSMhFElQBvxtJ8iGeYzv8rkv46hj6lzxWDcLEi34eDqWB6TX
xvjTK7ngEOVGCvADcnUVA2Xel9aqFpfAQijWYr0dmV4znQHcTuA4jR4HewSnVp4X1bEc122o0WlX
d1BaruJ7y42H4o0zyxrNUxNO7EriC4r6xy2A59N69yfW/TD7INDwFTqOke/L077ekfMjy6R9mVkV
LXTzGySAPGNwgJdB0SP5jSe9fbqMC3J580mF2WVetoYPOFlG3EOFFZ6uZtW+qxNaNXrv89tD4u9c
7bjwMbMy8oZwh4kqozwqlwwpLaEDqt6Aa2EvRa2kyYEpkDD6woCPiMPG40Oxr/K/SJi4Mag54GAl
0GiPy0ucwwhVjd54Lel8UK8iZdHPqCpmc4OmULTYebVYObxi0+P4r0zPtqUy2Nj1vu48jnCj8OyS
0eR5rWEBDJpJoGZevsKqI39Z99ns/7k284BuVXtO1X8dC8B/XQEtiajIlS1zzewp4uBQy6KUWeup
axaduMnNt53x0oBjxhVdJAQn/qE79N8oNHPgvNI9/MVONs5hSvPa5s5xmr1jCFovY3z6/k1F/EMw
ePRlvQdxnOY2BMqsMZCTdINBsoxWFg89p+j5GEjXkzV2vra4m8/1uQgGQGrZknjTI8IthrJ0Qegy
2ZwIp4o2DEIbb53dQjGipLiXOoA/Y0kIcfLPWmaY9P2Oh/7B4/zq+wO/p5SEvc1B9r6zf2FNDuS+
uVTD+wO7oZODAsXUNqyLS1vgc5Ao/iW8MtWt6lOIkIsljqFYPLkXAgTgLWMgAMzEFvsxWXfLkjVD
jgej3g2eMOJ9qud2iMhMswvZZunJKeuRH7cXFEUyPG23b7zUQXzAXBVIcF30rEA9GZps5R9h8f0E
3Iukt8iBiH2xr6Otza31tFUqTpaXF9vdBfrGQcBKJ7Q0iUPNfbmhSIM8gRxGSD7XRBruVILlXrFA
oKzEhKveZntM+Bc7aszgqoF8fQPJIrfUvtVW2EqE782SKOazKuwXiNGZcqf0jZb1/pEeiyPAtTl/
jvuzcAKeYN75MeLC5LXKaXI96YvdOho6VvfzvM16aY4ufFutjx/cvw0UAfGPZ0sgvjmsqGF6JEAY
1WpxhtGW1IfMvjBmXTDkNyFl4t/ya1Hl4v4nFOjejyqZYMvFjp9GCofnrnDeMS8rH5NxrvQZAFG4
S8xb9JS2PY1L/kXnxG0gM3Ehy5OiUkF9D47CDzdgQYuq+pVQe4ixD7/cbMKNXM9Qf3bCRSNl4Hsc
E7hFLAstxFOqAXbnpbtPN0rhHk9YTETe2gMKih7AIyJnwjAcDhX45a1pPChvx46b6zny/l09LDYW
Cu198maVAdnAyZilCaRq3ZwB6EkA5wog+q7lNTTyZBXPmv+u3vkstntOzjKln0Jaer2oJ8yctDtN
DrPN0BtBYTa0iWVkydzSQWoWAuCFQTdsCyxPRWA4hX4iTqI3dE2rUAPx+yp+7BgMT0YgfnO/HhXs
wFuFiAqfR6c9H3rN2QYhplZDt7C0lHx+W9JR5mbBIR0G1gzYQjaqzNG0K6C1tccYSnaEUD+/CFe6
G7fsGD48wyVGunU4Wj2fApp6SjtsMG73IYd2l4+G9t2OCquWKcG6TkVGokVdXZ8hnzu0S1lZlJmo
reIhGqVBvfUsPXTXSD+ZvfvtAmE4fDyi82xhKPZwSLRCbQrwVJ7lh+3tCk+Iep/Kf2AOAxuyv3e3
kT/eBjD+iwQomrx4lEDjMtHNoxUKG96p472ZnRwvjdUdAPhkMQaazL5MPbT1MDjl/LrvCJxy22oa
GhUR/627nolmP0/V1vYvo5dh/S+7JHL+BY1Q+dzy6Llaogt00Bf39tiLGv5I1D8fxFAfziXzx/MZ
jQn7V4xieyuqIYr4wkaprkeJVnuJadtU1VUEjxjdKi/ya129zvuEJ2Madka670z2RtOIoeo4/b0A
EYZ2yhXuIjcSxmmETlDzNoSNdOn5lrQmIiEur3pog45Hrqh+6hvSbWO1MuXkHRGqV4bEDFTrVwk+
oeYMOdQ5sDtLtf1HLTDL+ANzAA+uqN7p/qCNEpZuG8irg6OBOjthsfx5yqZseVSXwoLDm4d+8i3G
ZaRzPffNmZC+1xk+eQifjgzcOEq9VC/ZOZQ6kp7EypIkIT0HfOdh9fr+kn4wSG4GDWBHeDZwMwng
1/qks0xMtv2BPgjD4bucqBGXode7gWEMslpps1PI/dX40Gqiw54CTORIMy639WsKql+PlR1XgkkF
tZgFpK52ygvsmEV65X6g22+NmEqHzJLLIgdHrTCoZiIxBF0S8sAuB4KWD5XAFhj1jx52hjS0YI/L
ysM8he/gDBpd880t5pg+M0cJhNfVdHIXR4+Q98kf4Lypw0ezCeHqY1UF2YHK1ftGb8i34lwrY18S
X+CMgQyeFWO4UNucStiS0jckA0xGuF2rBX3ZveSPZWyLlewXzEPfKkasWMlpZXx+Zl/eOd0Q0bVT
sCPrtY1LWVAqQWeUDh9elGClIR654uVPdu84wT8ctqlQ02+j6gTK+Y/zK6nDxT0jDciy5lNPnVs7
tjWE2lXqDCweA/+U1xk3b3I0n+mxs/jZn5cDsBcyPRqDbdpdnAD6CDFGRsFakaKmgwJT+r8RalPZ
r7ddL7quVdsW13Wx7JGzwBzZtYB0Iz/7rLNioAvqjaTiJ8tNwdQ1ERWNwjoZMXO02oUhOpLUKoOQ
4ArbdqIIhKXIHHRkZDohIL0HhdXPJ+kzlrgjFn2RiejBbs4WxoxZGC/CFRGp/fjLh3esc5LXDqbj
cWFfU2trfaaFpa32D8g5EexHQaC+W+RvMfRS0jaSZ+j9yTo021eJXpOtZVGhs5BZs9/5gmL7kQ4v
TkyXkpp6Z8YtSjGhyAy1x3Su0fmo0yWIJX7wcw/4gXFtRXqB3At5QsUnTzH8u1UG+VtJ3f+ABDaA
25eOQm5v7u65rJdbOnr4pC3nVzU4oWuyBT+HO4byFzHDhT0j4IONGZgdwsg2fSMK7pGbq9fn7mma
ftq/t7p1vyLue6BbN2aEsMyVLMBcyH8T2z3tWPbfnWd+jtClBO7vzJxsyv5Dbm7yFyCjN7kxC/lT
k4AcZOYFr8iG4Qhg5DHIKaHNZpTkOkXhwJs5ljxGHvdJgA27KgHnpJdhsJYrxbE6yJEk8tlIbuH3
AM7/SW2jzC0FSHjEZH87rMM3zX7dlJBCiZ9YB0LbDPQmcg56bh5U3a0Iskzj6IsfaG51f7p1bGo0
6Z9NHLusNzqb28zlcQJ5H+F5ItKpTuDmSOJETZjGhJmFGdMg0tcPi3pu9Ct4okR4Kb3By/pA2KmO
TfXngi/LqinzcwggvAr6VFarN38ZNuuTJja+AtAX22MpGeqpqyMN4AK9W1ROZLsBt+q6CfAV3XEK
J4I7vATpnLM1OQLYgEQfqWnJ3eNEPSE/XmqrNDRT4BuOO4w42ZVfLcRfSNu1251w4EJY5+RpQmJU
k1Hkm3+i3qRxp4hmCjeAtgHlPb5ou2cR+ct8O4b9z5/aBf3CCA53F1olgtuYfsYebqI/tcYcGKRt
hKypNC9548VokPk/3njQC0ZV7N5UcApBzZySKCjD6Iw8a2m4nvsj2NMOkQSE8P868U2yIZCynFNj
Fm5jWSrdQsHSHn3nCTe2/rtCLCgb0Xeef8AGaR25YDDi5aHSa6lFd/gtmcjfrXB5qotrnfPx26Oc
cP4BbLAYDuv0uYG+u7HDV96hW5Cop8KlWGRBE8i05+fYyLsrYS9OAyQzqYPI/UbRv3NyeIVRBfkS
uW0ClbTfKzq4Q47RqygoR0PJMMzBSKhKAVXyQFOFLECOjYtyYY5YRA3L/iqmJtYY+UgWqEM2h77t
4IBaujhmfeJhl/IcBxI2yJTxtxyZIl2kXcNCRzci6ylTrRLa2Fn2KjNpGhwCHvLobnRIskj2TbZh
dS2qvYIfvnArTDv5GhofByBfUhk9A2v6GxQqcFnged0kZju43kKHhzYYL9vsi7LpxQnrtSsatz1j
Lje53mmVUfByQrJlWCVYB10h1IO8P1l/f/yGTpPaf1AXsoav5CxR9KvC2I6gXbTw/E4tFQjsLtKd
zdSa9iPvYkGOHkGMRv+uF9Z5N/2Vr58Zz2FvU4UNxwC9DzmEfE70frIztk5pdWAutnv9dbSkGJZT
818xbXggnsfOCcbjXraeku1vDLti2t3SF8Xq71LWMkG38HUy9ReFe0WWWp57RrRjR1pbHMwvXUzO
IVyR0OAO3JQpA41ie/gvlShP8QHogzno7DkS6zFRRrBimlT7cyxyA1tnNveAL8bf355SdIIsZ8Mf
k560pUkcw7bk/phw/pqBonZZRQZQfWMHDlTQbkEmnYToR3uMWHSyGDcdLrBumqFLTwq3awLIR5lT
RyXq2z5XglTvnOgxJPy6BIzE0Ft/nZ6ELRsKQRGnfCLmrUm9r+4rWfCEEPApXodQuT1FgK7NSMHH
9LtRD5mbZbaGlSBDCPCPXo+8tvGcV8VmKrMiavb1eoKWRsQlBwTaAIturVP6wmOMbOQIIQUgOkub
0km+Z8Xf+fDs2Bwh8lxgenqxwj9xOfIe+XjqfIRtFkCKDlhbiKYtuegvrsZ5C+X9/nkjqg+ONsI9
ehiuhdbl9azCWcyKICcWx03VrUU8+xLs+7hmVUTvv0hF04ljdxPDRKw9z5B5sKnS69MuFrn+0601
KQ6yHF44+3bQRuyDzZMsdsm3C2moOBA0Q69i5XACCC3Ifs7ignZo3R/tSfgQq6bv4l8SZt82YhOu
oyc5c31iELCc8+he8AF8K1BrCTCGnPgTyzBeh++RGN3p/l+FOoGYN7GYXmm7uLAoTakPjRSzf/wu
Bh8T086gKLKbWmvc9hNX3cNQNYVDKojof2ZP2B1qRejZpoNrKNeQcIZgx8GP3DqQPv1GqnjD+vTw
ql6mMWsdDGislutwIhbIUTij9EWXjQVnEPglsQweZZDB9KFBuOVyY27qbegMgDTR5fLTI8Pkb64b
i4XyMZ3xpoDyyw7JF+6ttAlufOGkpb55TlcQp4Q2OxHYQbu+1Ywlp30AZI0TQdP+t48JYbOoA7eB
pheU7FsAJ9nPZTsqcneVJ5FOmCAX4h+QN6u10FeKtrRmiJPZW2y1PfVW9E5F16llWgNMPsommFgd
MASamWTzyxwNUTH+y63crQPn4r+rfFSQiJNVYSw7baEJ4gyNzndjQNcAPSnc51g05HOUNTwCrlYE
jwO2xFKD6rl5UyE3g2tifH2cb4Z0oSS9Jpx1OJcvYcfQO9L7Xu32XTD4CoREhPTtW+8IMM6thf6q
wvXkWe7LOrfBG2j3ipQmRPEY+yGGauPpCumJGi1PWP4QR519zFe4EK7bnmKKfQMAlX9jCq6QGKP7
0cdXV1+o/T4nd/8YXIoo4LZtNnur0PivfR+HMwR5JUthDz8tUBAJOFqT5azUVr1Z8lGOVcCVdFSt
R6WCfIekJyv6pow3A2BRfuDzdn6V+n5T8dDiedRFpe4E5XsJscPlauGi7/sZHSKFqAcONArVKLQb
UocMqApDl7dn3y/JPI6jV+Qxa7tnjy5tSmayLqFi4YX1ZZZi8tfK9rOmWFdOIuTyk0ErXik/zyhW
Jdi4/dOzWzoJSC+4mNwl2rdIbVp17GIbECnv9h1eD1xKfzMSaK/bL3UWvNhJI++gtXro0suHb5zO
BRhHHgR5d8bPCQWZ+R8k2Qlx3gD+2U/VonY5zhwdB+qUIimuJWZto+ScYcUB5m5sthfbV6hUas/2
zmdjXQlub2utQW4CJklKL13565qSLy+pwAR2Yi4EdYJbyWSROaOfcSW2qK9H6VDk3UBnbcX1Fj6p
DCEtEpI2LFS6Rt8KX2DTwxrupziAUrz7FJ1PveTLcJJXGoYC39jakNFijLOr8IF9FuLcW9g03czb
8ApG3z9qlWsrRum76QOauGgMzVh14HaBAHorXvdhsqR/cWFZYXNqlonxCisHumhRO+Id3tuZZYjO
IByD/WOOXe1E7N2cOreq6Rjjl511FwlMrP1XnzBSYcl30ck+oVQikiL9XEvRCSS5jk6Z0Mqb1myM
lrgXdtsg6yAhcDHXd4TFhdydBkYqCMjob1ikK3xoNAi6b5ROzZ7YZG5pUm23kTCyUjBgIkYkt1GW
R29XORiAEjAhKmMjO8SuNyRCqKkj/7gIokYLGjcsC8QDI9InjzDfBEnYO6/fpgA37nwb49Yw51Xv
zZnYRgsJ1QUeXLtuu+Ieon2a8rIeHJYaLAyZ2QH9JbyGVzrdqkfHQjbyJ6UEc7dGYBLk5MxALAGV
MMw9YZZzllfKVp6K+yRbg7S2W5N0x1688HZMjHjK2hhwj4An0+ULKYOZtUNY2314tlwRvXt8c3N1
13czJ/tsRG52KJUxYf4SVLm+mFFoua+a4mb1VKpUV7wwarauRF0JuOVk8HA/Y81+Xfhu/PYv4kpz
lZz3w995Iqiw4nGzgu4sU+bLXJIv5eXjwr8BWIInJStRoJTOx54YNsKhWsbiyuIoUdjkhWTPz9D6
RyWOjuWSNSE5RD538IiPzU+Uali6gGef1us8maIgcUI+gnR3DBS/r5852vOe/imPhkh2EdxEWNTd
IhpPc5xcU4Pt8OF8oTvJAKqHfrrww0o0BjgEtC7KXb+JIA6x/pZa8uKg/UVmYkTAEyni+Qt4/1CF
SZ7BxJt12XTQkbmM1Gn7PD/v0D4Dfxjw81tbIWKEwa6AE+x6ltE5DRT0h5PvXHz8jAwU87LM9lM0
aOBCXL4Se7R9/3OpXPjLl7xixPB2Q1AdcY/yTNLyIsXiejrfIL3Y/njQ3H3l0yapEqCCgFAHZOOs
NS+266mKgZ2yxGbdw0dh+bBSqNRax9MoGfdbvP3iae9nNU+vP0VVU7xbKD+AGptJWKQblhNGcMO1
EeEFRydscuSuqrDjUZw+aeLugRRriGBFS7o2FtH5zi8UziefZ1LbOFhEG4Blma7d2PFRRPvpoTlb
YAj/vMWEfmz2RDhYDmL0cvaE8aJ+Ya5tyLS7awLovZ7ENsl+hQMp0/KaNs15UD2Nudmzr/eOt+MZ
xFgOcT1qE1JKxM0X9xVvLJ2eHGHaB3A3i0w8/kAv2FIeZ8PFfQMkKSutv36voYItNkjX91eAHubM
cCJ/ELfWT9n3CSGBlt14M5Hqqn/CkkZGsyHjU5kIMzkKfk4sjnQEr7tkDA4CgMcjVbp78btTt1wL
NyENA3P8wO7+vqES5Yui0u/RvfLmW2tATi1qvskfTQMHlJE4xz1aKCPefp9IxwRj39PZXwV9qupj
pmftv6j1RTKqOJA/IonpvJ6R/USyfXhOg/GDRKOtAZbQlgGizlMW5fCS8B0KWfXZ0yMKAO/cuXbH
74k5rcMFsUdEMRqgUVOghDDgnG98Zy1QAMQbmOrwQjG1gk+8mn/WEKswPCzKflqdGJrRECvH11GH
OGkD6x3RXsSf61P/9Im7DFSDUVDD+sAQ6Xz53D+iQe15hgodh0d+mpL1pqVN45KaelwjT06xEc1g
EqwyT+42xaMYUINeogJD6etGvT526sZbZndAuMofs0h8M1vvhDj6SjycXvKrufUCMRIJK3QmIiGP
Xe4B4kgqUH41SXiUscQvxmFdX9H9Q4wmgBITJcmNhZCmW33R+dMyrMClU6fvLajljTqqznWy4l5N
gIM+3aGlR0qbB1ng0q2ccbhMMVRxWE0guN0ervWNDuR1dDVypcoTNHRQ53cVukToNtqNPcyiZ4O1
ZGs4cvFJvzs+e4KV5/40vM6OhRhOZRR15QmyDn4s5Xr9tv896Z81bMzQJPh/b7mgx2GxlJX2SFYU
hxJSdmO9OZFdL+y2cYBfQ6yQ6LyJvisBu/qC6oKL7Qe25NLnjOKa7S024DvdjyFggbA3GwYYUN6K
MmmD8cNTbNAKhmCqp96eu99UyKaIOF0I2ZBUH+UyIQf4GcoKAJbnYjhW5+tbACQXOcjBuoiuQXEx
JPBlEpeBOm83HlwFA1QrIuR0TBorb99iplCC8entOthHqeTjotAH3ZP4eyDXtbjgp/F8Rx3JWe3P
hgCz05jmvVsfoD3IVL+BovkffHGBOwC8iOLRBoYRGiS/zCxbcJ6BKVtTC5uo2/945xdNTE2mIsCw
OGgq6gUtHkB/KTfAWoBVUbKJ+lfPJlnij/hNlaHu2KGe6J/OeYp/tne0BY08WIgcjtqDSiWquwWA
7QO22+/8XTudIeSY2HePeYEBvpIv83p1/tY6eDL3V5NG4X4c49yhpmSWlp4TW+OPgdBJ9ZRZU6Zc
ULrDoHg19BxHO4QSGfCoTAkQ9oR6UnklWy4nhNTLNAQDJwH/mylnU9bvwIPwUJZ8/QnsusV/aqPS
c4+Fcj+3gI73AANop1KBfadA7OFwPZ/nO4Q3UQkszfriieY+E2X10hl3NOSXDWUNi2Hhc8hGfVa7
eAgNZcFii/TwBA2KU/TNP8lIXOugOXKn5SaMj55u3SrHsNaCLZ4k/wFjN7HQhr3JOByeH+DNux77
lcO5W8zJ9nzpiTrh+DIwGt47i4iodyOhoCNiVtY9NakGv3TLcURNDZ0fgNAQgze2TDAGDXbk0ZdW
McKy+P5OdFrARzI0A5a/chTWyg3hmloTu8z4+jVnf5ridJ1GpebN/pUlOo67fkSsONXZ3w7o9/0A
VT75WY9X4GecBHd2o9SCf2JhgFfcPGplnspMSUWj15kB9hKP1DOl4lYxte+I/LibWfTchJ1bOwPr
ub/C+gxWGaG7gjdYPkSX10nJlk09Hn8s1mWykXeWf4Y9rFNAotJI3rKzRce62/6C3HPwdAVeRkey
k8OXdWHrqIhKE0M8864UaYm3KCij5e2eWfSJGW7kuiWJnYuYpGHQEqeSDcr5CSOb+sg/IClqvNxT
BIJejDfRd0R/v+CYFpGWKSqL9imlP+03tO7P/Rezdwo59k5OBevLIXmdOoqrfskSl/qRcYw0cqJL
6zKB9T2AAs/bfhAGzsy73RhIXhrk+z/AwcCudeFGCUQ2OZB6hGi6SNujTjgdgmorDsGjN6sjb8Bq
oXy61OyHvPCKjm2B8/wHJEzujF6sugh/ONd+y8q3TIFO6G2WtIbh24uHGYfHeKSszhaTsxOkNaP9
DlviKotkE7gQeAoruXBlwNkTVznyVrTzju3u7Zmg71iX1itY59xedsQxveGkYVf4qPN4zZCiwznz
Tn7cJWsDM72UQCfMjbv6Z4NduOk+sAm94R7uVTdbqm62Q/BlyLGtAHFsI5GYUZq3x2lFcWtaF3zA
eklXvbhRV8h527+/LViBKR5HS5QKyX6uX2+4Swyf3c5jTuY2gK19prmMQdu8F9ycueK2ML57fIF7
AhZdp5D4QB5/WGWjd4cf+SQqzzB2tmhyHbwm35rvA6dtCwGgP0x9DNoZP7DOW3SN1vsa33OulD9N
YN59w6sV7Dbx6Zlgn5f4IDiHkt5FJbhHHqJ5O4Og1EZpo2BA830qnfxTHLe4JpmEiMKydLjjjl5E
L833QR4OAgw1zKVwL8hep9t7fVlMSH4cvgUap68rL4Zp1HwcXEGcduswG2G8e63V7J+ZRuLy4cwd
0IaF6Gz1INx+h8oCWSLFgZLi077V94T4jJbcgPLFDMfOcaeczfGLvflFUJpmNFuaGsqSg12aLSVs
b8dIuXWAgOptpupQU7/VZhEPKQM7JTLfgqHJv9SPIBsVH6YttiXX8FCYw/XCihFhQIMJaDDIL/dm
8ChEdSNLLZr3YPluwOSQurgejfYW0EpY/RkJo98trW3LbxpnXhtiXPj2tWRJhjc+RuNoHDjx1riS
ZjDoMyY2kPE51lm0b7TIJGx1ufmf6cFpCp6KSuZ/IqxkPlffnUt1QyVrUSMLsYNi9s/Q7Y81Xsy/
hEzJ83QdqZyzlmtXhsKW35tRGalvzYr1gdgKJ7sCKD60EMMplNCfXs643BKBevjvfBdFDoMJG9xU
Uf8dT9If/trXKCS2iTXHLJVbyDf33fvN3PITvcBKszPdbc2ZWNuKWlLHj1bGLlwXUf8jhZoPl7Tv
DQknQE+Eec+epozbFq7Yh8nPISTEe7PA4CejlAA4a4vN7dUW37Ntxr0iJPCFBZ/hIjDxbejFOXOY
Ls5wNROQo/JvetnRrO3VWRgI99/WDYPuLiJZOPxr70T/42AslOxo8mL7J3O4mBLWX/xXo4xdgnrz
Y7ir9MvuFhxD9zas99X+HEJid7LvxlNdv7PsFBuOzTkZA92hJSRKV8Ai3hqHER/pggvzlN+oDCDo
//fadMooDeAw25nsQcP7fZlKwPpvjRx4sPvG5k/DtxcxGsT6P6odVhbTcIfBFK1oREx8EExu0ami
dWkqsVjTjno7C9xuQ41rkYQkTu/fgJpwdLMjuN0NV82MynbW1eLrf1sA+6R+SoAK33K2jxZSdV0M
IvWVrGfe3c59GbZ/hPbQyZEveyIrA36mk2X80GIwg/SJuoMnop4om0qWSLPmtGMDskwoDOTiSgNs
Q5YHln3BdpiP7HFQExWX1QcrMahSpHiFTOF/QRVdYojHlZt+gWguNDKVskP7OvRL+RLmBAaHryMQ
0z3AZu8hvtqHCQ/Ziwyl0Ow4nqyr1XV1T5qvK42/kPm3/Vie/0yO54WFXNKTDtZ5CBvOKvQXrSyI
wdeXHNABFmnWc2WfYZk/F0AcRzfiiig/2BqhBK+VEx3jAB/TCAO34RWR9c8w4XyIxR1TKE3iHd6G
XZPgwvnjJhMotgAVOWvmrywF8uMPgDGsf61d1RxFnCk5SXKDhztlr/tDhZBXWhK2hmZxvjXndvds
0+Qy19lu4MCQHF14KQvtma6oKgcmy6ejI1KzuZpyuDmZqkicwRL/V6NgZIF3xWajFaU5pkwStsJN
FS4Q0QrOev2xE+5nIoM67eHgNAeKYnPmsg9VkU5QNqdeIxBTgI2/ERVMGyL+SngL9iHrjffKAOWT
K5LgMaQJKOeXnUcZ+vjshx/H+fvJNYQcqYOZ58KdrS88WZ9hMyu8HxLKMUIR8c/iPyv8H/OXrOFp
thx+9YNMkLgQQjcaFvU+3HNSZi9Bu5DrsJdroIkGD0u0AI22caslIxAnwqr/ym+kklBIoXnBENfJ
xZqeq4J5QaaWrqcqPMOfIFfHHAzjIKAAE48xU6TgQTCZ4Tv5Cpqd6bZKGTyQama27vGYXSejjHVH
W6lnrSi2jFYPb1kbcv0K1NgtngS6xcpjpB9tf0nplRHC8RsT3D8V7w9mzXBNHvY+5uJ8MLxxeQgq
x2+ZktfaHU882kI9FaSLYM9ifdUbDr+eA3UYANh7E4wMuCWxQBWIt9rGy7NVF3kTuo4Gw8+LJ/Nq
HbZd17zEeOPlvFUiHtSHx7PyIa/SEHdhVSBjQYKWIBf7nl9W658X7TPWxr0uMe63yS1QWLZqfPZj
nR8lXFgC+6tV0cv7idEK92bn4Ox272oYo3dBsGzxmECABOo4ScMPpBvqMAvePURWS1/dgOFwTd6k
LqP44ibefoZ9idgpUCgGfxUlaV4dH3TnK5gLATADbBY8gf1iWiDs4pzF6ar3fXe1Izx1zweohdKI
271vWhOpBOTvRpwuhARs9fkSBCr0Wo9Cici0SeavHNfMjvfTXpqLhDFZSg+GnNCh/vikouZuuqwb
aQhLm437uQdJGnBFrbUOvzU4iWf9iLUYZhk6wO098qp1xvP23aRTSvT+rBgsyfYzs4sMzwlfBMvJ
jB/T86Om81lVmT6e1OBz/UZHNXKUWXSR3YCEWhounqzqP2mMVy2KsUZbvcYEGYMlDpO8Pfny2/m0
JabR1aRGlIYWBYlUqsAljSYgg6TPRu6ITkGfEo5iXrV9jMqKh6J2lh9DIh6pRaxKRkLQU945frdo
/tKgEyIrkxrmwHmqzMFs+RPF/cnKtIFpNUpN0N3O4jDhIlX7LSg7v3XdMyMiONBrD78QhtyKbRXo
0yZEoMkzThxvk6XkI2CyHoOmUQaZZxG0eEKX2raFu78bF7EhOcO64vmm4bHUomXa50SOrfzK0EOm
l1xCBc2wVODsLSFLJ5bfYEF/iwwypDER1OQQTcQnNGOnDYaX5YEis34fTHgpLhCGXftO9Y+8hErY
Fotf8Ve7pNZ5BPwOOip/AuHE1GdpfkDrNga23p9ezeY2iak4Uzh483rE3jHfYhCoDyMudOAm5YLj
GViURXymkZ5CSAP/G4U+smytbap9xbkn4TsIQZPQeRfoHbxxBJQNC9wEtPUHAjLRk/GAtV0g1ke6
VZ9nWzsiyzkgSJbTWittXIn4UL11T7PIY+TPbMOC/s8HLMJ7SBks3WpwPNJ8MBs74Z9p86pcEAJs
plxCLzdQnLJxxMBb3tKZBfHFLaFSe6QnWQu2lqfrm3ZR/8kfhAmRhmcZ9VHYo0kDtLBQHSsTxASI
GUo8EAUq6CpNVc9z9va/Gd19DYnu7hrh4nqwLql4XZJqiNPLsp9Ow0Y+kaH2d5ysqmGLDpkOb7nT
queQBDIRPF8l5MLZR7yssfg7gsAcM5rx+mIiNyNAr/FxGC+X3Twv086BCwaGJaFXhuij25rRqSZf
amD0iDK9xPZijD4oLyj8a+1+Ih0cji4GW8vx0loLnsxXzmK2ETHmotxxDJAqhSDETiQgArEt+FH3
FhWFMJtu2uOipJQT5YDqAz4bg0oTr8h97+feKE2l6CBAf3j/PKEfnsRUyWNEyPt2Hul4UgxSWwMH
HaLCrrNVdI7YxsPxxfHYhlwpH9wlXFg2E2+A0gMF//q1UWymzKPx4f99I2j/VAYX3ZjQjl6KzkAP
h1HDS0vy1AH0+gQpoohSoz0PEsUIFEedpa51glEHW+SmOd7YaQ4gYRMfAopa9Ml64UMjTwst4Hne
x3e6+utjwaRWmzxAWRYXvHPT5+R6uCE4DoOq1Z2yeGMA39iwvVa6cVQIo9Ih4RnBqpDjATeseCjR
838kTI1eit5TWiuZ1kPo5ez6KJbVVYxXep7F6hOsTwIM2/qVlNo7OTtjQ46/ESYJJSCX8WDrGBEI
/i2T4Xi9Uk3QMzl8hylkJrpdIaYyZYoTyU1ZphbST1+raQmJeduvqrLJsVXrIO15emi5nXlf7G5s
2e80DS+b/7bA4X7BKZPyYctBhIhgslG04/4Fb92Wd4BwQBwvPyPhaFZt9YDsO6AwAG17B+zbQnsl
olMSLxhRFmv4ahVEPK3lL4JxN9VOuq7PvcEFZA2DCX74qWKifOU0vF5CSpfTm1mCa7ye5Zx/xkPO
FujENHZ4Ou39kFB53bd9+8YNlG7UnR94wgnKt5EkC2TDKDS9LKST4UEXKo5wqFYn9AESU/JfbEAU
qTB767PF2CkNy51tug01OT+oeKqaJOMDJFHkUVn/fLNGansgCQdY64o6Zn/qPETLbTfcNBJOLNwa
s0LufrHp900qbCUEcZtquDaSgexrmWoNhNij4cZZC3k5ht6PcmB2f5iFxDwmUPlto3Tn8ywXrunw
1d/S7lesyD/IyTRZw7J+XUjEsgGkuyo/KAPocZP3IIfcYkOuHg+16UkC1ymCstbsyCGiuhX6Rdm8
rS/iW+bBeLcC65SL34bHOOBxBVspM9WV1uUOSnIjhGhHBT5CrlfaYjOTloE7RYaoa+79xl3X6gyR
ytP4bg+kwN/VBJXX/DzpTrmZKMAyqH4TRcJ/Yk3me13lUAqPXtaGwAnOm87IizZ45nbFlFmfuIXK
yvDx76qInRm7d5t4mwz+Zi6FCmZOKYJ6TPYof7jidQrgk9/49rwvXu7cuSarmOWk9ENe1ZJ7IGIp
0oRGb02QW4dWzfDrPkjCXiELb5yxP1yVIdOMOav9xm58HqtziK/Ie/ouA6mZkgxou20FSyG9acUl
nJp8oEy2wdRvFrGkumWMNIbCwbSb5s2wTgtNjgq2JmmnMrAQp86bSn4tsQcLLtxVbE7rpPqethCo
/GAFEVTbPsgI4WN6oU8gNflIL8s3SI18aLOVRVDMwMqkve+X0LoxEIHoj0P5/xEaSBbUApLoVPAo
b688ghfQjjZzyX9F1zHtNscf25U+p2SU8VTll2N4xOAVdBzZoL2Qy9gMxaOUThC8bt3JDxZ8X6BT
01FMtKfFmKvzEnlkU99URiA5qxIf79L0vHVZQRHPpKpLmHbPhAQ78ROcV86sTHAuVVuTIoEnIoaW
Q4bv7DYEEUxU5Yb+7QGgIuqSoFyTqL/yKWK+hT1edl3jb2/yxNBiWrcmZSZWelw+x8CUO70IP9YF
EtUbGsZ2KJQo9idupWc1ww8DseiFCWuGp76PoB5nENJ1Z+H5VSW0EJRXlF6Vi/ItGpI/FZDc//t5
D2xudnsUrtwLFT5EgtpTwuAztzwVfZCOKBazNFCangewPSf6oQP1HeqhbITTxbLySc9gCoNRyxGf
JyO4QSHmmmIoHatlM7klN071IzZzr1m5E9lG6V8pZ7L58/rhqFYYAI6vx10Q9mvfGzfUuwVu74MY
AMDfCVavMkS77hEY1sJJO9hOVSx4W5JUa4Jhg7v614rB3Q9HKRYTsG2achnPF5CpEF33DakMjeEx
Forp8zb9slwAoSeaIxg7Zg3p2PxmArOjO3QLkwon5EOc3+OOahWlqgAdTHypyeiopb4MqQJhUteL
fZLzVb3NKYQQJg4CcsynKusXRZ27s3nvDh72qxr0MJMhHgnqHxNlOwCxUGw3bc8Xk1jSiMVD1sZT
Lr2qwRrtHTnPU11AQ49mJDA0I3ge6dAFr5c69Ch66Hvsa2zIrwE6/0R1wxivvJRE51YmPBWS2Jig
cPy3asnE2zxLUF+PKSEY4XmvyxMwt2IrV6ep8ozzHpTe1MrPLo8rRD6PpEmkdcOZATw7kMubnaFQ
seXc0u0rBeOhFiflezqwCuMwZkyel+EZ1Zy4zKBTaGI7BdvoQ++21qKMXAgqfWTda4c02T9AdNdW
BYki7V8A1aKcC4ysmoGMmonkA0TuVeTKapmQ2elnyrWDia3pY6iW5aBQS0pGeU4HtngnLIWxJyBe
9/94vu+nh39QdNZsIhYS01mZRn3sdCLqYslFWLYRwz10HHwmPA24K87ubBmJuLePWkH5Z/a/U8Eg
U1PlFVie7+ZxkUJKQS/UchOo/iCFE65dt7rxDdhbi0uejCJZnrQkRLdoyadvuTMqghYee7wMKuqY
CPz10gtrs/1WMBYfUjfkqsXem7BBAV7AHlVAmdB+AzXXPdIlwyrqE8IpG0IL2rotFVPzcBfqSJeO
Nxy+v3rj3yoRIHB6SaqUlSRlTGJRSiYgZMlnNEk84m6nAVWfXz3IxeTlGmeFwg3N/h8g7CZF+4zI
betEZZuADwvCnu3BjKS8/J5yEHM0APMt3/sk2X/3yKLdTpVrHvhrMMBybFuU/oAaOZYf3NjSIFCm
phsOjmalEC0tYBc4YBW1frGD35pTGnZOgpCiD8mjC4id8JLHOCPzCGOzqBuLLQz3hAfHXuuJnn8i
1BhGfOgZxSqPK0OJ5gasC2N4Q3vAyPz+w4n4yy0hFP6WZ2Y8CnwYSJ3ps8YV3xUOo7faXKJ6Idth
tWVUFN9EUzkKx8hHCjH8LkuvYUXrClBBhnYs8YY4yhI0OKllBGiQshR+R2QMVyNeSlEd/CfXWJOV
BhL+frILgs0V+mpyFLQYDCp6TiZy+gCfmzOoCavQxazOMKYxucGC7Jq38QyTLKb0P4FQc73bbxE8
jM4pBxys5gxP0MOV8AjJU+65ndIJPQJOTATNcSDwzrH6PlT8dFK8OvIbn5EUIEBeq2kIr79/y9VW
/geOgraOewHoYnMOoXnGhxtc03ZJe8FIZVbVSnyCwy9ArI7D/PsJ7bo5JYTA2ShSbjKTYqPEHB2n
WQbg/KgrguEc2l9ZjcQmQWzsY1u47QlYPwkLsEtxsTuNXZq19Fa4GqWkBDed41Riqeta6g7Flrgd
NjSnouXzOlMjkFdTsMgRC7G7Anlw2i15Ias3dFIrx9vTq1MMrhZJRYVmN1q0DcInVhzvrW4xICjW
zJbur9HQa+plp47kOLov/UFeIg9EFIAuEu245pczsO7GeGx/3O1i70bkY9WaKHMQC42smSO6YyLb
Pa+EgthXjh7agU9AmnGjqeJlWptiNfwOmBYCv5J3LcR5IrWVnbdWB2rul406YTGaUJHXQa1xoZJW
QHm72K8eyLw/o4ojh6SzVTWouAcJWoqpMAnKzVHGuUADNB7IUYNcImpDKNogislEyCyh4RNuh8gl
QFj8OJQRPqGfwsZ96L/c5X2WcHizXfFDyRFjhbxBemU4haFQtr6etEgax+MvAewGMJy48Du8LY7z
ivD0e2iD4c/89zUFvwmFnZdacGry8muPOYq9dlKMfHGM8mvxUSxFakxh7Wc09xfKkyiCmYmerEJJ
Pb7C+0A+NCcbRWtnF8OXT4vMihJyMcKOahLkhCew8G7G/RglHid4Npq8Q9dn8QAvlkjau3Pdi8vB
tpBlSIgCg3ilJ0EvBQezH1aKuLcQTQt4f3/4ifGsiv0W/7xVDTl+3Cfei+U15lrGq82RZHRLVm+3
pnepvHQ1S2KBkHqgwb/cBiYWgsIacR1VFOPbOH2V+Qo0K4SHmkMs+K/zfEIFT8RvuaCXT7KNJtJc
XzJkpkd9L6w+t5ZcfxVaz10T/PJ4x8ptSkZrc8uuMJGC/adfbJqfWfP0IYj50JSRsH6vsF0UXxVU
uU8+brDzTlwBrjJfiQK3EOweQJYyDL2HHPdEivu3UAcYfRONY92frLOeXWQiloTJzIBSKZ7vSzWK
fiYa1dw8l5LO6dmLbD7qzeWi9XZ/af2l4uB1UHXCj4aBqZmqLbSVr+HamtuUZZuair6g4LB4rTzC
pkE9HwpZilbdnRLyki7f+7IDlvN7PsjxGYQ4BptFVuKQj67cP6lXV9f0iZqofKics3igYXX+ecVi
Ql/k9nmVV/h5uPItqP58Gs84yCUaUsUlUKeIMtktKgaDojMkAbztmR8lR59Oq8UlGkZSm5+1pTE5
CDKrWuith70My1eorIn8HmmPnwv4wI67j/qqlB1ro2/RJVwp725aNntYtFdmj3MTQUPjMF8GueCB
XU6CSQiecYLK3YXwJY53BSFFihCs1IkjIOtLCSmOshSZDWGNd9T1iQiJFQu4OG7qp+nB0S5nJaB+
7LVdBGnj8q2ZKckfEMEW3MH1U4VP+D5oDd88MBUk46sufilZHSsjINu+WxsyEV32+Ue7uoDVzGbN
fX5PKEccss2RKpdrVKIpimDV0HY8UqxrYEXeK5HbRYBxxqGHXbqCYCcux4GVXrYnK5rnHyxRnOG8
/mZMC29kWget7nyGuixJuV5Qgo9rmdvm/RHrjlPAa4b4NHVBDZD733gFQJouov+1cmqGq9Lu8nN+
o8wP5+bJsPwiBYWsa4tKP/IgsC7XbWT4uEATR9Fwonl2rbiZgQoA2/jxL9dRtU4P1gD2MDKbL76t
PUZqsTHqM+sXq+oJEn6y4B0kCKq+9x/5OKhHaOagCPb1gTCMLIAOxHfw1fPJL4ZwLxwhTyko9O6K
BK2U6SnH/HGxAWVfvULkmKprKGmDtBqPgKPV/Veaw4p1Gp1Ivl3uffGhbDLYAqaKAkHI7pkauNpn
1tXCH0GmjxuTZMvzLhXo2VWNQ5MR4VW2/mF2pd5JB7xh6LpeGhbq0konKeWgIuXnM6bomyLWLRib
sRgZU755XfJwHIwCbHbdSQKCXTzWi04JthXXRjIRyNlAjVDSuN4KB+vzAxEd7hLRhlervJvGtd4i
J9GAHbr2dP3W69N22XaLJXKDU7x7XVdtCGbKwkfdyTakildveJdxFLVv51HHAfy7gzeP+4EQkFX1
7JT/4P0abMMxEOyNH8gy9twOo+PU7eBwe1KYOWyQH92cFYXPVYnNdgmf0A9HgHjcmed5kjbEQUsB
gD04GkBHq6XZHnXYKDKXJA9sj8P5CDJFQHI4+xJD4NbdPprBm2dRLnKjNSRv2aYq8TbeC5LSdu6B
ACQCr/WyuEyPHyIj7bGuFbKePHiC6LHroftN8DCn622VS/tUR8aJfjFvBvM4/Z64WZOPcJuFBQ3C
onZB41pjVj9EUXdziZ8RGaFeg9+vG0Za/TbepLHsGhrDL+BsgZ/CwHEhUj4sb0WmUbEwPU0a56v9
yOcD+XnOibiiQxGgIld8MLG+Ft/CgIXivhhn8tXuQADt+YQEieGsHmHHu5MuOhLcT3Qb0njUh/OB
+LKJriH1RGrMRuSdLP8X4JEui5hA6Cn9cxdyvUUjy1DciR6AiawgjVkOWWpgs0njFHuFfdifeiEk
dWjt6O5OfJ1XTRlVDUWQa4VKz4AkTNIy3/D6K+b5Tn8YnvgA4PXgrl/Tdr7dRiYN1L3584kcuNnr
4/bJvJv9rF3PsAjOdHtDgzxlloTbE2QK7iz5H2OoTIkfD/AbOaqyE1TGRSMb0OQXZIdtqwy5aO2B
EMC/1HW0y6FMtVad/0jo6mN2Tn7xgleSiLT+F1x4BSWM2/noKEwfklBom/y3lBgS2NufL6UG8X8Q
BPaSd4ey2ot/oi4lEatsq24CnPL3yTMDTwFF4OgMqFB0odPOLehs0Tqz/oH/KHB5anonnYBdMNYc
1zinLeB4mIpsfz/8VnX2g/JfJi15M0vPX4umOOWqLTuEv3ne5DY6uMGN0n8+HKY8i2P3paHRpBrD
18IE7z3Rz0f/5ND8ND8mMOgDSenTOS0YLk3YIWP+W5R26yuad6KSrL7X/ig9EQ94hyJTzSqbVXg5
I0Q/ZM1kSsfNOpYeQML7gUCjoCWKJ7klnohNT5p3Ld7Z6o5mEc1VbjPTyDNeiZ2MUNleuu+uWLNj
9v5K3Yh1jc+OaKdbL3wof7oq8R2hzAvf/BXgNecF7JyIb0P+uKvldys9wHspkwdUNvnODwc1wv1J
JR4+PuR90ky0VW80JzmFjP6Xw+SAXBBAVcqw/6pmP10FABG9Lg//ADEmKS1OzDxbI9r7NzIw8OLl
axR5a0DJiQ1krxtGmWPShto0QHCunAUhflPJqfTgysyLatviZcjzaeBK4o+IqsQoLBNUzpNaI7DJ
5f7S5jhZaKxoW7XlH2HfWvQlM258ajai6looT1KSl3P9jadDfi7StYG7Qw2RuUaeP+B1rWlWIWDw
NMtGm5OApk7jDgPNfP0Rx3hUzbPfuNSqiR97YqvTkhl8IQ7exCttiBHL3BnRssWrxVz8P/vQwBun
rmjm7rgBPyoUFYj/wozTdMzQgnhRWl2f4kqcqfPhQVRPAkAcL7Fmms9DCXgCP+nCGyEaowx0jzX3
UgyFBEsU6GR+dW/Wfn9suR7FXrOUlyEMII9qaPy+1RmZnF1JxRrXzmy23REFUBvnrgr1Ftnn1pTi
bVGL+g5nFFq5Fes6s4OAGYKGIfeqjNrLlWBxJOAiYVgH87r58o0Zv9QdYbmV/w++tAwlBGkMMhIT
KQ1gOCZcQgGxm6uFYdk4uMnAUrmrpH+RsTUTnDeFWLDuVeyW0rb6kUOeL92IYf/1Ow7svRhoch0H
10J8lcMNxeUlFH6Q4ZQifvET93qn53l0T9e1Bt62qBBIrMJfQHLzh9s9zuR9lPdn9n6RDGXaOctD
JxBdwLpTowj0pR9EhpTeiJrZ7HPwMKNoWSWm6C42dq53s3LOwFxP0iqTxf1rlR5YuU9+OHAKHdGY
yFxm+q7W3kqpEAvEbuvvGhOa4qdsdT6iP9MVqY16oBgrv2eNXdyDHlkEnUoizwKmpFUQfu8sR/+l
kHzYekQIodMF+nhkxIrAazvgTDLfFVhCo2a5rnKMc9B0awQ+D0+S09HW2QgKb+HkocUVmFjMCKi4
/kgua3irxkx9CM2/jcvNrkp8XwSH779h+SGQQfoZLOtbr/ywNZFZaFlKK8qejXqv0tfIvCoLNfVH
DDhqWpVmWe2SZUmeyqMUmXGFhEJbcVSDUfT/P0bWbVOqoeDZzRdjmADvrCntguLhaZK2u+syDBD8
sTPJK/30JZpbHGRxTwLabHQZfL2sgcc5XIdbjXaxQaASipe3kek1E8BK/LSFuiMZrH2bfpOJyGRM
03+y77LvGuWl3pxzmauRU3MqDeKrrsp/TyBEQ105ESud5tLiX7ff3D1aUQksr5uvfayJpYV+qy9n
4SFYQElbNvLmV6gZoZYWNf2zBDL6pA9dRqbpMVr1taLGT9bjmQN1bOp2Eo5aydxDKhtNZoZOue9R
tkMJIj9vWo8bV4PHzx7xMFgeY/vvvyuok8I75jVdEt9x8xeGLHa1CnuyngR+IaFlHdjTMtr2NPRZ
2E+S14I+eOllpnVZU5NDs4RIpQxX6HTp4Zk6yQRafewWj+UoDbBMTfoZfnflt52vezoWNxILrv+F
6j4z4SV9hhaQPiFZUgvk91TMHn0igluFbTuyawYZEPdYYoU3qUqkoT98aku40p8v3NTFnxJOihug
IcHsCmVO7nbnvZ69Ono2wLrV5bzBJO/6S7/5XYStT9j4jCdLIFLVy6lFFsp7heQGXocaowEJ7nEO
37Y+SmxH8mkknF6ZUEtO6aIQiFj3ttKmeB418BAaWZgRPLCRokRTp/wwCU4rg/o4kRkbbx6v4IlQ
BC/dw9E9D1ylWWS5ryvoSVC2nm/cTetVPRCr2Dm3Hp6lKdaeHylVimhBJgtgixFhz8c83CexoNqn
b59SmpjGrTWNHbouiJSHpCL/uGntPtwDUmWMXsy2nhkVJoDXXEnR9NkkVP2JIk53DLOG0P+1Norz
3POoqGDLep2g2BCLjksNISfxRFzRnVjKSdICA+E8rWNgjaWmHkD8kyHHSCNtVCFhTxEAM/5ibeE+
a4AaRo/XYTgYfw7Pg9riUmqNvxaMIu7BUTuG+G3BIJuXro1SxyJYC3JFyoTWg5QNbm8deoc11aBw
I579QerQpr5fWx/8qJaBE8Gnm0AwqmLF8BauMSRNselcY3BEhIKkYwQ/wzkcntMlV9dqdFqkfL0i
nwg4MfXPPmh1015Hk7FdrAH/IuA+G0fl1cCoJfr+X8ttljewfGlMv5kFXD3tyP8ER5lI6gxR5wlB
p9ipEVMhqVHyWaLWJw7Ie3oTI1krQYF586AquFb5wz/6cDJF5s/5sCghTW5ShqPB6PK35w4pwk8f
rRaOEPDrFTRuQE2mVm+Y6KMWyleimwFHfWhCGRlu5BeJptrv8Y0ekkbv174OZHdR9fuBTtVlIRYL
cHjgRK/F5fvPodGcL8v4htprgVlyoZvi1WB84Nu26ACtxUL9KZMMH9geJDyVH1VTGjm3N0oB68xS
qE+xhVfkBOE+ZOS0lX7r8varHUYBAiSSq3YQMakha/8gG6dmxlWZJsJwnmgu99NbsPWFnuxY8UXJ
BIs4wh3JzSyJcLeBGnrYDsVwcCCRYupm6+MKBtrhRFNCRPR6d1xQhlr87itlv12drNoEtU5lzkl0
y0RwOVJTNPt3c5YoMjmOUHRp2GUcgqnErYy00gIi6Pko7e5CwBVZ+gN0zk0FO9xQzX+x9EHBPsWo
7L3Rspo0h4bxI/ECO5yjuKEJEHBNZ5OCTYtD9Ff+oJGZArQ/LLy+dpco3RIhtJiCnUGd6cgnF4Pw
cYaO+hrqHG+v215y6MRODe0VQR2n+Xl1LygwYZhLbMrpFtPCf4wsqx5y/2KjOfSPPQC2XmWpGXUh
TToMSWL73QVDnv3wRNXMBzK6pKGy0Sv/lQnXBEmxz/AKcPJeLAzY69425nFIxgxU+xKWs7Bc9m2X
2EGQWCz2putnL4fAY9uj//afTKgEmNWIof1E2S+cFBbg9rc98vyKPwN8QQjm85e5994OH/3yabs0
tFByPyxvWo0OQHDnBav/NKc0cSnJ8SYtyhVcvHru+k4mxCq8KLxGpCXWqrejrAooFUCYXwUTWlCr
nC0hPBCHzbKF3GqO4d8lpm9ZdNGnH7kzRPMQUAljrjKntXZ5zERiku32AGndtheutKJQwwlbrThA
x4upnjYajumiWnYaVMFAYEm//3LIV+2dBUe/aJ+VjpjYc2i4oGUPMCRKoHDXcVytivah3rh7gzyJ
ZL9aWOYtCmKl6sTPnxrqmpdGvd+oNtco7z/WMtrxNG73UhxDss42wxr1wM6mnRNMPys6NHzuaAh4
3+WyincOUKf7o8NJwI958CdHxNVe1ohAfIKSCP2w/W4bYoCxaGdkh2KcUQ0b3NfLqPkwxz++fuTV
l+u1p2W5Xk63F5RWz9XUlHq6kuUMCyXLQiTYTzkCOt5Hi7QBTPY1d4QJIWKKGglHLeNdJmrrgQ/5
sNK2WJlqdJZO0kKWfwNeiRpYYNFnXtoJrGRuqtBshZWADeIXNmeyhCgzdh6Qi1r2cXPQuY+1ZjeH
O7qyYO/lOnaXd1/zkJpAZhLt2j17ewRbx9tDKT/MRjSeDDZ/c9hJl4PXk4u92xft5kZvgIISKTl7
9e4W522BZSl/w9no4Kz5Hm35iDpH0VFKi+HqOFK0I2VW+4Qaq+httMbF5VXgEFOp9ikuoEYrNPHr
2rxuXAak3nJj17htn2a5I7P5DbNzHvdq0Zd8FeuMxvUphsBNzpjQYXyJCqIjYrHEvZNSbP6SVcjY
693CNmrxAu+VDpKm/7gu/nRywKuYdkee8SQLeaT/waYNQEEkkCDRyHfZhc2ob8a3zJTULG9dHHIO
cohiabk04RLmgFi5JL/PEfrMFO+aSCvh5DAI4ls1xX4os/U6uWSLp7a2YPGFC01K5P6MHErv/7V9
6ZgjhYveX5BQxCwM886VDoLqyS7zvXu8l9BkC7G9sHcJvUpwn604/7fskBnxqoifUFN4N6e2GcQb
Qm2kw1SHLP81ESQr1mOFC3RI5fnpFTANYmmaNZ97QM5D6mYMjah2FnClTsHUFKx+iJV8Z9F657ly
brlTSgr0IAt0ZCImQx8S9lPLUuYhov4dxx0eI0wQdezuaFsfnjDbvIvhR6BjlV7tVbFmzuB9q/qS
8lY2t0/tcYkQ6uRY8JmIQqh76gqwThmIVPrdQMKg1IP50Yh+AaQl0/+12WaRT8vBbmOJW6r8cRNr
mHATyg5uvadJxEK8tNlo/pG3REz3MA50rew4gsBQdUoycO8gOuT/geUrzwRw6A54MQf8zabcz654
DN5M8mVOKm7emlURLGF51KUU8ZYV/HUO3a1Ynmd8kBkF6DOxvynzwZbNP55atVDxrbDEmA6Xob78
Q+f/NpLBsAwic3SXL6viM/WnBxLgWspaOiV+uUJ2VEm14FPg/1Znks79ITGYFZV/7BiuVDJli9C+
xbXLWf+/AEbAMPi95dCWODmwwqgy2LXAoe5noXQKDCnStjTLNKNtf+gqSw6Xa8tJXHCXXsTAM3pl
zHDEMsaIIHNz/vnFilcHpkjmofb4d9aXqIUbp/AGyAmmqVpwpHeEdrdTcz4VdUXRcJl4yAZ84syb
HAsmp9p216IGWEh4GIGt7duDX1fl1bxKGVyck9+36IgH3h/rkl4VJOxnm8rvAZludH8dn8PXzEhU
hYGyJCD9bX7BBWeEFOke85XHWuqAjwbGocWcEj65UTzJTlVQjsLOl9MPDjQvsPUUo7aykeSVkaIG
+ykGgCfme+gF3Fx15Qg7z5kjksYfXQXntwXvegxqeZq6pyuJFbToN63WA9eimg0gAuT6JjdYGUPk
+c2IYLfEdLC3w2tbgstGo8C/2oSpRTSYaJ3+XYPNmLxCofPfLlKlQgXkuKbbsq8A2NaIb7xMV90n
ZWF3iolJoymmvsuOMJy0Ycrf8icfkkvgAUTFt/J2qRcQ3/qCrPdnKZeI9i3sQmh+Be478dporBpL
9p5satIRIrwC9CMol2eSTPKaA8s2liUjbJxx9nFt/TARLLuWJax8txK2xRke6twGMPlk/b1BRHGe
SZu9Va6X1C2yTH2NTW0gBXZHLUfPc2iAhO5NAS72Nh45mBWp73VziSh5gtrR+ipUFH9Vf/02rP/D
WYsjFEEK7NBRvGCUEhE1GauqBMw66yFFjTsi70Mu0eNIK7qfGMa8hqFEgnnhFm+W6F1aQtxdg0OG
IxjwUfMzKcOOkJVuEkbq1RDWn9OkLeNMS3fuGfWV+SWhRAzGh6fMGlE/g6N7QYR3QIxK6dVqcQtM
MlU5+xGY//uYTm0XLtqaPSRlHjqm099yu839gAGhxWL2Ijh1HUR9ppRuwNZpMvpR/rZxz//dEguP
vKuDF0/XXIQgy9ROpysKYsFrx6f4L35EZO5QiNFMFB97rIcHQ5dw12eILoXvmGEOliONIwR7yXqL
16ToBgKMYhtpx0eQTMxul5jnATdb3vD5AP37HdQrS7mmpdwx5dPOpkMsgt4xiVgmCWiWfH1Uj/9h
+Bioj9ShZLvzTMLJmk3N2CL4eovOpdLInY+K3ign/pmHCGunBfzFESpseEjKHg3iehkCfAWZ/VUi
3o4yMoIKVUfymu7I26xVSPCyckOsMmUaTr5tzPS8BdJ1OafLJOUzagBgCaBFqExnVGjt2+Z5i+1I
5TT8oIeYY2l93Qp3eU3tzNyjH8bk9GREeaWNocxghO2wP3Cj1hFhTfiqu6gKp+lZjlMgmSDhXfUx
UA+CFN6gRtbBgMoAG79+uJ1eiKjCOaK8W0W4gReHaCXCUJ/B624Fa8ZkLHCZJ+larrk2Yib9FvoG
AOeuNIi1+NXvPwdKqopkGg1foszfZDjxmyIlqrOXoy/ylsSPwI6IrYZyKnP+IgeQvyuSalcKF4QH
+R7vikiKvn0QwDJh3/gHmihDPxgJuLHz/bsEqNjskL5yDtER91ULq6P/ZYGHEDg5ff0ZUfbGoaRM
mehQz6WDIOJFkcdIku8rjg/Pa9/TWgDl/pcblBiDw3dbEmAnbe3iYarQqzEPNEO9jRwt57bxnZWA
4319IDGUZfP1mm4JDyXMfU4DAQYPkB3FbeY00QB59xjgbGlG8r1NO7Tb9PJ2tinvhWs4SOmzBPgG
7kptMKTGfetsXpkLZQlUHp9A8VIMKTtmE6qrFLpb0U+XWVP1wBBHo3/NFXPqZOF05EUiIxDbG97C
H+5AbJPvycyKXyra7a9Je5Z7O2OYe+QVSi/osZOTb0fBY2jfqCf4+JGPiq/G5zm0qstigoPpU0Be
+2tjyvAzzyuGvr8h/eumgpmTFen/vbVHrebo+hkbu+923ZRh3vuWytrwlWepcHgfbPDRKwKhoUJX
Lh7R6/uVNWDiquxtu9TY96p+awrfe/O+8mKDs9bHrjucendZixk4Blf9DRFl45ChEvonNrMRTUsO
6/2H4Sd1neYdf2EEzklCGaWvjQmOIZkJDmVvgCtaMC9esafdJ8uhN1Kx4npLvvUK6lZUoWwibQKh
6+UfLpoIWUB39MjgTD4vG+MvZpsHxCeljzx94f99vlqEKgMnUX8wirktz+L1l+K7uikt7th4NReo
uiblBEdzxzMF9vgIoh4bahlDcA7GhXOo8bPrEcmBT/3CjvH3yQN3YRcQtMyx4L4tWgFWzYGIi8KR
VVjbGPUlUQX/P0eIS1HH2KrnUOkxsGWviBZjoSFp8nhwTUSFHL5/0X2MIu9HPmH4T9GIWe3whZF0
aJMHYyQ3SyfHgwn9oxn74Ef5BV1zyPtESZm6ymd1QyIGIdNJ/WyDfdiroIVfW6ShPTtWX4cLU+j2
uE66a7kCMtSo/5rCd2kpqVGs0MoaRv20W7NfSTmCTnE52h/2OE+w7MqwoIbWNbDmnvBg6/QnuR7g
CJDHnEtYUfIUVZODf/z7kdNcKSyXvj74LocqhJGru3yFWMpYahsoyScpExjysciYy7Q73ArII8As
oYJFR71lwwhQlCVujBtyRbJIyUbd3eJCffIz8Gwb43GVQfEPdJRYYphXcfqDtMtT/ORtowxRcG50
G0BdXiboq/7cjRI1a3Sv8iYbPCCVn8/QbK0Hg39OZ4fSUoRle1/ayoq7Lf2lkUigJtxxdBQt9O7L
5mmfxTJ7vw9WkutKp0O7VSzpCY3d1ZSvGcIITYt2Pn7oEGn+cZxJVguO93vru6KJ2cMfkeTWJNJd
/sJv3zfP6HASmdXzRVA3SyhKiNkFKcthU/Pt9r4bUymUZRg4iY6RblptrByHp52NfbsnvE20u8mB
wziR6FOsGLDFcVzcnCuovgo9f4akCGTCYmOX85hrpZqWnydj7Q9hLmqyzho8Vo+no2VJ6cgN1eeN
teQqdoKGsocJ05izIfv0i5//XKyWUFvP/QCZ8GndY8BI3fsgbXLnfcPrR4WehH15/af6l22rWFEk
fOQmFYLAAGH9Cvt92PfXphH9YTtx96TH7X33AF0NEMCpsYiDnTPeDfIKybqHA7TLHByOqx5dUoJs
vK7AirIjcLuxgKOrFd0XcNHT3FA0/1+sJeolvXV18Bkn9hPkUau2mZdSqxXjTqukmwmngwu85+A6
lILGF+i38dOUENvXH26NM4fYdd28jI9DhIF0lOpkispnBaKpuJ907sOdjzk6pvkGHIuME2Cigc95
wDHdUXzWH9XojuhTcTxv3xnr9Qj3oVMDBFPfAP/gBXKhBWwGfONZoXXv8SzCH7UuBqDqGfWHk8mh
KV3R5cxXBWjquDQv/RnDTU3q+yJnsNohEUYE+oIg0bkr3J1vS0iUqe1+57SORabr41Z62pDVc8sT
46aoImvasjy/doWywtnGyGtdUag1xfO9EIMY3+z3Qn2LKJTDCni+KcSFEGjUuKTH/T6sbknUbEGU
KGdv2tUcRC7SscXxGmq8OvaCKaCsmyg0woHtVRZAQh7/mSEzV61WyN6/HQkNqQ27Pg7YQFdnpSBm
PK3z3G3I0mp6gl1sngvoArbASh24jDLoK6pRiyFaqOAQusKP04JQgN5BqKcVYiAfg4c5ZtusNskK
OgRT+KIEhWcAyhneANQYMCXb1dQjvHPRr9dVOwFDI5GxvIxgo+QREUUokc4oyY6+l5d1Y7fTiPA+
tZ3KJ/fx9ZnwmGn+6GAlPHxgVql6RO7qnlaUgwy3qLw5VYestpvwqlahZ5T+G9N/l6nbR9uLU24c
EpDiYUgZwDPHdkHqup10TLEa3trGYy2zF2zqALVi8HySzSCW+d5/XZkX6sVibjlDqW0GVEbeQssE
U+gHDTS78Hw+XLjmrDYb+5Y9pc7U9ksTElxiBfwVmacPwIkjOeo0212S08fJYQlPgSQaUnmRQ+Ug
qVMPs6Nr6I3F6zZPsAmp6/tm08RJ/UplLePly5L1tGFtw892MRWvxtmKMXi2YGWjtKZhPLXD8It8
6qBcSooHMDWTz+QsK6XlRgi2ppcX04qItMeyhDx+O7qsU2goFcKunMS9/wEax7ruUfG+N4iB5w77
H5UTiyXCrMfWtSA8H6TNpvWKNyjS4l3cVlkbgVYsH7hweqmYwe5HYacN30+I7YhigUdp0VGi4+xl
4TLnuEUZ5uSEw+eUC+iGRPcpM99gAyb4cZjihM+xcrrkFXZXruV6PDp4wZGCSPN5fxh2x0UlJucp
T0embA7O2BsaEaZkVWSx3ifJrOB7D/kWnsMuWXZVq0V24thnhXJzjH7Dlbk8UKHh+92bzYqSe94K
4OP+c66tRTiE+9Ctt1dOBxOl+c+BhKgRMS5PbH+9Myva0JYHLn/UQjT7ppinpiZJ1ewWyVnw6OcB
q7dSq0d04cN7U8Iuylcq4rEL8z9EPyt+a8veqX/GWHeraRaxTLYCb/MeeRbZFfYPWS3q69JkzANd
ZJkmlDKNGKYLWSyL9tPO+Z9rLGQ/E1dLLDcUSVaMjJIeQbXSxWkNfI1ucV1HJHjffXHG6EMyhH6Z
kIgZcr6mah5w7QddoJwdt4NYi6yo+kHSrHT5FchOekNwB3e0pKT07SXJrXhg6UpNnK7Kz39eO/LJ
fbWzp5HZYOTkRSxjJB0cfKZjyzoHZdf+Qq0xq8VlxLDFYPI05Bxfl64pYoYTcANy9C/d3q8LNygQ
rwQUr3SaWXjZPYZTzmjNoVPY0/rIOvL2G6xM0kLRgTvL3a3DvjHYBoFnBJnrQaa+5+a5WMHYKIpy
7BElVRb5379d7lTlkpr3VL4EEzvB54xCtHUMiWRrQoVUq+2SrLVeWEdwLm4wi61Ya3iknoQS2kbF
zuAZHERyRays2parxokqWQsf3fbhcGhZnc8E+7Ztg5Ea/rYIcMOP5VrPwYvDdvK2749y0dUxpY61
OYhql0v0Ba260QC/UZA2W1dlSxF/ZEhoLYi7N9Qjrx26ozmqhjJq41A3jFwai6O53C1Qdp+0v4t8
2AV1Cnb23liJTN/bWqv4iURxdcWNrg89qBJFbLqiLMA7NHtcAd5XhX4pBvp6SmK/f3HHZgNJ6AZ2
9wH6atDYuTGhO6zQbzEx2G4/tfcCYCGr4bGP3oQBP5xR/w9u2z0Fcz7dy3t20tqU2o+29MMSaZPM
vyB/hpbMRecFmqDo4D8zH+/dZ7FtKxki7WJYiO5ItPu4p1SUy8GFaf0n7Xd70OvFEuu+pyu8FTEd
NuRobfLQNXp70fkga8qISZOWJZwrHNzvyQPt1c7KqXwjMvrMjBB4oXJu7kGyxxNsNE1lJK2n4hIA
ivNn6QGCjx1ACbOfcaBb00yceRaPpuRHIi+BHYY7oqUJzMVyn0xDrTXUB2EMJepJ4Agj3RrvTieZ
CxhsiwaKl84LqlRJO4G9PWnbFsszOHl9y9QUElK+30/iXUoyGLkrUYEaYj7xdcdFkopKUGUDWtB+
gpsOnsrs0AlptkyvOma8zXCodn7LKxAvDE59F092yLcJ4VmXO+ucBppdpv0qgaRdqDYAtWpUjQ8G
vNPm1915SIc1NRgpYyVHQx065FGiuYJ4ik+TF+gy79fy0yXPgulDjnowPIgNE97Rl2Tctx0undvv
BJS9+WUzItupXRE/g1aV9e3yY4MgrZ/ugroFMLONiGrl4Bcw/vyzyJaLdT/HyXO6aRtSgRvhlrd0
1ubHhv2u72BiANMIjLEb2yJVD7Wp5R0cgPrin+z3WIhaRm85OWtIoQfr47mY4jdXTtg3f0CQT52+
LngzKA9ZKTlw9QN3K7DiqygIrYvBv85WXXs6pR1IaKo9EAqhQZZ+LQQ5d9N5z8U6bUGwXuNRGnGk
6qtzmQfAowzD1UJGNuwkSBNMFjM6trIbN0/WZ+5Vk9IIHNNwnEl0eKLAMU8S2WpPO63xd2ZJv5La
ZmpjdootzIv8Y9c35ioS3iymFnvgNdKJoe17zhaXaQnqnkQW7Ao/jkUzBJszrpdE3VUo6XL6VAEG
sar6IselBc+knTOd4DsTJcWrUs9BbCvNn88MfVy6RgT7BfZZgF1sdsRSIeEeCyp5zGkM20Jbcfro
irJKBg3lfMtQy7vNujc5D/y+n69xqlTKmuiMIgFErRlhERJRQY0iL2HK8n6MGkH8UU1Gfc2UxFBP
nGaobLpM52dyJXS2DrldS4t6Q90qTSyuTXTv5zQaJezxELZTz75wvRQsxMMDwEDqPK6pBzq+bMm5
NZzeYNkRlswatLGsrTBqRim31cbZY81qV8q6liOZGxkkmfu4PShr6gIT0ZMhfzkI+yYloynLdTa8
wmdZ6PvVSpFnc/GP3rrTZ8Z4HAa/7bELGc50jjgnJnkEuhZqOdHQoOpfoS7zEIEDc+sgJoEQ6CoD
yDLj3b0YE2o/HaOj7l3mSBZD7Xgbltgb/ntE9JsZQJxBXDk9AauR0ceZuI9PNXYNliFaBwdYbR6Z
hjSn2ahscAXCrqej5bD8Ji0iVA/hQb1g7pmqLK68IaZEmQhWu83I3vj6ZIQNHAl1i2SsdcXluFqh
0FAI3ViaUzMGsDAy+dzKuHjcyUJKGV9t7/6Ai6OajH7hZHcOX54QqOzPykA/72uVC72qZ7c1NEsC
oVJUL8XnHI/wG/R7fwhwIQQLm0W94jt66SsqFEnHP5/ceIJS2vhlQtbyk6QvAmKnpjYE4NadBP0d
6dVGdFGUQPBPlQnlyAauKIU986uMDx2Px3MuJ7c0oN/g/kk40p8Ozj5+ozO1wUHbCc3oMpqgLOQ5
jvGP8GrgGyl0OnRokbpjpDPqLIXjLhX05qbU/Vs5xdykagDTQdm0oUtRtZ0LdUCHzfQV/UKOiP/a
u19nzXh60DLliE7RaPKGI+/lIZ2cTY8hrCLU7p5aMTm0MWF71oWuM8fv4kQqWJOSZyPoXCx7v545
tsI74zGZ7R5bfu76Dgj4u5FqSI+5GZXJlZj+YuJR7aqmOHJIEXlAm2hhPm5n7J9ElhnJLLJQT28m
ydWDsbLe4IWOpGkamV9v/sa/cG+ef7z9Nv5ndxGvwfMHaMA2cR8bVIf7NRUuRwIqHbUPiRUYzlKx
IO0ufzQGZY81PGl4a5hUmKkSrRHUdAx0ARFm42C/n2k+wsT7Wa0h1d9olgtiWdYZQAgvpnl30MQY
vga4asQqNpILNkwnCEBS7QdyNt3VO5UJyPWgR317yuBG/6AWAq+69MBAOaT6+qDOAjM8EYB+8ZMh
s85dVP8cnh1IFmIvYXKPbOIfIipGDnEiWoARbG8fdxsEvAv2jXmanAiF9dHPsdklkPMCIfzncSPt
4gDDMuqFf+VTP80btMbtKNhe/X+jzziSbShy2S4kh/+5mlSU6/q/0l7ORgHHsm4XZC2G5BIykCcz
rFvho/QlLAKFZ4BC8gTvygDSGaE3vMd9zfzezPxNXOnV3hDELonwsh2Mr8gxR6dPQ1vjMBmGmtM1
GxbLxYLP8EjbyTVlqqYNM6ymtaL1YH32qnwqwSVs8FQEOKpRbshWTcY4H1oeSzZ6iv4N4JijthhH
tIs80880+noYJfBLqfnIp/yeDczZ2XzqWxvMuJH57C4nRpvg5mMP+q5l8XvqvYqwSVsy6mLynsdj
MpnQnj4p544ZtLcz70Lhoao/TySZAd2vAZ0bdS0cOvAfsD34P76WxkX788Mj/CV/RsuTebaf1yGt
84TRiF8cUQe2c/rOtogjJlrCSBgRLqS0Lhs4RA82X/OvDHYDugi21Vxlh1FqQKLsfRT56jRBtnZR
LJOMp2PmLcVwGJGUANnbbmnJRzU/TinksBgdfz33nHDmCCml6/y9xf1YWChR+25zsOsOhJ0iUgDp
Qz45tqetc6oYJK+P9agnfjVE0aVkcFKIN7PoGq4+A2lcTpqEP5M7dlC3umdcovrIrh60yL3znV1+
4ybt2E1fsfwVujrO4Vu9/F78ke2oydMTQ2yl4kZvvsN6g5s98sSixIBCrutY9P2akUzIslh7jT2N
HTQh+0hzkHh4gbaueqQ4hYgtNT8GB+Er//vxAA9Tob2vpEupDT5QD5BeyEWtlxFUDpDkvZiIDnnb
I4b90z7Ulwozc3QphmQUxBzQ0Osrr0egxmDnH4nI+0Lq7/ueFwCJiD2DSd7ROWjuUt5tf65vtGil
iotQQgMXx5VzSut9u/6/RSb3xfBL2rFyMX6uPDYXjmcN/UnhpO4kqgB7maQdyzJxR6nsDBiFju6w
xGalJvhy8AfkwNUL+bAzMWdzXxD7b1Lo7T8NN1+WcFunxVZaadYZTQ28HoARtNOVc1ljzkH1z6xP
GXm0u91GxCGrVu1jow036EoF1C0Go5KECEV4qp39h6Ea2Hl9jedr+kRYYngFbAqCPy8zd7//eutx
2WhFxrlhazURP4lWhtOVHoOrGUUXxPWYvDQV3qfkBl0504Ybg8i8Y0jYO8NO+nzYrNYmJ2EctXmf
OaX8gpkDhyujk+hHRkiYyIV6keVy7jA6XwfiXkjC8GkLVHN9LLDdGa37si8TjOWIton2hylZeGMZ
hXzCdREtm0hpiRM7eczR69DlbDOP+ON7UjaeC0yMGTpcRJEGVsxZt6DzFE9ZEQQ7xNA3SdT7nfO9
7xSQ826iR72mp3SGr+1lpB5sm2rbj57vKXlNBj0C8fWN8NiAnakRLNUcbNxhwIs4/o0JRivIQqxG
oP6hImuXE47s4Ldd+J2cynlSiO9SmB0HfZvxtMZ2XFrb20y6Gt8kJ/EPbUcJCI+1juwGZkbgQpsI
CKs7hjYVGgYNqeUB4wL0md3BsZAIekURN0W69fgNIwPuByqcOka5IgGCTB1dHYyXxiDXU2EtG2wv
GKwyv0kfQU+2JPqcS77T7pLpv7wNIcIXyopVpSVtFcZ/PoTDvkgH9DTH/492ImRemCkjW2jQaCfx
1q/jU9z9FoZ1hcB8v+SlbGATPDnQRQ5u+bnRTTLTFCxeOKcXl3qcO6LWATW6mT7kEncMbWAjVeRh
nHzYbMx6RKCvppE4vRoRTUrvQl2aNgQbXYk1VOyY0QM69SNy3SYgCsj3MTixndMiQxfrV2eyY/t6
Ma7mRvCrQOES8CJO7KxS6D9bBW9DV0V5DSpQE8wnNvq71jGyCLiN90q7Ky3+6I55xlg9iq4c7hZJ
t8eRRlbW3WnBZ1vUn7GJb5lxKe2q0JMFzgEjfFQSh2r7UKF5+kVTWlWn9J5JUYUw9/xHO3l103ue
O58EZHjyFSBEKOOyWqjqhkOHKJAcUKwykx8wQAfH08nj5sDGJcu8ymTQRrYX92T7le40RTk59RdP
jux4crhWtcZWIErMzhtaizNOKmFjsm/3QN0hW0/m0TQbh/X3MqP/XUz+3dFOjSOpgvnm9lPUse7b
iKQ+lzgr/NyasyMA7CvAQMg+jgVj3F8h6cDoh6tbkjE+H8g1u5L1Hk0FngYv0zv1zh/wQ86p6o8M
z7Oibz/PgMYMiPQdOybPMRCZMjpMNT3Ih7i23RV+VixU+yNQ7TflkDCgmEwBb+S3s+EBwypIocrC
99zB7ioSnWzWVwE90O3wjL58xzoe2rMQL42Ybx+5Beh6j8AfcWdVrugbYpkXc81fJsMQ7KSm1wuW
KZ6aEQRCWwTkZeZANlG0LbXMGjMB4JiE0GHMO79Tmeq2zIw2g+ILHWpV2qM1xJc+o5OjmyynYvYc
yWzswmIo/cyyl1CvpiMDWIyk2p/PyXXh2pdLIgzWHMvKeNKCniGKidH66AHllHPaz3ZxLwfNpKAD
FdPPPh6yOzLlAXgU0sKjJt8svTAY5phMvNRT08YORrIRqqDZ0RH7Cu7NkoSWNNQW1hSfvg5rzD1q
jTmWFoHU1RsqwpVG+lOFdRLJi0qJoM0Tk/XYl2uHlezr+T9uzLMLHDbBhA/Bp8bgG7WnpVrHmJ9Y
qWKRVkaadvKy5O0vepN/w/d2XVvDbpOdW5oEYLkacb9+l90D4OsN2FOKk4IwKUyY31y9rszLuV5n
Vulo7LvpGO7ox9Cp+q6HkPU7YwpaQyIL6104Siyb3Lt3jWrTNr+CFKHFrWX0Gvs4aYCTvpeTc73Y
HzWNobGkKCYnWKbJOXkA0ovWOXjDAUhiXAz/B6xdSUKf4LuJ04g28he6UsfvZs1K12ftdCNPC7lP
eTDUIkSVmzztqx1Tke8yoED9Zf2SP7/jpFLMG8JRkGF0Y7HAoKQLbwbjYkBdPNkDWL3yNvhXVmnw
kaV+884nnsJxPnueATbuqn0TItOlMTFIA2LVP7aYRFtwdp2OUcC68eK1aLAh8P8ONR2yBz7mklkw
vrU4aWvKCAVLYbtIc7R6g+2pQiI4Npupzg7G4CHRHZXyrHGqhvgMpg/VUon4Krp902q3HtoSUyAf
sdGW02JHfgjnKO7oasZBbKpqPOf8g4ekWjnw9MToBXdHOV8wRahALrCrJ1rP+YpPUhiJCDfga9/y
B9Z4eC+uQsf7ZYiBT+IbfWsg/rp2oeahUrRiJZizT/+nCuh0DCNMkUbVmL7jkYo9K9GY55SXo/C9
Cpm89JKJ0KtMvP6Q9asB+JNDqhk1OgnRuVJyDH7eJdg00KHlBY+s+vnMLsH80acFQxvM1djBVioZ
TDZezFXv5l6M/aGTz+UMeKBhvv39KZbHddL0M6o6gD6sxeZoqqI7xX2BTEwkGJBMfwFE8kgXoe0A
Urv4xYT0PrOF1up3L+eEi0Js0zBEP/3ZcHnYIoL6s57HI7u6JzeFOJZ2frirDlwIz6cvH2Kc4uQe
OO+RAGwiDIptsWx4EjjBmtcsf+7OIM556AERbd0Z6sxD+Gi2nCNwb5g3PDf1rx0KDpi6Nkge+IEM
2Z9Dujv8aJG/zUB1rK+e1BZvXGQrV1TtGXFs86U8RhHUxqceoWgzZAitKc1K4WgH2hNKNXIsi5mB
CWnmVbaaMu4YbbAWpC+j9JUlkUi8fmrUkl36Qq0bcFE3jvy19GzAHwzeGLZjbNZs6uwmB6xUjK6O
63nHPSijoaYZHsfya8f8VbqcYh80DsnlfwmCDURdRAB+JnLEpNhBOp55MTaCiwB47P6zR4WXwXhQ
vtDF83PMFkLuHu+51lxyefc6Tx1HN+ShI50uxtUSht8BvcL6CL1eBP+ch7KPu2RHCVHfelW1ORS+
M2YdScrTrVPCnrx1QDLYoZyvVgk+T1TxVcrf35aNOOVtYT+vkd6GGUKn7oo/7GL+D9Q51B6d0wvm
r7TzC/hvVA+2fwaXZRLQW5iBWeIJTeeWggVSzZz/eGO621UP/iSutBHtAUqP4/S11GCINuV7GR7g
Ua3UOgsQQE7cj2L6NcO6O87BMT2ru4xGalkVZeLCTQJ7RUbb+lCfFsYdsIQEUhd7xl800B51VzeZ
KYQ86vAGLTCqyEF8L4IiImyhjRI0duICioU5Ql8UKf25unOq9HjajHLaP2BkYlJDkOJQ09fSTAbo
rxlJo02pFLK8v9LT3yC5Y4Onn8nLdVDn2b8KV33e8thuPKk4iZbmiEFJDq5p2ka4a5DhZp1C7RLw
krUG2Bu0C6XUXUl4qd5MepArf9AZs8ZXWsd6uYfNtz88LgnNkiGjXSRVLYj5/D1d4FlBHC5LRSFj
kxuV1akm2MYQYNeMngfjnr73HvW1GmAZPt3jhQPXc7CP8MCfQ+o3DwoH8Ql+hbJr4WGMpLUBxlkI
q/px4fEFM66duGtGmgTvICv2A15gdUxf1utzfsRJgUhNcOGaU2qbWJldU9ZOAWGsQ0L+ceG92Dml
o6OSgVY69nxdAH9n+F2vcwXUCffzTFRp8fHsopPx877yHlW1P7u7P1UjrwSLb+mm97e3S4pwIbvp
zXNBg1xEmNmdZo+pOLs0JneMu3JhmsmeYcX+EYKCjQMgY9w3WA6voIHe4Dl+0ZaZ8yMvxs0cHxfe
WCuGQu2jjE0K8v+eeBYZUsjtsP3vmbT/ADLqJoOo9mfVTkWEQx4EHFOvUVpiIwPz/2GTVTpeM2qw
mFZGJrHEmivU9HvPse9Osdn76faU+EAoeTfyqk9uG2zYd/MnEczc9dbtGk2WH1Va7WfD8W1C6EPw
W7cW5rAF+xpRB+3pa0Mvfy80Qt7sBbSip1sN7ERxUh2P58Cz7KUZHlrRSVpkYSH4h3syAZBjyqQF
jjzeda06Ey8ucwcOr8GCOO6G57NlpQ/x7SoXiGWf3mEtY2yqK1eMdWFODC2qgM3FFnsasR5WatZK
XJqgFT6k4lXGtGnh4IgnracgSjsB4MwUZ4UGNr8zsZCJ4wokuV92uOxAgkr6oAyp60fHHV6AP3p2
VaFsrGtBzWGj8G8+FvGise8IIbHCJARbONLAJ899qb5lVnWFUvhMixuWUPPeAnmtzVeEJ9gKIZ6Q
V/NJJQbREr7WmNaIyBUnDOqCfkir5VmRIEDrs7dSjwWCy+RyM8XFhdePnVONAa7TmMd88f8O+14I
N1OcnOajg7HEVEw1X8KMimY73noct+EbTq87NijYp7S30cIe5nSrLj4PZSqFoDP5dxNJh5mIuhV8
pJt/3yO+PnQLKoioj6oPW9MbE74u9PrehUAGHiUWZX7hj+FVFXAJU02ziuq7j9hm8yQVNsFf+Kyn
/SOJaLI64SELP5EsAeaaz78dHQqcDw3HiU39Op4hxgAWy5hMcQ/0ZbTC39MZdYwD1ng0sj5QfQB2
68IzXhKa1aT8PzwUj/Pm1q5CBghmresQ3qJBcLC61LUDXwKWRoCAEJnyapNAkmpjh2KqxwRxKy0C
MwHw2GWmVx8+2GlQ6gzlpmhcP4L2j993r4IOvG2jhQOP8OZKlvGVJDk7YvHgbqWdxqRQQ7yIR99U
EXDpzqqOHCUefx18RIDFipBN/7CIKTZOAjjNOEkf0W9XfYKigtAkuhdOqULjn8oX2voCOzpT8z4G
HiwWG4vh4NPMfL2Sq9vnS4tKk8kId5c6/2VOKetARDxtQl5JGqS+YTugZ1OYrt9iYA87cl3iQOMN
/J0kljzQ2/1IAOo2BdfM/MgDLrt6/wSl6RWx6qzWRc+ve6yrOB+cwqQXSOXjVZ0P+ePCvbPqXMWS
VtXZM21QJWW+TgzFWuOeAjC7FeFolNJaaiPkIF9pzu3KYa8K2Xjo/T1R0dkQM1aY6X6VlrKvRJej
qcne6jyYqmYjJcv3dH+fahetxt+RRzOcVYzFYpjfg6fAVXFQSJm/SMcW5j73tcRLbxO3EGqny6ka
JEVCJOL0Inz85MlZVtIw9PYC77x4K4Y9aDHpepmnwlXyb4Fqk1N4E2oxxMkjUoj6aOmEi/SQ6YSR
5noAcpeYu85GQm4Juzm3jnHsQr9b5jzAf3zly0wVB4yY03BjmfyUMDyfngG4s4onb4gaLGbygpsV
BSD2hu4bjZ9pSGr5VPJPU2+pDnsMd0B6tHLSx3bu+7zfMXdNv617FIoBMIYxoKU1CVVc+Zp87CNK
f5XuicMKLqU0706nzqmu5PjfETJhbJbsvQp9grxva6/yc0w2DqBUzmu1r01vLDjjMTJJJjLCeDk8
HtiQxkdgRx1aqxeIH2Y3hyk8AlY7yWoAQz/ZFLkfrEuEiu9RbrJrkAbWju8Hoq5d3wMzDb5XUP5F
o9EFk3HCUnNKhUL7lZ4qTSGKH+6G16qoAz/AwKjTepzdnY7+okJdRxz9YL63bKP/Mqauk9TICrq3
mfIcl/DIBTLWG7jAHAZz53cAOVhm5GVu1qj34zNUk+M2HzkvJZNcM4rI9oawKXL24rMS8xnt6h/X
nV6Ix/EqIZZGF78lJAH1ycHh7Cg7gvQWF4To/he5f1znL3fKjwUKfdKhDyx6c9PAZy6GWq62Xocu
GIrshJ3wqoFpd+JSJ3bGDMH2rYrF9AlSP6wZd8+hyC65eFC7HCSqc+m9jPvfR4wEWmyUf8Nm3E10
7FqPE0DPSYTsk1SymubkhMSXzS1zUd+JKsL1xmgOx4fNuuAIpGMLW/lFrzexH3L+3FkWIJg/T+4M
QKInNS/UhhB5PL7IbAm1DfRavL74y4ERzVdOzVunnYyDxS1sFyarQw6MfyVBp/3kA5DQDujcX4Lm
5rhPGjlfoT3ntx4zM4cOJdnT+QqP4QTpiRETwD06OOZe9mWQ3MMEaa6VFKcbQKKRlvOQfLsVliOe
pGiCR8nr0mbrpiXWiz0hpKrRrpQKdIK7cwyj4I7TaUW5teO7JuhsXJ9h9rEnO31lP+8OpvpveHVt
3DPH5dJEz7zv+sBKNYvMc1G30DTf/416fm9Kjl4LeCDgiQi44hojmq5AmMhEu1xLfcfEZb82WD3x
YQRAAd3v33dP4oUQ2G8IwDEDTrCMfQ5UJVOlWOU3ObjUkCY0Dvz7GuknTYf2Gtre0YvJ3zY09K1i
MZ+nydvrlTD0yIlM+bzhZJkgB3bvvNvPhed1IhvTHUec2ZoKZvp8aZOVeSGllBUM1+8rJIz+Smss
5AFiqiSmHTvH/EJnqFTuSEIhoVBedOk+qV32Kx4A6JamjhrVvD4M27V2IRZMQsgBB7oCeNe/szMH
+OBt7mRj3AdHAcPtYpXP3dp5bqlVXNDbcKjd9lcdxsAA1NRUZz6MUPbexbXlt917tVaMvzVEcALI
3kQKiuRE/ZpF/QKGa7O+pNnDphmVPZ1M3/dMQBSyWka82GrZQKUo7IylBB84aNwD9cGBv4hApCfs
35QafdShxTqj7vL1b9lN3E57cdYf9JhKnR1dWwZSPyILiib6+O4RnLW8owwoJVHp0XbptsitdiNq
bHGwd390WGTuq2YZ+sM9gb0nhqDDAC1gDYo71HU0J1dgrmKMAGtpijRQleW6rJotB9Wf7ot/cpbC
pICekS+9zBYF1+H5G4it2uCY4//momG6COrSJShmxL6jltJZ1aKT6DTa64zRszR6wN7bCrnj+LsN
mS5BgFREOep8RTGwI4DaUB1YgutnprtOBHiAfcd3irb0ibsEJTX0FaJ7A/c8MU0VFsWnNKrmIbBa
MaDk/AhJTGeYR+6YJbSOMoXeqpoze6Jw5mlCOuGAYbM9uQGjq5YAoBjABvEeycGV/aEMDKHpDAaa
3wwaOc43Cgq6EVYrk8sKBkz8TKcwfgEAtolzI2h9UNQpsMcSM3HnYdp9+IWuvSCnYRrB3OSr0VCZ
zMESGHlUfn5AZwgn7AknZejuCFh7cfyDOCm7dTTwrCkhrjrbWP5AxTMDj3waSu2VMbns9M8bZVwY
FwLHoa/xcdGcpIcSl0Rw0Ky1f1MCJqHIl+6O0ixCdiJ1P+7w59qUlEqK6tEtJqWKMw4Fu79MC7HN
8D2DrDe/bfqLPhTG3Teg0bCxWUh2Meka9J3ixeUpz5DUx6otJV+PPIGCsSGGizc3YzwLSEhaD/8T
ZHAaMzCcpr3beG4Gz5/o846pZvoaoOjr1pkvCoAzB+sAg7g1LYmGQNPuFCJoxMMhyOVYGKt9CxU0
6Yye/rgbdTYrir5CoxJcflEFGYe9tNWoRrVlnguprFjqoarKiMRXZvZfXv5uHCjx+KbVA0cgQtwX
YiYHIIjduo0TBvDRoNuOCiTPvOImMkxPZ7/TsPsHUEKnheZkyDQ0B6+Wc1LvByGGZjl6XJMLip/x
l+4MPQNqByZ4YrL5GOabogEXJjavRZw1brz3t7yefAglLTF8UZMmNi6P+s0Dl+eQ+0m4z3Hj5/cT
sDUCy54G/enQPOXLeZIw6T72dElK+9M6A4sx590LaAokTWrBIfvvdD5CQtBlOiCHv8ozNSp4ue06
IPKNnMDwV+7XAdOWa5okkR4ZAsFBGKPFHTG6+5PuXoX5y68ym/mpJrfdiGRQNQx4dES6zu95BBiV
P1RRMfQ/iXZlvPa/vnPYC3tFYKeygbNLRYrtPz023X/WAPyCT1cMtvBt6uomlMEVVdYZmmbxIS02
/74c6PlOl57iBjpd4fB5bjumDcCxPnuoUYSbYC7lBBfzneQ9vwk41GGPL+dzOjBjXKb1nGzafJ29
G5rgANtnrTjkt4Ko7NdgI6IiQplvIIId2cRERl1v6wie7Hp+SxGdOyWsi640SXKOp2jHQtRpjuma
45pAHC1zQ9wDMhbtE68auTA9JOKSBZAGh9ngs3lTdv/8e1251ik1bBdqhxJf2EOTcNsOmHUwy7km
suK4mVch+nC8Uq6sDL7dLHEPaXvxp9GuNvqot6E7SJmJ6CTd6Ij0sZR60j3DjMS+GWwDZ5IFXztt
QshdHh1sj8gyMfj8u2lab2iKl7L2uVYI85vbSS2l7H5J+2grIXPKzhma3m7e13sroBlKW7UkQtHr
F6gBjVDCFdyLClco9CEIH+Gg0P6t0rFxTewIWonCr3tJ1bPV+Pg6qP2RC5wddoaK4ySpF30taVr6
zsdjKBk6LsFia1wmvquoP5+IYSCuGK8ZcVGGEpOwp3hbdS5iUQiTnB9Fa8ynO689Ri1bTvf0rq3A
MclXtKTul/TcqiK8iqguB/Tdq+BEVLxkmKc9fA6zhCJ9a5+Ukie6KKaLQV3ysPmn/4umQTbj7U+B
io88NvSysvBVMvKbaqfA70JtaG8jt7+PNx/yug5D/bJzrbBH4OD152JiiGwV8ybCECqtzbcVkPe2
Bne7mF7Zk4CvHhNOkYmUws4fTn5FByR2nFazRvHQnhLv5RnwR7b/TWImf+nicnk6smB0cHyzaZpF
32gxKvn9GYunwlgtqwO7Sagw6TI2hipK/O4W89lGh5g6vyE1cdASS68decADdYP5OQjdh43Dv1yl
Ag2W83fL8WcIcLrkvz9hGyALmruCGH5icgjyHGrKc1Hmu13lwki/vroO7iHgxJgbaipQrA0YFoUI
7UHk9DkZTbKxeuvMLWpEKfn90rIvOB/Whyr3i7peVJBracBTEKjJvAraU4lXlD2YXnvSiOArFfjl
D42G/sCzn2wMwCJtzVTl+Y0pXFNwGcO44xPvmdvlPAAVrb3p/JCEPqDWM4h2pFNsSfpu1IXNC/LI
V/ybRWy+PXqr3rP9yKeMSPvG4UNjheGpAgomX1pPMsFr0ezn1CNdh27SwEYUW9GpEf1C6na8e3Ro
K51jTAkYPCOvXm3Qk9IV991/hITYLKdy+v8lQndpI7x240afR5tEWSUTmpJmMFQSVT9dZGQ4hsxF
cOOVJxUZOUA2/m/xUdij6wJgaR7QUBDjLgRBnoQfW3HfPNmRyLAJNlcIl9TBrqdFGKRifBo25xpo
x5tWGW7cWmt5IX9vqEO25pZmsBXOLJBbfUOc0Mc3haNx08avpfGWmRtZDqY7eDHsmh6H3KdJOuvg
Jx5f2qWV2VEhRsRyVy7o4W+EyMOn8x9My7KMQMkvbFIfc4d13U3xn5yAelICm08fNM9AmWn64Xy3
wpY7DqLXmhTgvW0vvlmgEUegnl2mafelgkGDjksEvw1PHykE1QuZYmTEq6Li/jLVE3cbWJjkOXTH
npSQIIQ7mDGM8f+H+1/K9p4Gp7VR+GHEzhH/HbYVjPw0QGcnIKPKVUrk1iYlrSkkGzupXqwZwYwS
ipqSg4fS4b8xNFXuoUozX2cuHfXxIwm/2CUcaE2XLoclNEx0b3cMBNAlDLgBZS368F4gyJcqNde4
RQLOo/8hxFxXMGBpMR3ITLct0WY93xdzFnFo1ONjV9/e9nXhkRGhyIvtkVUmtI1W6anVlXKlCYzM
tTQlb8BiACvRZMtyrVhXnJIMuJvBn25TeqNWf6HrOyzEVCkWa8Nwi6HI8BU9OhOVXIGaW1SptO9z
kPQpf33AA0A9dLyye/oH6i9SQhhDPRAXXMDwKIen49YFn+rYFDA609suiTdqeXJNgX2Oo4ihmKSJ
PE7XoDUKJoIBgdsJO5YzOvtP/pInDrLmhfFXgdJGNEIgzyAO2xQ7LxOFQFyPjwtmZ3fdnqbv5TzX
UN9fawakIMksABR2ZPV+DmgmIHlWhMgbOf8DslldKs7wcYYROXNKIPRmJYH56u80XpnCIvSiFsTq
Gmu+M7GLmE25PIIdOFcv02LDNR4XoL2NYGXBpx3Car6u/Zne7vfIb/LMCU5yuTH5AB3YKfG2CqYi
/0+iwrj+4efpA+NPo+AWMDzWhpOH4HbaynmWkDJVJQqF0/GMxZtz+dWPauzn01zTpue7b8ZMnGRS
TxQnQxZ8eRuikdOFanIwKCTVfOaUptZ09vKRRUF36Cngvdkk98PhYTIl3maOzHEvZ0yMMvLBUJQ4
Wa2VoN0Rlk981o/c7Dlf6WyJY9zFuAzAFIixpn37ZF9G/1hEK0Rosw3Temb6k8RBK7VTEBGysmD2
N7JWQ3b2LdSatUEgTr1BLUhOAL8WAx9mEuuq1ydb17zMSc0PaHV0i1SeQbaWiJxpB4LMZnWR9g6X
FWk/zS1BO4fH9rBV2t2SHh4qlEXTcwKB8c4889/vuerIKQc6CXas9Ze1pHdAIoYQBzPtuEx1x2G0
3UJeWzW+Bvfid/beATPWU0nxUwd4h9gPz0e6aNQZV2BG5JiJrLUfRMawTiOdgws9P7v5Aody09F1
FSWc+mNN65IAyIXi9lJGwYm+yaEeIZp7T9h4kOvb6dvMV0MwQaFgXrGvG/h8aeUZHfhVls1Wfrpn
C64f+F93tOHL7tp7otkA83apxVEYBPfffSCNq4UzhswVOtuEsofrtpUwQoYSSHUgq6rCLyveUbGE
NpV8az8MMAecX/lZA4Vj6+tHPK9u9L8a8izd7m2RdYbn9T4HHWf3Sm+/mMz1CAxpXpvILUsojehc
tKfjew9pwDXY54SVL4mqkggNcyqOyRgicTHV4urp4zERhWODDtlAqV0Lq6xWHmTHa8BfVpUjvQbC
JPRBN0Gd1ed28CXfYzI1kSOEYpXKTBOrIWxzdvXY3mJrWHphrn/5AOmyNK77BmHUb75HrrnYgo6V
ut7XQ9cRRWP6HI8UKFIesBUqkV5VVn29GdVDud47oxGpIddIL2qz7sMD7rjytq6NjO2TvoacvQ6M
Hhv0626DfzbR/RSs7UtYsdQ1aFWUPld4DK2Fi6llZqGUo9xnlL1J1lIl7AfE7oVHSN/8VaMDbtbv
BHiNr9jffGeeWk1jrsMZkeIBi7Xb5qb2b7PjrE3hJoSQM9BYo9bhs0a+Afx6kBi+7DvcFPaVLe0Y
2ItHkdLrbqsk+wd1zC9bTxfo1IZmFllK4/ZK9CEDPnnkQZYcUuD64+7vw0VqhcCTsWHzswznxmM5
r/tAEtE2TjBIc2P46CMtinoHYh2WTG6ceYoMe/TQirPzjQjDCmFJn54aPyxTc8IWko+ySyeBXPdo
63LG8+Po2+OgGtd66KXYGOBKyJBE9eyD5HizQ4qDgr05LOASs01Xkd/hiYUaE9HjiF9suPUI7yDg
JjpIBhzbE82Zo8TJ+o5Y4HiJkiRxmRkG5g21Dt7Nr+Q4NSd5lu7rpVUenBfOeaklh6Cw5auXjomt
MYSfQhac8Hu2odnuD/3pQ7hSygSPL2wdAj4axEVexHlwClxmd6FDwnIQjrX0/mTF1DkPsmjog0fz
6o9BEeI6kIx2RRpKTwfq0Yqd1yBYHH2aPmhN5GDelhXLn2HuV1fhc66VFn0CaWu/Fw3hZvpocK/x
Jjbyz6rlWgPSHaWZ2Rzme0HopST2bVRo7tQ6LriLYO4QiqgcO7o6R1NhhZTUAiWM/wSnRgyBii3Y
pxjb5mVaoJ6tECllJFfjAV9Pj5SLpE1RmTG6WIB0YV3D1OOhhzgXI2szWZIT8B334hKNa8hcowOA
WDFphHGKZRDmcETThIEygWsO5sIKkpFh/ecDfUNnIhGUoMFa42VM4F2MJJRKbg7/NgDzhK0W4G6b
Gqh9U2r3db+iIzWxqLgAjpeSUVAHXJ/ePy/DPsF+6XV0Z6UTGcEgjwWCD+pTEi/cg13GcKmuiurg
I1AElTT7BLK4A5iCyQjVX/+6c6mFXU7Erg42znW6VY82eaSkp+7lHqb6Gf6Lsvgzlyhue8pUJ2jw
LXee2eJhslDOyuVRONMYEwy2sNbTPKBlpPvf/GDZ0ZqyDzE6yni9wWBTv0rlizl7yRn94C/GB+0B
3ogMEWRMLQMe8K/dwc8MWDynm3+eo0hjrpH/XYgdorFZYasrB/Jx1MbRakInJwjnd7ueeDyNlvyQ
fd9Uj2z2L/YhfN/zH6BThIAAJhhyF9M0Y3G/L6YT80aTOGi7LLPckB3H0mcs3LmrDojjZMHTHpkM
AJS/QXBKxC95kKLkPKhigwFxiBycgxEPIrd3D6F99QGmxe5dO3rIU3PIETS5lr6Ne6UxmJOhRBab
e/3igv6y0xqZZz0lLL2ZMyfQ402Z6dVQjN/9wSEawgYENMRrfG3LoymPYImzZZkZ0+fjOuYVIIvr
7T7/iryp35XPtJCFSWjI8OrgAQG5dvrtY87VVT4BKbTbGtN0ydcQduzJxCduHXk2wfDdilsl7aoS
vstwvVsiLTBq6FRMvV6tVHUwJ0TLgu3kEQb3ZmaXfk7yhNrKY0wwiqfjbIBHZ+rskhcP+1K/RbFu
ZFGUUltL4n4lLXtz95WDfk7ziU2zg5g8gZWSC5wnL9oLXau0eyzRdqHZaUqiUsxN+KQgeQ7wdTkM
1GVUBj42nn/ZEU+p5kjE27NgU2Fga7DNr6NvH3OtSLTiqM1JlzIyrdUGh3s1NkjdZRwl1i6DdFS4
QRED3biDcPCFF8sTGavWaBvkKn81y4bcZfjtjWiDKjCB8OwJxLiDFG1Hoq++yFKG3t+jZV7W+w9E
KOvJWmUrJ0cuSPOGzn7e/s6MJkCKzqxh1QgvtmyoJswpg6wwfD3usni7TaASQPyJIhY2SLCZsj++
am6m8BH4A0TGMBrnD1FKm+RKJXTbpZhEm2my/XPrf1iNNw+IEO6xrdK4RmZF23Id3f+9s+STjJQe
sKLXsHpyeQOsKiYh+vCJ+wZ5U2AhhaX3d3DXmPh7Sz8BKYWEsWNtoTOPp3Z0iO+uP3DbFL79rLPH
Yq7ewaJUcbR6JCAglSIfJtoRmMFfoYC4+j8nRB37L7lWYFKpgJBPinwOSca3uM+qhau7cjXElgp0
Lm5Dqzxdkkytpt8BWP4xjtejFi1FYXTRcMDlqUeEyz/Z28KyjwuGW6O9XSuAlA+ZK4YLrg9Dant9
5zPmZ1bJ4Pfr2RUACYdrsG/1Tc3VTv+1/x3CUsK4Ohs22lJuNex3/RsQW0rPVI8njnHg/m47g+gO
aA0loofmAvAsQNRoymre1Y1oGEmkk1g01Wg2j8CG/eNYpUfqu6386KAVSd85WZv5DxBHuKUvdgdJ
S+qZDRfK2zicZVvHM9LEiLABoZ8IkKBipHCU42sqQoRfjgSo3JqMuSV8bk/dAjqrro72d24G7FQ9
eAwkJ2ZjLHmluXbOnSf5s7Tv+zqqSxmmpWdzBunBPcacgF33bs28N3AsniqRcYeufhLmUworBQpk
OFnseH6egPI/4OvRz2xSIj9ddpuQKdF+H2gV0kQeqLyMkeGnJsSkF7QSsBQMBuRth7zFAQgZKZXW
XoxwXkt0BpQK9ZqqoAs3NL+1Q/nBzB6stcgNpMjXA3e3CSApWSVwmiv9MZnx4KC3nDX2OUCI30Ce
BozjBcp53vB/emllmiCV2evyL8BzEqssEMKxpcwoAm1+E9bHvOLNGyrb32R9HlEAl3Ezpttqy/mt
Ugm/vqJf/CUlhJIagSo0hf3AMZObKktftgg7NBJLI4maRmKewTnDK0sfO4gzMWmSqwekmJ6WPkyr
/hdW/DpqzAGkSkvrOe7Nnrj9RtoAY+gboySbrK2/sBBkME9b0E22W8ZQLEhPgRNSAVK/12O/to/M
EWZ01qMqFPpItxea3RcCE6Gg1eM6wBVJB8hu/P5j9ExWL/uhb2prpl/95+x7gN9n+liLfyKA52QE
pRVDhTc+JY7jwTs3ovYh3JOgseDSJDpNuwlyF40916y63A4WkWPsvy544S4APkPH5NoMofdllA7u
Peq2xFsMaoGFCawXtlTLrkj1AzsdAeGvufepBTPzq37Z9ung87cJ3FOiMBJHMWBusN4Dft21vzMs
TrFPrUFfHXGbjLPw4+OldvEFwWwdduhVkGeSdPxNaU7sAb7DztrFDWDeO6RP3fgHkHmKsSaREoYP
wLMYJJk3T2OTIJdyjzwJP7mH1O2KvgN/mc7Kjb9Bx8IIGPk0pGLccAsyj/gx77t0ckoJdCxrxKQI
otYscqL/av52xnK7Y2uZscTehIBAbZSO94PfNMZZgY+JkRSfFxIgg+sqUtc227pyH1w+MdGb1+Qp
dKK+RB7bMzxBVwaCgYO1/ty08oFohlaSkA0lPcWUo28SHseAsgFyVeddTtyV8wQjgI2bxV8d0J3r
mAmHXrthDk9AQaxBylDAQE5SDQby9+5CiIk9pf0lqVpyZRMTLECfSJ3l8Oa0gI/csvCn2oNr/rfN
P/3GhQ3tQFI/l2mzmZ25Q9QYvhy/d8OS9pSNeIzgzV2wEv4HCT5icHzknpwnVox2b64dqZXnKQAi
wBc9xUvnaTvwn1h48ihgFGWwef9XhuInxH38PmNeG7AsFJlFDkuVzMmquS8IhVor6dLTXU4tPR9z
SPEw89t0S5whk5XaysTiqAhiA8XYZckvBTo0ZWIsSyOUjRit4DDz0gn5a1Edqn1nJMQ9bTYKWdnw
TUaoHFaMBoDhdv/cSDenma6iQXbGsxBKyrRHPz18vmRVJRTqPRJtA1lzOr98bSqLAELwIf3d2X4v
T/DI9GzzPcbkc2tw76C68LacAp8+ABLwDBuMUGtpqfUmd+bMTth7IeS9PsxJnr1flMjUD5DWaB/d
Ql5voAMazRy3o41kqCgYTIAmd7/iJwuU28EAZquT/CHiHO8ZeFok8+TCXQtpi2A2BdMULlCIwrIN
ZtWOr+4gvg2E2qHhcYeeYEpIZcZaZ5tjFks45m30/Rl9YHFLFRUf94jV6aG7zsDZfdJ9hQgYfajU
k69dHtINyxYe2+DhkVOwA0oKdkpGvVu0zF+1psSUdqMK/pXVub6PtdJxwH9mtGjzKpWQZhKpAgmY
FQ8rdT4/kLj5eLQYX4G2JsjKF91MJDuEg32+A0AN7iZ5pjOQF3vWhzeIJYMYmgHfFbp1elPqfYqL
5lwWK/X2ET8zismyXnbOTo252KY/gH4vLcDarfEZF+XxHAOE/15U5pwE1U//H8iim7/8YRDDyzPb
iRFcWNv33nAVvRXkzXowwVTkruItLNjfIQZ+hIPSILU6gBwwmPA1PXv06QPUP8brJ0kHrATkPkMR
pTv0Z8spR/uFg6g8VtrfMGjpfmEjM9oA3CQUi+XHwX6zVDLc3NCtZNQT/pG50krHx6C4VWngUjv6
aHXjfObBweKYGpC/g0z/pZD7+ErHiGQqWCOh3XPhMZSQNX86YDFrAzyGalFXS2MGmIB0DGnr9lkn
VBbfYiAo4UcqgV3b6tjlFihJu+lB8XgE1o6fyKA7GI2yH2u2Mol8HbtaTErepgsBIpnz0fC8YbX2
f3OaJm9mvvtSkP0wOvkW3Yzr7Ffc14OR3+LiYhB2pQR5Opca7qLfwfjiqV+kQbKP/l9wSKYDfQil
6MjXDTvDmkjVN8Wvlmv1Oyfo2YpoZb9v48peGn8sYABOw12xyfvvMAYHKOht2WB+jrK9fNyiuYAu
+OlveeLjxh9FYIrwE728PMlCs4E5sWIFVQUh2n9ox1CXcoeGr5AF305F6GsFg2RZ00zfhpaUfFLK
3mGVvkdQ5UV9VwGxFMDztLy2eU4jVnUwHAKIYTw+rUYGgaLt0SD5KMgfW4m2Td1Guw3h5vmiD4YD
0jtFyDzIG+EJeJ/UB0baPQ2J9U/AzGbIPN1hbwdMiWkRvlFsMgBs36pOBs2PHAyTi+5JcXtypK4j
TIQAOXLRR+wO45/lLUYdXOOBl69fGQ7oKj8gEm+olP06tjoUlo57Vr66kmecAFBcGzg6/I1596/A
KpbYZZfsEycMRhurgHMcTeLQmhKv2MoQiUnrSrGna1EMS2MjAejL9zAAaLnV3jOonN/ubs0TRnGj
MKJkev2VhI8CFdniUgWRgpA73sZg2EYPE1RXCdlQKqbnqh4m0sWyLGLHWiaiZj5/G8yaVVFRcNOj
q24EUQardZsYkRLBL2ImAVIy0FcMOLOl0+kmK4LgySrOcLyRPiUrVq2u8BM5Oku4T8H4WX9roYq+
JPSVxN0NuCH6k3gaYq588Ymh9pXxliVe6AWwbWl3W9oG3gi6fbtAbV25YzV49EXG+JIqksDUaCa3
2U0vrpmeTBprVEWUtcB1Tw4S9R/imsAav6jAFqvyy7cwE6rnBfO4m/6k6bXjFIAwLpWh+llLf8Gt
u7ipItPx+q081jq8SE2TyZ4KPkj+NYO2xlpJiF5SuluaKLPpJclp7sGE5N//axF2+/t3rL4GBB79
isA8ADACrDihOrn/FtQVeSCZSFkiX1CWMk8bfwsVsazfWCNAmHEIJRbO2uM5nPbtd1PKqI3YWYTA
Mkzy7aGV26cJvqoajl3OU7YN60t4+in9NmbV0ML/YY5e6gLgqqn3t7Pswy6Yp/uXBNuHfUfs2MzZ
HkNFOs+6kwU5OoDqvdmNQuW7T7BBcia9y3GJR/vAtxsdYKFUCJ9mpoDPbIv/f94/Fme65gGAi+H1
El87fTwf1ljxXE1gGLpyHP21LqQjHRQPYLvHRj2x1sBkhhdVvdPPhaeD1PzPkbm1EedUrp0C7z3x
D2eQgD6I7+pMCB0IfFTuKyjxLt0HN/u8vszyEw/eBp76HxIAL40xz+gRAbT98uMlDl6Abvww4K3K
xOIboKMUwmqtEDjiP8jehuSLANO4ZNNcacq0OfucDsL3vSHVi92bg+hKQNkPWiTfziJ1+q093CKI
0dvYpvh4DwK+KNrBtScc/+fWJqSkZLpOyyElk4denf7lYZYdh28xHO8tXdJpyf3vJp1b6e7bZcU0
g9hz7G8MNoiL/ndQcZJLDlA45iah9PoySGruD/pNmiMzRTn+qyzaeEzBNsGDpEZWsoiI4tbLeIo/
hwDdryu1Cx1AD+HzGB1yGbFp7UT0HsA6+JALgV/OWhm2QOlgBelWFSySedcTvzq//k814Qc9MFKs
JLfAYWBl63t/J+l1gJ2NXTRJfLG+2OTv2gWwtJpaJ3QcAB8LwDyMrG+9OowpLqjz8jigQ5ea+RrR
/oE0C+RQpmT1ijv+XH/1WK0g0q18y2ijpnHomlf286jG/QLWI1rwmfDwcLrmuIc5jiZcTszd6/V7
vBB1UmOh6onTfK32DNlamNrEdo8iWmB5jbIcxuSE345/1R719tVNAnmUuqZSnnIwRoDyf4aT9QPL
nDq3247YurL61Wl55J68zJY4Nh/vFzK70aJP6DHKMoERD+HtPqS//YPKigQlhVGx10zaUVpHXNat
s+dFWRCBBQjsNppEUVdnsDZejdZznhaggWEN5j3jnnrQ5dxlDwJUMtMmoiAmDPpjQlJtuCTWNJhG
h08jYr0HMSDjNQp+jhUklb8mz5hLy4dY/K65hESDmYZpZPTjqcXpy2zi7XZJ0Ov/qLiXUnMZG4QH
BvNOGEbr/UhuojdmajVN47amQswi/btpuWt3eTUA53wWdvEvYkAqGhfAu7tZjQqAlqnfXsIVb/LQ
ldq1nhj9dMpB6sKu5qYjYGK2PDBuxFRJzvUAUBxIwQwS0/p1Jfccupz+Jj0A1QBgg74R8Fvbjn6M
IEvjprDZGEc+pSCqjpojtVjwIgzgWCUE/PSy97aaLSG6IcyWAF8x2J9wTK7/KFUQ/NL97sClq/EH
p42SDoDIkQdeyRN7QYeJOEqdPqinrQO2326K4Htkg2nDc6EQQ6QOwAz1Xwc8afVUTXcKF1GA94on
xKSb2xHKTXY9U6b21vK8Ut3B+JF6NzkJPOde8oalCT5C+0X5VtkPf/QlqYn09FjuHP3vYqnT8VZW
t+LFDBaugRJVzh2IGzLwDk2ZrjO1Yuv636++BwxnOLjei+iX0ejb1cdUEs13KhfvEB75qo/VImw1
/1S0XydvMMEY6MeNnZxMT5I+TxfVchqoL9HKUU/9BNfHIqEwR/Of95SSc2xUjfk/ujz/kWAw2f9i
h/PB51Am7GBgPtS0Eh3irhwRWE/2NsTPj053otKgtWEidO6Xr63WZWq8/RCXYghgV/pe9SOqsmqU
LYpDvOjWhJ36qYJhFe6HNbDoMqJY5P4Esi/7otQm6iOV6nUl01Ce0rvGQ5pAXK+MFT9kInxj0fdW
fiTaVH1bAlFDEdGPNPw5e0QCXxY+rD8taIy69Ffhvml6ERYE6AOyCMeWdUfQJN7xG3+klnEKNtpF
lcuvu7zDL+y+kcPH+w+mndYJFwhJImgk5hxKWSr2cXWH1J50OeD2pGq3jPpZcwdDIfB4rUiBJK68
30gXnhmGrc/DuJYtGPTiWtouINfJwqyh53aZVoEscLP1ExmqHMZjgQrkcoe8C7VcpxPyzDTYBnqa
l3/aUl+oHDsj+/73nSpzY4e56SZzENdz8f8KRNBcRy0j2olg3+1A8j7K8eeTPng0JYJaSvN54haW
LoVH6y8q5yW+5OpkIS7uOdz/waAAN4cDvQEGKBoMRidfHw90/gA9e3lF0VF885lucLQlaSF0Rumw
1unrTT9UymPsZnLGGeX1X1CUHRIPqW16wuJjMpUxNjp+CvIniz0lyhD5iE8kngiqzRBg3mYeM3cd
1K3TeMcyDEtLlNKzgjtqujXdMa8+6i4EaLr4g+PtlUxtXzRKXZZ+T86d9E+XJiHrswMF/Jg1jTy6
GNd/UzXA3PnB5RgnM5ys6j21Y4ClXdDm53miv1mOicriPKPQRpeaRYgxDlxEKhn1g+PbpHv+9gLI
MijKWpOnlsZIbphsIJ10ZMtrv8lLix6P53IosRtkxi7wC3G57FsmIlId57xE5MpeEhqhlQtA8MsN
45MWwAiEgCqtX7fQZS+rXm8T7M0WT+nSLoqGj6WL2UQebc8xk3dhT8cNbfsm3y3qUITga5gTLnct
EVjO2buaBKeQFL9S6yW4vsqvaBvVJ9MIyBRhwT2LbieQH9n96P+UiLD08cvFyMvb1N8Xhg+YImzU
6CZNuZXLmevTZCvc/ye8ADLrKUpfI+NDRq8/p9kTA6w8Xnt/b7AJAKdaNReROFFm71SmVxpXQ/Ec
ECUgm46yDyxEdwAURwTt/RSRl9zUnFipiqiAx9rWXVllRkZajizSmAWIgI3QaLWh2Dat7Vj3at+s
fFrvjo9dSQQ8MY4jrgu177oO8VM64t0Kv3pJx4WYlfi32d5E0hyP9ggJXc+3VJlDnFPKGAx+CbvQ
JEa4Ttbb7seJK/3mxVuZR4YGiHmUNgdMOUfWJfWWXpfqvCaDHM63VSZcc3yvFyf856HjwmQFQ0QK
AEmJO7xT1rnnAf6T1MPMwgijTesLXX9zK4B7y2DkeM6fe3JUrFekPFyX76Y8CsVOoBs9OEJ9uZI8
/RH6vmlWPRUFA2BTsu4QZ13dg/B0y+xpoH8JUhGhzYdg8azams9ZrJenUj2OPEl8mccTzDnlJGH1
+AXLtS31hxRSA9JXCm7M6l7LAuy4w1ywelQFJs+UikF7xEr9dL0RzB81ZJG36QYlPqFZw5YidFY+
P+mpkf55ohAw/oaGl3W+3eCfOzXoDKluFcYjoLiJI2ZDbihANd6fyWrfwF3HLhU05JVeN9uFKxzy
0CFqMWNDjrO34qQ1R9RkArv267v8YZV6tExkoUmfDn833zX4ImukhT7dsfambDkqfrbnCQMrGzyh
4IZDnRNcAU0xPaWArMKxbNMEwt9dl5OYpQ1gRu9sc7TTxv74OXlEcZJWicL10UnBi8aHuu7Llmo8
G7A9JbX9QVgBqks7vtI12WVoyP1ckP6QC7e3MM97VuOA87Q6ETCXIo7U8ki0gGj+oBS8VbG/4yin
/Gt2Cq2UD0fvk+xcGikbvCK5HfXUMgkI/MwYGzgKTmo0wWe4WCk9lzBD+vULtd7OGD+3MqHeRlqI
hA7X18Wgzg6yrKT6BHm3IN2BJDN+tVvF23lZrIBAKufTTIR+SAfEcDexz2Zztrr44TIoUkamd88a
l/yBr8hs19f5UsNbgc8sz+EovqIaaqU1ozoGaapI8EWGDblVWF4k3O9RIAE30FRsmDmMXuD7Qvw8
CXWUrVxHAl2rMWkYPiC4RFuNgY9C5hSQOhUyiVKMhPErsEMjlvBBU0Ii9VBX4NMmxsKcZH2tRtW3
axMkdCMzPf7hRMA8yjHVtbeE2Y2Vgo5MkAj9W+Fesv4TCyallv+3wiu99/CIR/DN2X28v62DY5sg
eq5MC6Sn1XZYMxc+HWEah1xOUg0hYFAPc1sBMhuxJoybHtHZH4CuuAI5vEzmfKOU3Nf149jpMQNI
QrOtck/zLt3C0OaC64EJwwfbpgPPEiGGydkHmRuvDdEAFRTJ+/RejtNdSmOek8ALC+rtPa5YO/qT
5OUgK1Clmd4YzuZ8MoN8/+lBf0T70FJJomLguq/CDlfxEGtCVTlWB+pXp86xc2fmgLUX115qj7QQ
NFdZ+J9tRm5hBq53YhSWefblMmjgup3E9WA+fMGcrH7AguC/XiQr2ExbZoEDGyQ1ipQkcN9HAou9
MaYp7pRWkxXG9h+ZGKs2AaDWLITsCeqWu4nPWFvjrRpIZ0OvE6zQFIuzwMbFmWCrws7y6fIDc/1R
sy8GmM7XNX5r5MBCPZdSMaaC3fVS6THiNwyC5mXmwHjcwg78h1nsRmQe0FL1hjRHannblyYhIz7K
LmWa2lrx+jxe373AZSQK4k8U7Oi85lHsOjxtm4byf8BJNxiNeMuX2cNhDj2keXdT4eLAr+RnbGUA
IjarI/2nLCIj4fpDVcZfkKP0Mh8Ds3BHHCdRjSpffjP0TMTQatYHYOgsa4FBd1d/ku3zHbr6R/W+
qXC33Mk1m4qDVDkwb0XKZAexLmY9h15LWPVQ7bC32oTcS6qVz3hBVjI14Tc3IgIZW9WdwK7C2Ehv
bRkW3KwyOFn9/z95tuW1LiKgB5uyZ7S7/gmUo2HwaLelf1z11n5m3PNphfZRMWgLURy0vFBLCQgm
pS01Ols+6AF170fNCKIDhyfiEJbt6xOJAyShYR58vftpOjadlu6qeRJYVgoaliFpfYZAUi3mjuQd
igK892NU7QD75KOeYHZ4d6lQMTniyapJsAf+x+wm7XfQnUh9mFxtGLWh8YWtC0iekcWhOUBYappQ
Do0ETV3iMV5zkxqgqp0JJKssBngbR9ReNe7Dc39ZkDKaRhdi18XUX9m7ST1Vpcn++QlOBYTpGWWb
gtlTjxDgXDw02VT5pzDY40N3IQJvpD+eqaSjgfegEclUTfZH0FoTKXmdMDbL+tSxsPx188U9ngdk
6/6mv/uP8pLE45ELeyoRC56mX+l/KwTNmJWg6JCIeB82wvUEeBuWsUrKCwJURHrxU9/dM65gryZb
o2edi98hZp1iQ3+3yRa7zMMYtSxWiPUWw2LSYl0lOqd5PqYQw2x4r5o4J/OYXh7HN9NeRjjBpB4A
4S53QNLATXsPKegVuk0fl6EyWTspIXnVCNrtCu8EhVb0sEMJc4pDYYU/kqgOx3iKKs5kEQvI1CvH
9uScXvG14cM9lvSgK7SnrxWLXVBFa5ZuJvWicDrUmEGVnkPu+Ygyoxzn9YCmKbJgS1I5bFwWdPKY
XQF7kUFhpqShz2jX+tZiC/+v9aUnWx5O8Jxp0WfFvoQLpjfhVKMRGyoUAq47pfXv3rSQXQzreiJc
d9dW1LKcFgJz4muNXT5dUbbeBJG8bnh80EisDSTnKsQbmuYo58AGeXvEXjvIAKp59607f3FTfKBc
6o23qaKzukhSOKjC6JfCqmQNkhpu1I61t5RJIg8ZNRxui1hHy7KlAZYEeJXkK/Kuq+PzLthgKkYw
m1orqNo/bkGEsv9sN/4DXkhUJdbQiVK11jPjxY/EWQXIJpR3GlU+qaOi8dEcPiEQip8Z4zN8O2ow
s/oGetvb2vZVLNAlIY6jJ0LkGvxfqwQYkAmC9+2oGlc0+1AN5X01VKulKDfPTE88N+xpn/22ezrE
BLM6x9pRlXE5CZrcKJuszgKPiqSehmUg89T2YFU5XRenSb1WldmDLKZwlQdGScsyL961ekRVXNRn
bMrFUHZkSIXMoODqSlGCFlTxjJvlF3U7nLrv40QVsm21mxPWUNCMTjF+0RpHhH6lHYZmQuMAA4vQ
RoraEvhC1Dq35SGEHoutNzLDk6gEZf5lFqYNZHb3l9TU5ClS0H/CgFpv5aVqcr0WxArXBSQ873iT
jJ1TsbCz+8PfvwtnE0FcereSjSQAF6sfXiOA6hZmPBJOExnTPAtvMunHx4/4cWhuh41SfVG/Eba5
NX2xfROawfdY4X1Aq+sEcZCXZdyz44ky0mTAi1f/Z2PFguMR5q8e9o5fY6Ne1fSah5BXBej/IfMQ
AcTyHxQ7RHqW1MCik2ZnRYLqJklOGrOV/PmFzvQrG0sl6vnHCx3vZonf5f+NluhC1xJviX9oNnF9
8GCsXvltRUDkOKiTDVRqeIPQF0PCXgLdzZVYQjhj9ehC4Yd0NqoaSgYHadCevVdQquYVjexb1ZXh
f6Uc3sLuGeosE9LHAuhgBDvNDF5KJSBNGjTLT3yoCQy3wZn9wr+2CDicdX+DUjn5dRrrmSZrmnxi
kdR/u3QbKLvn9yRNA+ouSjth6uOn9Q1fKnOmnQAx022jgBVFeHMf5iJVsgFM0XRi9EB9wYvLzY59
KGJf0daTlQhSibOeWby4BIsEblYYjq6AM17E8+4icAI3keTPedwdgAYrogNeCHfr+mFgr0m7P2uu
QR/8ruX33OJHCXzlVEHewMeOPj3+b+wpy9KXps5M/T5a8uVG69WuRLaUIeUldutBHHPkiBOtmrpq
PZzJzxfS5ljOV1+IBiPjooO6nzI5c2AyCosLXB3FgWIt85sQIW7JlGDqm7gLBTomaNA8rTuYkY7W
uxTLqG2zJhIgzK1Br0Ug783ltnan5kU3U/SbV5XdLzqVA8VvlUV9kR4AxafJXexOXy31IzIs9iQP
vWILSlDNp+W8dXeT9Cb/o5LD+Q9YLKmzXdQ1LuEHxgrpxIM2pA/HNKrCGDZBMhIV9n/tsksD0kAb
X7xTp5PqQ3Q0OYD+uJR/jHu2vSn92icVI4yoy7dvtnlrBGtCedoWTYJDztSaIgiwrYIYNndfhRSJ
aYE/KqKmrTRGLyh/EbdQlKJSwVPNtwTITUCerOR79U+T+HLMmDOTgUZivjK7TBUIDlLfWpVZTuAk
1QiYXn9OVPca0FMOP3puemcINdPfo9NfvwlTHGMYoNGrwtAPZkPxnNPS2WgJ/xVx4hFYearqUkro
ImIGWJd2l4d20VXn2LzysQ5mZgxffP/XS1NiNR2TsMbB3nvad/ZZeAL9zHrUqXszb3RcnRqwGOSa
i0q12AXNB9r+s5S1Qf78c4TtfnzRtGJa9mQDnMrQzdfVBumaZ/w6fnxiEEXq/8xi4xNixYYBKiae
/JsojTEJ0oVlejlK+83xLmui2kEijiQSWHdPFjlBXT15HV2g3LPZmwloNdO4xildNW9g73ZZWTAD
atmQUttFey6UO4TbsrSdbAgAS1RVjYZtZwND7jwOLI6XMu/2V3p54kLI4qvRKKlu+rtr2PoYNHi7
xfh6loPlYOXxxcTzf0CWjKZxkS6IPxBBRnOoucS6EhVb9GoNp2qaIHqGavtFf7vUGRX9l0j1U0K7
M3A3OKiu/KiYJtDNLUotZLaROWOnpHrStbD89R3G82V+PXPl961o/mxf4UdfzM5kzi5IrCUaifgY
tY1TeIaHaE2m0wTdhC3T9o3Wja3KIiq+rzwhKFolUP2P9fAFKWREQutyd9LvY4I18FLfPYpY+VZ5
ez6Gw+wL7MHGfBf32sQnz7TjGPD3RQ+NFWn7Za5dzriNjALH2BjiPpv4XAUpRr2GO538wS4pAmrO
a4gHSRhRlY2WNgh30mzD1y5Uvl2tKNabTHJMpuSzzeSKFnm0HHoxJLCX8CBhKBmAHWoero9uxWv3
YPpTWC9VId5A8/FyikxTmn0FR4hkdZ7hlPH+DDjle1jfuCcE+O/Rx/+hB5QI6rv7/pOfHNIIT8v2
j264DPGrFRhOoH5dQZkPOJ7tanrdGqZ6HkmSUaW330GunYLDnCtckQQTg+BYC1cVmWCzWY46b95x
kiHNYzPOmcXTpgrj6WMQ5QjUdOUnynbwRyo+ZkPFaw6rEuZlAwIapQX3AOx6/VWhoGpJgKXNwPbJ
FJYB+IV5FmaAttVbkjbeuedKObh0XC3LIv8AwAkqv2zg7Cyp9pWVhjCFJXKJ5JHpLoJEWjORDedC
9bdDe2q0h2gfcMq++IGbJqL9572jdzD0GMmXrD6ciKncrN/OcdAy/mgglJ2qHmgNSMR179cfW9zQ
ZBh9V3/Z8E2ISqBvAmOoLupLnIBzpsOT5YdJTMv0KVEtZPdGQnfwrBFIE5UP+hTVLHlNf1FSQxeL
ydAmSZ4ZmW6DqesbL5ElHD8imAF3EXhEJlRQL85apTJaeb3npdZ1mKTtUaSLoMSjEeLB6RYZTfk5
iCZ+lasuB0ninpqtn0JUS67HZWcMe18y1X4F6fU9kV3r9GFRlKdBEbYmqkqKV78yHyb6j6qZDROe
4VgWXNFvw+1oPsUt4YWDDdO8TTFqZ++PeNsnb7FmoQYPe4qkdAzAq6oporw9bnbCs2YhlLilaZCp
k6nNpY3hljSVdeyiq9z06XYay6Gl+I2SfuUjLcwNfGICtnYTg4WoatZvUG98rjpqsftSFTGDHV1h
PaPqVDeycm1zG7kczsR6JRSV4Gz9WmNYV0xx66qpdHbNRAE4Eg3jIN++M/ST45Vjk2R/CWQCs3PC
ItRS5kk1665N4z7E+F7FS6DAbfJ5ApB889JggxZYCX7LF48MzJDyqPZhixkAPbav8Nu0zDIwuXOH
EtU20R4OWxndC+A61LKdoSThynDSkh2Upqgr+6oTyVpgyiEdyOjX4dv9+iZ26ln4XG91rqRjmjn6
/pAQ/qulgAeuiiGuRi5hinYwRtqp2esZa8aJmQSGFMTyiEYGv4+aUJ3QQuGnoTEjwRuTXHBJndHa
NM9ILKRpdJdzPv1NkQd25zjUdCNtOnJxY7xdz/FblctksAo9oRTWXrsHolyw6fW2HkPaygahg3kv
YKVZNSy061QIKjDIKCnbdvr10c/OkSWnNoWsWSbZmJQmW/pR8fq0rAS5tC5+2ay/l8iw3fkS8cIX
5MfWXcYnMrNQ7dz8RWKOKhAIu+Ou7I3IIJMufvyRmwxjlIN5/VKoo+Fw1qWnRWC+PCCsXoy7WxUU
uWSqnZ6koE6rn11S5FaEZANKa4ngnmtKleovpUy4i5fvj4+/9Mn8FUYJmFG6/KkSXzIVYptD2XhQ
SxjSvv61iH7kWXyDI/DdA6yvz4xOpge8s/qSxSgFJqUehFJMycht2FTMalXbI2ps5krlC05BEshW
vU6R5t5igdfyXRkfWbNYOHCduzt9ER2LdvfijqIH0/F6PVpiJgSveMzaH4SAat2D3hO8m9jwp4SL
YRljzt3nIaLJFzp7a44vGRlKiEsMbih33krDzrx+Wzw97FC1CRnKtkZwQZKy6lOmiEGHNzrW6ymM
zAwR7vanJEzZh7JmgRzEVvPzronnEqMhQIF0KzrAMo7Fs4CWhIdspklRWZn2EDvnX+yuRKUem51n
SAozrREN9kTHqRdqBvobypjLic8E4d897oT1Y5WeQzi6dmTAnYkrYltLP5aUsrehkrS2UIWdlKP4
aFtxn7LFWF1umSAcCFHlGM2zVUU5/dPeF4Gy1/1PaNyEJpcnGt/G6yFGtmBicXAme1yUzs7HBe0t
bEF4ALThOz8yAA1JwX2WCm4aZaVIBBzpwW50Y8ayWRREC9UNEzbNFrzLwCKmow2DAu6IPtuYNjtT
vDxAlW4i/3K3u6BDssRdKEh/ermygxXlD52M3yIKomMIJkSOZRe7vKXXRT0EYeOO4I7do2p0ftao
VFE9Nw/pYoQUZFsF5WxoH1iqnINikPoT2pXIF1NDRWJtDNCzgevKW73HJu7t8OZP/ZavPZcAkFl/
bGBPoMJv4vhoYn8ICXtDnZgsiQb07r1By0NWgmyCISNBP3OiggIbDF3BaNoWongDLEJcsoK8zHXJ
CnoZtntgU90jcJtHSN3yKyjiHhpJpkJha4dTKLZRXutodyWE0fjXRkr/4FqmiQl2PVQrLOG5gj1E
zxZuEpd2zLf1hidzoeDgo63B/UdY/TQRSHIiioG3kDs0+iWpqYDO/rjuXiPyVYT8t+NK8Rev7TrK
rIdkjr3FOInYPJ77BmI49nGc79lsN8F0wypnQFgilVD+bPlZtYYoy9VslJMnHDUQVwmqQ8mCSQax
8dJH9TgwWmNkdB/Q6kXYs9matL9enwbC7Q5TzdYcK8LaRXy0t1KErWFZ1w1LsIkm/mr3lWv2DkVp
WX67e/imP5HIIMTDIOZbICFbOFZkL0Li5jgNhkFntF/5VYNqd0HmziNdlXAq1yr/1LcaL/DL3Xmt
Ug6M2ffzOEfBXz/IWWeyiz7T0mUH8exJm7+TmNBUt0vrelCBehjtRB57uJUd1sg/UGOkzv78NAlB
XprcL0k61F5BOanLspWNYwhQxdKIB8PfNQGTXq1r3wsunXTaPM9UYvj36D9pvD5b+PXGFgxO5nWs
qYPmhqWOP6UmtUKT5Q9IEucop4jSlZfytdKOqZp+dGHjAyDfBaPgKFJG8EThMyCO7V0S3d/wBJVa
KA1+Q79b4bRYj4DpTUjRLJVdeptFMpR3H2YOXPo5l3YHT6QxzlGSuu99/zD8NC3Ko+M2PNSMyNxk
Mr0+ll75bRBbHlJ1r9yRzUHrfNHggo6HLpoBYCTmkvGYHEN9dToLuiF/9LLYC3bOsDZFaIUWDTLr
G6MFQZCp03zO0nm/seq7lfsRMx/hjEDWHrFPJKrXJB0C6HsBo7ob0vBhlgrgQXfKjNO37i1+xZdp
GxiwNvTblebPSuJpXfhfNUozbiBxKicme4xCKv7SIajK1fWuTyLx7i/qYHrKLQNaWOoK3UkdbiDA
heCDEtp1NPxHVG0wX9lk3RwAJ96OxOe3Lto3mRtu5xUXmHNJSUC87ccEB1DfQf08f4z2Ts+eF9ft
tbVROZ4x3H8e0fxPTKDnblRAJUKgqcuEzBGfbAbrWSHqesvdKhkXCYiEdobiMcDcceCMkkZ8UtPY
h9TDhdlGnb6Yn89IMdHQdsRiwa9KkM+qL0dSKWaizNsZAxoFdEkQFhoU6rQWfCYRacO90feWXmBp
2Rfe8EBVTRrc7UFG8C6pxdaC3nrXIzvtZUYxi+61jDQlaSpdbKEYkUobBjJoAwA0EgEhDvJkidlG
kcorCquI1vBG639L6su+sCueKHgkybues109r+CWB7fgOYszmk9CnsLw2fvx/PH4dOr8TgffK0WK
nZocDSgF+T6Jj5AJJ6G3Fm4GC5yKjGQw/TnaaDtDn091mwEEKgTRyH3UL3hjXduM5eqBvJp7TE2w
+MHcrwTr+qVBw/kd1ok2YOpiiou+Mn87mjNn1V3asyqVW5AmPPmf7BeX4DQoS6simwx/ek++Alfg
jOpIqcapKUEFZuVl2eM2/fEMWy0ECseDHwjTRSwAEQEmyDvqvQ5p+YhLJ52UGbw5cdE262+f8qA0
MUU7C/f8YkrdgtiGCMJAvcNJzMArF3ivEIm/UGVHZsxdp3ATWR89rVWx3WtcqBghsZOdgDKvC8l1
+Y9qpIGzhOIxsqjWVcIuyZRgNg4Sj8hDkhE1OWsD7BRWlpIC9TtTkghJMiWTrfs6BphrEvxgzUoK
7vJrzPnyGBQExjr17UlnhZdLbelHnBZfLT16OCBCI9cXVzIJL7WwozK9GeSJJe2CZjS0bw4FhgEj
SDyQm37CJsJYkXhaTZGcrSxba/5b/pAAhga9aIgUqjC4f1LszGTkUXMJHc2u9F+6h6IS6r8fmqAf
HN6yVAyZa67RUagSzab3vYeq7wBaZ6Ixe0LvrxUbZ0FKkaqBsgjCpABCEfoThzCvUbQ1jZoCtb94
VmpDD6sGWBVWtzlKEYodVEC+CBHBmH91eb0y+WScGqxIiU7KxRlYOKSw/UXd3rv96ItUqx5L3xCj
PhAtLoi93aKOexYtE2l94AwDC/dWDPEFFAteZoeQgKuVwrR/+y/iU3a/07lI02QnhulkEzQX5CiZ
gu7VuHOre9oM0OJAJaR4zp0tSFMwV3D1tbTDO+7/6mtw3za6kyzBd4s2Vam2Lu6HDxhqintXVel1
va3BrDmo58D8bIvFT3eF9Z0Oxrp22snJOt4Z3D75Yy1wORmTuFjTROEvPNCaJrr1Jn9tjYaKzuu9
zoAPR6zFrOgsxYF6riOhp6fc8tdzxI7ofgiO8/Lv2PQZDoF86eTwpQwCVKkG2KQOGzh9jHg36Wzw
1u9fXh8OY+lCOjjCyUrdT+C0Q+2Xr86zpMNLkbgdU51gmjzRmJBP+OeQPxP92febTkDmsDv16eE8
jKNHGFCH7WRKg/viEd2koKW5Kmr3e+CZV2hi5hdPR2epwIHdp9wmiCIXnCWor7eQkqo6bePT9iOp
MtaJgeX5o2LK5veIFHkE5USiqvyL1I319vczqN4ZJC6symUYt3u8ZBOR+31EH1EZtHrXkZJGXgK6
fLQOZz0mqIY/dJ5jDjnPwzG/byLjRIGi9WxF993jcK7gP9ROPOWf2p7bhGSzjivIzBzHfnev/IOr
/DWZijNKowPa+DONu1kPeRZOhr9ra44O/ymQv31b4FDLh7AhGjYc83ZnKgKz5RrvDNXTvwtdIwAj
dkp0BzyPv18ZA9/3TAMak+nD/GJbYqTpDaujnoPM5TkbVTI4o2q55HvBozXpTxMPltaEnBJaQLJL
kQPiwxLX/Mqz80ilsvgcYr0+P8neMaEg4wjjwjiW7Jd16oEwg5j+w0B8tih9oVlUwxG5wg5r0t9X
uZY7KhgDNVb2gElCO+rN1zdGL6gewTnVS7ggg3QCHINyCEVxLMKqDCLFLYTAmPJuA50AOSCZgsvv
tInqUb92Pe4dqfA1wtsapXz/tVwhv9aJLKh3ofl1HUbJTUczgSkLBF3j2AkhAv1s3zw1upao/vO4
dDaQZpMs4JN3PRk0KVBD1p3Z6pLkxI+FMUVfhJU7pffP1duq9wop1ZtZAs47OoaqPvh/0kMc2Xcg
rHS5OOZRbJS3gP4J45HQDjrxJBmfaysk6dzXlBZgck1GHHQg+ZLmd6jsFLcJMjEkEKj//Gl6NQYz
gbvnYLnTzYyn1hyDDtliTGo0mV//Kyczy1OL5Wejot4cbgJxdO8ckNVIl6OXWdNvIYLDnAKLJnNp
HwZ/YZ4EBVEz8D0KE0bFeMYmnxV8Iw4z6dQ1ulFHLfxnuRwler/7MjBI1rz1yb6QeQF8UGwmA9BO
uRu6bluWpR7QuAxvWiQvqeBXUetgbRhwiJKtYaR68IxjGfPMrfAQ1qxWVtmHHKRCpk6ctXnLnlqz
hcDJ7yBZTatorwsDZULM+H9FwjO9F5b7G6F1t3DPkaTlwiUn1o9eGgJI4Waoy/iC1ZD5FvleFmXW
9bM+7yRwe7v3OK5P2aziprCZlxmwRXZiakI2vC2njBL6U75XWQ1VDHGfDevlWL1InEIjbcUXjHSd
yBFeGIpR/YXUeHrCksgae2hcyzRq/idsoqSSZLq1Iue/sMYDYkS0Kb1Djxh+QSXmWBd9b1jco9bH
5x8Lpt/Cj9ydtAFTbKZ2ouolhbXdRzE5dfo6J7GdpzysEcQmfptwmyFnHjWrnZju+OILksDilVkg
tf8PiOwGTpr7X8f9MZccrr9lT5Z44+fw42CSS3pGAezwv6fHC0eevVFBdlWV9iSxf6NN1RrLASyL
m+mFB032jOlWm8N9BCqf+qL9ugdb5tqci7Ka0clTu7UEDbK647RUOyZNAvQ6QH1zd+dWaWWEO2Gp
FLqWFUmu34AVf9oIQtyiwl6NdMGXFXKKSnZ0Q8sRN1H66X6Tqy/HppORnGu6PxolwFk8mXO97hH5
huOCEIub7ODJTY7jv0I7jIMnGrM2YfyQIlHPQZMwL9HZprw0lDaqaFWxr8wtoZf+Ize/J4LRouxY
ylw8RQJNwAYKqOTI2l7RNLbfjQV5rMIU6wYjjOpx5I/flZj/D/VNiccRwbHIjyMdbjpozSBuh1Cx
ThGE5UGmYOW4Wg3ru//FtUf3RYX7gFcNTsL7/ve0fWtgHIS3iJDbwwClpuMSUkL/JDz+bI+E4/jl
tw6U+sWtDlKIqGMxfvk/U4sq1nK0Bww0NBlSem0xdrZh9+XjO9K6rIKmMca+ktkag83nzQ31OVtp
11DMjnDtnVVDvcYGuon6vYFtRn3mLz8Gg1Pv2ANUnLi5hry22pjbtubplCuGLFxDB5p4MYwNcGpp
1P8YK0w1tlM7o8jng4xBrJoeIHaW6DF4QjIMRIIj2KBYEA1g4IL7k5W6HkUOtRYO7MLxtHLy5m34
yWR2Y9Kt+FmAF8nRVe9O9zBEn+pT3VWVe/cHA4U8AKsCWjgYv99eoX8oeGB+WCPoYVr91roHPSfz
uEFG9NH84FmOGQYXI8RaTizkyC+fsBvhS98Q9HUCKUrnIX/G2Wq5WoBYLXEdAot5VICn9jDZ63XZ
HTZHJiU0vkKYJBE/eEPGkpcglDp33qXY0vkiAnMAANirMJf6I/f/d7ia5ql0Eu/hfTLXwndpHnAQ
hanix6zltzVn894se8IWR45fAYzjihdZrsI2XCMxWdyoT8+36Nz4UB3Nxz9eHCJJ8jWnte+SaAD9
MpTWvoxNDvjSgv/OHvyL6nzxw+Gi7rPMt48/HeftKIJC27ik0Xi3DGc7Rig6PuNHHGpnr4flTRpc
hxgwAr2VNFs7podg3ikrFx51J+pKnOFDF0LnysMRBOc+osrniuH89NdkM+PJhPoojq5Od5Qcr7Rt
bEt5rUgafBw7wmThPzqUA7X72DHYb8F6svWjFtQ6Sn/IpPUNt4uaQY1gB0s6i1bjq7pzV5netHjo
lD5P1U5CuFLmtjcFgsmqwJKoKXPDRRtquTQXK92yfOYwyXfLGB2WdjCDku3BkeYHF2mlAS7AXi3U
UcvPaavdJ3OJopIWVp/0z7biZq1iYrAa1Uq46SxmWu2cc4Y/RVK5KgEdLft6xUVPVTTO6uN3nMb3
YxJwcg6Aw0YzH6vMDzpuJGCvyhwOYUBj/zQiiDBKZiyFfwYQcQtvom5MyuQ6d9UPLZyo9DytIh8U
XpKZorTHwU2tubdwAI3OFOxQkU/XCVaRlbMecQs+zOMHDbhq6qO7/lhLEyREkCVil9fgmzArYXtV
yHQdtJvWLHs8Fty6CSwFCxc2dZA/dTMppDMUT3YBQwRsJ178EJPMZJQRqPqkd4EsiDd9KbNPnCEL
YwDTsmc77AnDbs0CMqE/oJigRMDIwY/VN6Up0mNdFdmV0oVsJ3LXpbG/ZYB+vlialwnogXokw54x
q8HlVuf6DigLT8rs4pvEFaOieBvN9bhQiW6pUCgW5lgt+XmEnwkd5ncHhyNji7YKvmu3xC9vXK+b
Fz/u1ToBRdD6eHayjRgbIQP/55+k9rGVvAo573IJKMcgBihfdOE2AbTK9UgUnQO0bLU5Ky/S61Us
htwExoDMOIN+r8EePYaEc1SqoUvsGYSUfL0/NgP0dZN5/fJFAXPKQt12++7IHuWPezC27/4Bmle9
hnUdWmM1C4aMx66QCWp+6FsB/+nd69Ko2Bs2JYH2op0F1jE7ww+tm1hqV7HLrpMh+MZDH19JK+Uv
KysOToKGkFuNJhwIevdU6VWJpWUx+6/D7u3q1QKrsd08Ncwo5caVM+kQ9r+V7cNbJ3hMfXCWaddm
98qYIvtNkzbKPxTW2NHCKIOCFOEB1Q23Lvx5cl/1J6e7HpdRYjMTohdn6KWIg8hnnL9awIueBLi9
9lBt1+eEIcBz+0stJEXDGuhbSWz4nJ7JtEOMzDw3SqNtz8CNMhI1zG4JziZUjx3+eHwIR4FiuhW9
QYLzIixgvV+Hs0DUZNlQjCUZERyrjNhvLYZPhHJRDq5B6N/YULcLu//+CoG11r74jxMLChiKDvcP
aPtP18CE6Y/hpE+9qfxz3kFfkeqr5hMv2YX4yq+4aUQ7hXqL/AwKQT6kcPsGQH1ouimQ2R6KvZLw
Tr/COAvsRa565qri0Add+yO5k45pgbhh1BdsL+3uYzu8vfLnj0Tasaze5a6hHvMiqvxGZgIsr6Sc
3mbzgQ92ncjIilJJ3+1keF6NYgvbnvR5TTmk2DTg6fQ2Gl6ybca9/1zf+CREwwFsyZs8tpZ/AstL
xHE3nPHPdvtvSUIXe13opzWBIu4+GJxDvd3QOmLCIBSWBvd6k4SiYbFF3zDVVQvlTENMxA3uQOK4
tyD6SVn4rni3NE2BnXpozNfrMxY8qn42t67aVBFnXceRwLXuo2jfUMrPaPYII4DTqEPeqwMsQ8F6
06k2DS1fX6jHCVHn+iftzmr5M7uGvLLhtorfi4/g3m0BmdfFxQxowBUc6klmddrdDcsti0LMIUH/
EkvQ/6vxtcHyjqI4McN45JmKNK8rscK6N3zJglXaSzQTMRhplx+/rsESW75ol1cNpDJUwNcQ6Lpe
R35h42ojENsPdXr206lEcYUJHe6SYYbGseEkoQuheeyg+fRY02XuAwuMSg9nWOexfdZrELA6R6MW
dC53VNh57UAqkg6kMG5QLY1Zd4Bt7YbE/PB+4ISrcxoFk8cziVMbZHE0RJsGqB+LqBMODc+kD/Ub
tt4oZmIJXTwThZAtCtZSGNzzZeQYdQhnMm4PKQQMkpYVZmewxMGkFSEsaFmtwRJ5ubQ+nZC+GZZ2
Q67FnrtpXCmKUjc0cr48M7IiqEmi2jWAEdtjB51TTyG+5QVXUpIDzHVcLtBcTu69uGuUxeogdnQG
034mL9inZLK1gp3x/Wbd8CdqV2kc+Fruhmcph8ZAXELjobyCJSuJyl9VqlOciXT+02NfpxAWeeeE
f2RnHAsJLHXzXzNLLQOpoFTh+evREhasBmA0NePP91wGW8pkDEeyxN5Gj9daNpj5SPL86z3rzHRw
RyLNimda5me8AQtFywV3xvURhOuN+FzD4YGZ72uBF6KD0cePikiZs/7fbJXx8tSY+BYJsWd8oK3V
fXv6cp3L8Rwv5mDITa0w5PnJho2/ERVssCrQeUL5SfdtNWa5RqT+ciFYsKdnaJp/CkiZD7hoLji1
rEQcO0OXN7Ypa+VD/Tm2STKc764EBMA2gsELs4+ssyEdKUgRBASMLh8I40tXk4DkrGGCRY/vXxRr
lnST68k+Ht83XCmQxyiHtLN/lAxBw9j8N99WyjwLxuQTwYBR5jwpw2YDeX11tyR/stOwtQiht5sL
P6KAPIWim1ZAVuofj5zrpEq411LiXDDIxsKVDuFVT6Ki2J3+y/Pfrn2C8qTuIo40nmjmBVy8TUl/
GLssl1GxuIOMV3vQp28l7cQzOt1nUcp/UTbiPlSACUBck4AbswcXrVNiQMBa/9qMLhX/UM6RptqE
0wX50MyTWjtwN47JhLH0hMA0lc2boIovc+A+fFP9wr2aUQ/fCZiGfSCBw6R3mWjs92HQtBZ9BEKi
oKR/7rq0JYu6asoBX46Y3Wjmhv+WGPRnZw4KtbFWdrB88mSPuRigGmTW9A5V7K1kifKUFOAKkeNN
il4w0lTnJtofTX22ycFOX+lm3sOG7OD6IiN7pVWfUpwOWdeOa7XDTYbzA0XEoXymBz8NBrEyCORw
chtwdeiFOBb4M7OI7EYtxiEQZCd+y8EpYbzFuLL1rjmqfYifyS0dNZesfueMbLxSPN32mZVbpdK0
deR8nba8xgyElmr3YaX2hclu/w1WdVB3NpXV8010s+2/oZnV2afe6MKNk5RMJF1QSwh2PbNJjtQD
RdcKwbJ+TDUmkW7Z4MzTsWTVVKIqdB40GZbf5OpkXlzXT8pk0ipb7ey4BVgiVrd9Gz4cJGXroq1l
IorWpqBq7yt2S9XOhb7qc1VRzAShjR2Zkl0VonBUL/eOKkQSfqvkHsa3zF1AZMjGjFD6wNpZDsyb
rIc8Su2EBF3Eq1ECs+MRvNe6nLR0fISC8reR8ZKx0OJ+9zEQvIYRkwJ6aRdQBB8zFJ4kUzJqPeFW
vE/GFJbbk6OMO6WxlxMGuumas9e/G+IFb/5WpUett50hspnC5qtsUr1jhJaA1XY8FN9pDqripV4e
dXcO0hiuaKMDkchzcmQfOmeakngFuA/Nu5yodZbRwT6BHszEz6CanK8j7wzTdCPk92xZ5zvYE5h8
xBJzpmzl+MIXfyFmyJAc/pRiWL6D6VNbJfLJ6CxsTay7YQuUBu0OMPA3O95EK2DiTTl7eCY7G8eD
iyCSYN0jY5hGshwu6XhDhQhV+ZJi3zr6OPod4hqOCAV/BCiJlYUz49GvkobynGFdlJ7y458nlXg7
u2KvZwC4fkpE/mthDoepK0v9yFtvtrLso+tUjRocY/Zfz/al67cttWJrDwzt0fPCJ40eHYTYZtUx
oQY11i+1BPC23Gqo5DlXEyHZbP+2RjOoCDP8wr51622YS3ubKtiEGTNd98RwEwbDYdK5tG4ih96k
PzC1yrUYdlr+ITd/rjZy84SDBneI6a8ojuxEGNGrZ79d1KKvFU6Xna/BzhfZ56d3eDW5TSwBx9b7
SjReEXGsXo7AbOpLSvc4wqBwVKYNZYDJjN9xf30BCqbQdjgSJkuyUqYrPHIO2V6HBqpJ3+fwEBd3
TsrUHFMNgeOTgdfJSjhaEqoz4ua6eQ6zh3Tk9/DHSU2wi2+e1PMk9MU/IWBc1B8hb9Q6O96ELRgN
2BxRV65DvhNH1psJHR2EAvPKkOeXn08crkBTj6IDAkM1TQK9+hGTk+vf4gPqYMNnfqj0Rug+nkem
YOPGvU17jfmjBnACObFeDT6AqCME7npmDeRzBOfxv6sdM2Y0adourkBR8f8ESBMs4RtEVwuOqUAI
fvI9BjflF/VXZHLA0ArlP9dJ013y6uy1SfbIG8yxvgeuLZUHmXO6Bp1XAV7pNU7QOeuF/6/Tqync
6CLK/zlmTdQavax+effEm23Zs4sX8eQhAmyvZEBklJAYY2YigvLpYj6kbip7CXqfc6drInpOtBSI
MpUoGKU0gN/pNUVtraPOWpEFvojvuXwawFe1bzNRrqZPpZD65nQylbivzg+EM3F7hg/p8uV/AnvD
QNCvNxQJBZzLQnhiVIW8loJbL1bPv6UIuEfS/nZmU9vtaud4KN3XbmjnGxUFII9DkRoI37ZqlfAY
HSnK0qDD6/nA0RTFG95gqtFHHJLV5rGslrOTrM2dwnMXoaivwh4I9XLQSY51oqqrtFJt04DW//2n
a2G83gf2f7g0WHSQnMkIfNLQZAdH9iwjTUuhJyEdbSnOspL4MZ3azAw8hHkTjdV9ox6tzExEmLqk
KfZpBz4RnmbgaF6zU+sRKcFXggfohsUHS0RgOyUDl2Tfguy+J/bZ/wlP63mmQqhnRFObKinq4Gbu
FSH+AUiwszfzZGJaJ6fB0C3kpuH/mzKHS08+2tZ8/SLNDVF7+2IlQnBU0Hkzldc/07Ib5bvcSqCM
1a3xSbnfH/qVb1mkPIe+lf6ifD0xDsToAfl/N7Ux70MaVyU5uMFm8A1Bmb69tzRDoFsQh6nPj5Wn
TV6oAl4A+Oh/L1NKiqBjHBo+HWwn3j4WHZdWEo2qsVq3oVFb6ZOqd0MjphRYACaYrNZSWy+4IPVR
94H8GRMpzQ73dKEbiIbJFhWaqHim5PcPntlFwqxPBzAZTOYyH0E/IH8JduBzp/rKboz3SQNWXREC
5Z54/tPmuJbIk/8+/v2P60cVZDhCDvVoRWl471EwcHo/XxN8iGATpF6h1UdLWgSLH3TWYHC/KZpw
0Sxmr6eA+DT83O6ZrBqax4sPy5ALibLl1osc7NPdjbjBXn5PKyayA/ZLKHX1HLvAZnF1yiLjvAc/
wnFXO4AxI9qQMdFZyrQ2ny0z5ZIonDvkNAOyl2tm/SnkLIZw9ZXC/bbxHcnpKy0j5oNDr/Mav8D9
WB4rxRDVzcfbrsraVhG0BSUmweRxPxVKg6932SGkJzR/Uk1Tuxw7ffWvgzblZMdzNp86ZxESPA8I
oBgeCWUPU50HUt1dx3km0SF5KN/6ebmi9vQYDoAJ03V++EwPt5anfRu0A7Nnpwk0WzVR3/UVJ8z7
8r0TLA9hj11lwRldBqRK7Pza29PrmzH2kmFFRjHGbQOnXmYj+CFZMItk/OCZKdf+2pM/a7RXY4Jf
FdBcHKbEk5bu3WD28OonbZdyTTkNWvI61Gp5Mv3oYNUsSXwb67FFQB2g8I4DUPujZk1bH7ETP9DO
mlKdJUj2g16arpQDtqc7vCoZ9CWUyh6PyjN0oa4FpxqUbsr8hoBeegaKlWGfPAnE9KGImzLutAPo
IlWySx+MK93a+MzVrD6lqWTxuQxkcMVdZDY+DQ3SvkjueKpsYITfFI/wmZhMGwJSDb+eK9P9BzrF
R2rG+7AMtUelI+JzPMQTuIPfWqmE5J3kK7SuAjWVzqiTdJWfV3kSuGZznU6X9urGvJdpu3bauh8/
Fu4Ty9DGQopAOqMfLU9fJlhn+HtxuQuzU27uJIOa6q62FhkZDplmGgRDloS/MhVbAgulK0PXqx8u
Zr1fTtv4ldffz1x/dTzBX/a9XbU1KJ03gypmiMf8EUnMz5PcA6pLCpMSe1SCEDtJSne8OQE/a2ae
pVCWnhbSnh5EMI70jKEmqTGC3isMDPxJps6owRRco+qYne8XPqtZbG7NA/w4epc8XSubtUt3UEXD
gbDE6rWkVK2fp2KpArNg97aHibMPQvn/D19NFs1GyB9Ets5qq2fYks+YF/6N2nGlc6Q9VkTh5Y6Z
qvNShv7d5KxDWd9Uh64nGvIsukQ0wo8cnZx5uldO6AcwUeeA6JPHLUCjfBJxeJ+357navN/TUNjT
+FxhP6wLsPi3WFQO5dYWWa9sPzBdbtUjGFtNIXXkiXGzrBAtBnDBAvbmon/kRl+bDGx63eh08G50
NupZEBNus44uupXEl+yys19nFHDLnk7Hse1QjLJu1MlnJoy2xhe/lIHdxleZUytsOk7kliuapYk9
t4R54TCx11wncSghgkW+NeAmiLCB/V3E+QmsrxxGRXL0t3BBs5RvvI57ueh+ZVmkKq4T/X0LTL1h
FNMDKM7UVHidmhNVxzazbTNyVVkEbx0uqrvPDfh8sCuGLao80WPQ2GAUF1CccIkcnDNFj/UFUKcg
OBhMqt4Wt7hgM0+ZeHlfporF8+oR7aouTfC2k5643yIlL5FymlbGk0EwfWL09grq8EQA9YlBhfyY
iz/PHibhajgTxW25OFuhZGt969rb0we384vcdipdTfJ0UHGf4rn7ekEzV3XGySzqN2nwZgZkwqWL
veyW5tPGX8eNay2uJx+EiPdxZ2x4HHhzAgbwxa/mdq/iIb5QhAOBU+eICzS9666Gc3wzkCG1mLDu
ZW6EraBs+V3mIM3nKvkaQemUf5zrkgMTEjtbdq5NivOqFZCXUSAcNOgq1yLnw0nC8HW67+nKKvz5
kGNWmMfx16Z51nJqt+b1ucidvz9EAy/f6KSUOwZ+2qCoA/H4JGnl/gaF3bnuCrchnsQaDTSdM5Ee
wdoWhhAorjwb5fNi3ktMmPG9AcK4KVNUyjPOoMEEot4BhJtFMUx9Emov/4klLZTHW/SGuWxgFdw6
cjZL31Hfp5PPd3PQZlElTHn9LYR9mq+cPiBmPPIpzgniqfBD1OPkmCIDjCoX7dgRuGOTVHorLxGu
7FDRwvZKCd/tuWTYVkMwJCLPNEsuvyq+vk4a3PG1bESPRX/CHWZw8/P35UjnnD4Ah4a2KRDTA+O+
2YeBa8u6/BXEKzqiiOLGk/xhDMyx4CZOjkeG5bW3wS53NbqB50TAgInUkEQBcZHYuabe+SDMXSyE
lDraUiU7ji8SigXy8XRM51VUmd5PTAzRlg/ajmfRdhsTRb1WFc0schak3khBByMiey3h9ntmWPj3
9+AlOg0HW75kjT7KyPteqWnK0K581lNQFcIi0VNyXjkLbsKL8tScKITRoQyWqWON9ApJ4WdEeJMj
yngAXnq9/RfCW5Cegul0BGycn0f0mHeOftKFGbwLZPsk6c3fXDL4W4lE6qweJzMU7FvpaY78fA9i
HvNq5U4R1XvxIK5Muma0re96IzkXxCNHKwnYDrlOyBBYWZYhxKiyXtv83PEUcFXiu12VQlCzAXPC
u4hwH0LBeRc0bJqlfeNdRsB2cAQkOKHwMGqhwI31fkUH88poTSruaqMTz4MDQg0P60kGBeuYrY5x
2ScTVAjfvb92IUjdE72vBG7orW8Sz9ixmgvLtKTaKB0EQgevu0/WmVU5OBYbf9NNYsVRWFgib0rn
QMuFCz2rEj1dG80wIYLa2OIh65/saazPGTmkQRU5WSROlWBx/7yK8fkJ1Y9zeW3dltUI40cy5TSN
nsaeMwc7hLWSEEdE7sEp7v/ghc4K1NkGmqOPcx2XNYJ+mrPtCZ/3+TUW9OGHycZI0rFFSyNVujwU
rcWLYr//8YUbxRHloDGDntkMmbyukL9ZfbkslOnyy68P/RuUND4lJ9zffMdcJjTnzY6xbT3ANFaS
ys8ZxBIpd4P+r+g7nmQRyX0kZx7PXksyJCyplW2m0GveDXYexy6d5Ui36PKsLqsV0h9uqu6cCpv8
fCCAAVhJT9K1bLHmsPhua2g5aFw8lvVwsf3+2YvFVMs2pU7Vo2bAcoTT7cOCXneoM+90IMejBKRe
aKN7yoj4cz88K/VOQO8yGXmlB72FmSMnwY2suxUZ2G5VdWpJfK0/aUGpt3OqWDkLO/Mw3VGW8Non
0CROv3j/dfuhbH2Hln7lyIELHCOmYXfwLEkXV42HKrmVJWUE7+NESOxVex5mRxL0SFXs+2VbNsZx
kTgC02px/Cz+8/7ZdefL1ZLMiATkLNmoBM/oZf2DmgYHqijiqxZ9CSihFsJwO2HM/RtqBZdD54VG
VINuW5vTl9BGPuNfElIMKKkt6+wB0z4M8cIQX7uJq2JMfuxtTnndjY3BI5HLo1XjBIu8WxN++cqT
GXdt/0KD4ImJ2eiJ8/YAzNlnZ5tJVkx0jl0WHdd0VHEAME2q+3xD5pWB8DE1Sz6uf+eX/sBU8I/y
FJISPh6ohu8cNFHTaG8qpaU3YOeIiCcrZts1EWuVlG3t9NWN9+C2n7mkxhTUJlJuBCkHe/JQTw7d
cXykmj6XOAqttn9BbqQcPW5Yl5jQbjTu9WN8dXLmKXsoshmsMsWwv7360WEWCxYc4qdqbIlkzi34
4x4LDIKqrwoSL3a8ImI9DG9GSHNFW/gXe0PKcn3QptCQyp+LGEAqP2weMWKYJxex468R6QYb9Jh+
mj+iv9YKEG/m8bB1IhDvXh7BGLuygbebrBWUctMnHTChmhub9ReroD96NXWqJ1qProYj9XYmncNM
+T9IeIj9i3ThNHr7LDuWs0+tx5hmEB23wO1e7fC6624+uktWF0A1nN6tDxsa4is0KXstNV+ZkHx3
NiJmTV3jaHe5ycMVQoy41QFTVb6Lle5UjChyukK7/LI3RqRgX6H5e6+OwJg44nb9netaSKstijIL
Rl17nCyFlnxMphtwXSM9z2PhMz9ClPWPCdptvznPuNZZfJ0NJdQJuCL8+mNi3RKZzMK/9i4xL/pi
q+B4Yh6SEVTyX7iewjIgmOImORgC0HXJOrCSfYo1chFRB+ab5VN/TT7FRcga2iOOjoUoYt7WZgE3
CTV0oOG1cDtzq3vxzl7DYAKiE61+8uD+BxxeQcqb2KsrEHf3fqRUDnlFs06Izu/80Q5Qa9+xP1Iv
g6J8QCKQLGhbk66l7dYyj/w5Tjpp8L0vPipTvGVuHpqBUVWyPDuGLJ2Fk/m2w1Q9ywYBM0WbmMz6
PxPyky4HylCGJQZPFGely9Jrw99+6wF3ALlkOM/pfAO4ouUt4pj6qBmYcQtR4ehCK0lPTYHr/mZx
ErFnbfx6C8ueRR0NsFFBlid3ocH/wjMMOHfkX4cfTxaeLaLZfM4ZkOtGL2mwmRofoWl+IAdLXPyb
HcoCMyBkN9Enykv4yo/WdYGQl1o65znbJU6RA0ZhePvlWRf+KPLyfERdMn3mmuPS2rjbGqYMDMTj
xj6Ro8QHwQQ1ovgPeonu1k9Ydp04tpjziYPfArhA7dV+C1AtdVHcWK0LVwhObPExdFxpwT8/3Eh3
I07TZxfPfEX8eH7JKf9LOabC92JKPiQs5zuzER4nW72I8RwhzYhuDdYnpUuaftI+5IvwYCKuhB6B
yX0hKNclbTGI0DmIgUfoLCBOp+Vn9gz1TexFfWa0LXp87fuQoYXDFcRlVXmhzIKaJMj87cc2FQ4l
sIlhMxLJWD/FpC4jGalh5XvzlBOFCzyjyiJYdJPEnXST+XQzbXDqbUPjSucv19hK0y0qkxdn0Spp
AUcGOyMLu9XT6uN9xmLLe59nqQ2ywbQhjx8I5ZnUYgNE6rNNOCU4FjiwTHEtytcEkIYbPYQ84yhI
mwFUiFkY3dEe15DDdsYavJQVWrs+Xd3EkuOuhZtDTbFNITvo4EuMgLL59huvVAujoq1QoDnC13XU
6SK+8XRleZ/f9niwV1QCnq6IIRw/8RiSvaGm9TTgEFdQvqvXzp36X5PfEcvLs+pZPy2yFRq8c3vM
lR/fXdcHy8pIe5T9SPQnU30XDB0aVOBtBY5HDesXZX2k6WW/B8eXfbbMWnMQ7cqw+LwJLOwBAUDt
c9rE65Y4+b93nH6AV8HTdKFiLTfHwVpx+zLcAsRJIT6K6SiKEM02OVO573vtghvCPRHA8eHwjfjC
mcl2FHa8GMx4zNDrx21v8PtCWR5QrIxawrcZg7VbeCBoSodEd/sV8wqiWWBP/Qw7XU0E1maZTJIf
+yVpO7bjWmfSE27P1eKS+rJ1DO2eq8SFqK4lhZryaRB+I8FKrDE31LcxoCdkhyTZXmEvGMwIvXht
5/6pfYJBCUa0kOHiguImRlimQnYu9R6mCdg0ydiY0ujEmnC3tYElqwNypdIoX+TGLAJp5Ig7Ev8h
C6ueH7eXKDFxfOticD39FpaXsC+TUGBR90U6ea34dR2OeTE77//sSE8c+0qtM1ZfXyQNUCS8Rx5a
+b1rxCWsDzkooK52a+8mV7PP/xyx96hSlVy9/82YmzWPWdxBwpv9w3qhO8GntgizygzDVF+2v04X
bt4ZeAF3RCDjDd0I7Eqfpqh4ebGgPgM5g+v3Yxky9XOftIYtP4RFfxVx4QFmYbrdPwM5pxi5PnFt
sUHW1VIITIb0a8ks5ybv02gWlsb6kacE7Ui35caCSmdq4a/SD3ATSTbbiiNyIZBruB5lYYzjQ4HT
Jf7D/ALSCGNwjt3P7j556nzxutglwp+KULp8EAFdwTlbHMnZMmTblcqQSVcwagYobFNCAxO/1gfY
GHoSqVzN2LV81MrI/TsbXFvisvTllHW6KHi3x0d4NVO2+Zfcw6D4EnLjFetU6AhXJVfth73ND0r6
Tcm6So/AVQkkuw7e6WeCUIGcSQeuRne5OGps9oA+0dLdLqKCWOKIBb5vF42l+i/MQsszu258mzZt
KOtgiEri9a7Vrw/BSOivK2La0VfvndTbnhQtxmJmYwqngL15NVednv4rPnODS0CI30yXdeNf9xT5
IWCu+67FKH2z16sbxu+LH3WvBomCbdV0/66T0LzyQHWbVHACdFJ06wCcGeuBraZAVjT0uuOPUmVC
bmZejtyLF7f+5DbSc8EjAdJVf3mubWfbvS1HPyYu/L3A+rtDlrTBZEhNqOz+UPYqhZvvFyWx09Zz
bmY84U4MEBpm/vWL1AXu1Rgcl+hJ1EfIoNa6LBQIUpToyUwF8pw6PBGf4qtL1CCM/C8TZTzTXDFV
dGczNnsNkRqIvwWWHKj5fFfB3o66T1ZwoZtLemamPD1MegdcXpj8oHUpkEDoD8ojZ0PWzQOE5ICj
v2/ltTwsyuQsbnbIaARq3UktjMvmVsvnPk18UKafwg9g61Xamw/30X8zjmMytIjzaP2Qma5A5Icq
qX2eVWiDi2cfuC09zDQv0jFVxSnSSryG2GnJrqGu7bhxLPepZySZ9SbHi6BwIHYR9SEamBbS+eGa
TJC8iIMeBbqRz51OdiVAm56zwdf0XK5T8Hj+5E2qIYo3xMp3mOnESxB/sjJulSVbYmCrjbiw06nr
kVF8AmLA0BsechRURck0csRO+cR99AsqyPC2KM4Te/oXvU1F2TwHPnqdU06dh15XWuUZmjBHm43R
mk18N9z88xY82hVrWC5RWuw4GA/Vn//CCFgaE9639eCnPR8hifDRpbh/BMn5xVFNooyoGy0qLteJ
DjLU64r0enBa+JYmJije3Mx1lBbdw8YwZsLSQ+1ooDo/Q0jpyjUOTXZmk98LHrqF+uK1A38MT50J
8SGBBlehcoLnQu4ROZA1lUO02Am6/d5CkUA/dryZZy8pELVzvn3EtxmigLH9v4Qv2lmSnE7rJiHP
PDuFhewMJg4usJ02qwWEna8cmf5YTVt9jADT4hE4b0P/iEtvoB72rvc1kTlt/HrhWtDbD+/5qL/4
5NRMR761BRFjBkmC7omJtSz0mR1kRPvYbAvE5n6C5TuVW35Xt5Pps4isE6rRmn/xo8SeQNy4ukeO
J4Om16bq+G7tZaWpSM5E8x0mGoiPUnHQ8lZ5+95meqGMzEB1kTJm/FJbaJkxr1afIaav0ZXIiVEA
+ta0n0+UyjFNLmUWLC5N8d1h3Tt5DgkCKDtU848gK0rKegVErHzh1q8wZEETgFB+zX/+voDD0a8K
4/Er/bfVl33OZAhzAQZFFAK5OYlDEUCJiGDcFAZ7m1YS6x7w/VaF7bdtlSSEQDGlDayizX4VW/1H
NS1kkNK6fpDARyOFBIqUiI4XDWdQbn2qokZPrwXnTeYvCgUEzCJzOonPg6xJ9hF8VmS31M6GBQab
/ywJmOCoQJ+xN+D0BYSEqZy4Lvx8d1AxKzvG+LWwbM1rJGGiidXpveW2gsZNUcgheP2zKKnD6RGN
LdZTVVI/54mwBc1xWYulqyf0ts4xeUVYetjiZuLM9pHo/dvXTvRs3WN12sU6PDP1jdPQGkXbRC4Z
JpKEFfT9J/fIye9C7DtIvYAEI2V1vfgcCVbCVhyzBVz0TP+pjSvGC8zEpVQDKIh3wiJo+yhZU6S0
tibQuBekrpUhG2Cx60jlEquufwCq4bV3JLcGDLKS6FhNQ93BYGjTVRaOtw4GFAlCrP1Psz+7o2J9
XxF4NieKAFT7dxZrt7+u40zjUAml1RXWOhGhTJT1WQ1ojihUTbJqyit4U8ckX3z395+jEdOIBN8h
40q4+DzYjcx9yPV0N9klIQI/6UhSsqNeenZHc3EwAFix54wIhSjS1dVNFOu936x96Sm2WJXBbwr5
iI2nx77To9jzxca2KASBpEzOAb7CufPZU3ceeYquis7lqWpBmYKCvLJ+TFtprTclcwFoLeECke+c
Le6Bv482ZUDA0D4zbL0H0MU2nCQ3g9eOfGOdfW5p8gfdX6kj7eK1bmwKWVJQNkwsg4XV4RzF0uee
etcLXQggcx2rz0SlfpPrJD6e+c0wZpljxlv6DVh3ozVY51HhsVKBZ8rnTJv4iY/UWwXcrhO1VSg3
8LrOhu9TgwXWgBKPg0tU1QGx9CNLOj31ShirBT23d7dJCuhLyW359vQQNidCm2nRzKb91kj2+MqR
AEKZ7wQYHag+Ogtqm4iWDwyVXTXVQmCzXybtfX4q9xpOzykp9SqBOHpjzwzJ5xXJyTL6kDo8aUY2
NgkTzHLkXtSV3wKdumLxgcfOgnkZGObmP0qP63dsYO3SK7DypPgZXQN8sAmQdTh7bibbzpxslAI4
JbMT0NJbMYv0KxQqaduTITHK1ozKhc9qBW7UQB2tTUd/iS8N0xGgSnqIcP6oNXVpIbB9PpabK+r2
A6noXNagi+/MgtEJFZoFKkR9KJOXdyNWMM3o/z17wmJVsaMOMjyDJwby1Y4ETOX4P1jbI/sxjQGC
KYHuN+LyAehhsv5JcHFLa/Ni5gkq+kItenmxPYOftY4DryfW+GAD2zMcseNRlTcSmFLKDSJCELve
l+9kj/6bkxoojc3a/y1jeodtUBiS4qyZ/5OKJT4BSL/+JwqVjCEWaYj4YySsBokyT0anxkERscAz
wXt+HQV9EGh1eWJVxLJta0/8tYSZjmgREva9gRIUEyPeBjw0A2xl69fHc451UIptYNKe6w7kKHjx
g/MPpOtWjw+yeTsbqXUanVr1vqj0TBDWgEkj3g7B1EG0Xl8Gel56obyQMkdsQv+u2AlgmE+MP37V
nZnfRLspuVReWX5Gba6Fn838deEX9PDc4q+BKBmPXRG8Wo2Z4UfMGKcpjGdLm3gSvHQc4fQGxvFP
PDWd7WmoPR129ehAeXN5fxpQ2RAD3MQwoIUn8Gs/KHhQaY7HEV1TmY4Ta531DZ6I5OXYpYb6114c
HAYMcmtDqjDNrowbmNwOwVo0gsRHR5iZmmSDOgpcdTH1XUI4VvPHyBoJ5o0QOz73W/DQanVVA1Jz
JmvdXLMIIXmyHyoYtkvYXUxWHyyZoXzH5lSPexHTKoeX43KZmwaY5NXS4bG0DkTuzlKjQiDEqyTv
iFc0YgLo8A07/REPq1rM87UEUTYk/vHBMcNSlnpbqvk7mJixRu/lWQKfs8w0sAJCQGEtoQpE8bAj
qbDJtdxYdGlf8zGu7qoXW7YiuWbf4Wro2FyRDCAi7N/riMKa226Uxyx55JLSitcoCKqPf+2/e+fx
WuMeSH1yfUpiaaoHakETdjNho6PlemjulzQ04pQ9a6w/gPr4WF8U/miMpiLsvja7fYoJIzV+nN4Y
K2CZ/NjfFFnlNE8AfksGeCwkwUy2etXKFyqs5/dLJiu8+JOVRNJLo39TKNmKQPU3umFCEccB6Sep
PkduBMNloFnOhDWKMi0VdJqEkl4LJUjcLlaHJxe45E4Zyo+Jf1GzZ2VMJm7SjF3qB4O0tzcmqsaG
g+74OheYZVrNAqz81c4v/rpk3zDNQmDrSetZL+lBtbw0SBkcad1/TaZJIlib31a/gW6jmSGv4O7H
2fJoVYlOiiFeb2se+x9pRZntsD748ZkyU5sGsfCalIeSP7ddoCHe4TD8CPaIm0qbTtkfufD1Jyzn
khJe77xPe6Va83VrdOAnR+uMZn2UTeCBL2v3PwIMG5NtlmvFJ21Wm67IJ4karrmZRpLfgQSKEPDh
6bQ6re+vELRnhV942sP5qQGN5yAv0YFrD2sx/9YC+Jrs5BHrjD4rJ8YG2cLeQCetuTPHqmrrIiqB
V3sae59w7PCLE/ehnnOJQCRkuAD1a3CcQtMdtsddKa/s1cTLR0aoVr2s7WCqKLJvlPpX9Z+wFxQp
aXQEVUGvahjmZcNlFzwF8hxMskcRwQG8aWG9f+Hz4UsNcNlfGd4urO7Xtml/NqgPHHRZUnhtyjTl
U2B351qaSQb95+Abdnaemn3DXbGPGiPBmbN6f8kwl0RT/hYXPh8iIaDGm/FOZ9LkQhoiTLOOU8n7
1+wbsR9afZvbIHCZ8ZaS7uinaG5gw3lLT2tcGEv7Cm36tygBAHX6iJkkVN3lFAf6gMgaMV2o1YGM
uWH7qrtMRSBde66lg1MTDEvFqlrKOQMd1tawOcl/OMDIz/zw1Up1nkhfBg86B4KtSjSpOUPgo+AZ
g+fbueYw0DfXHMUiO1t+F4qd+/VnRRqK5TObJgdN09x0DcfnVwZApCvAC65BhEqgqueHQ6+pDoVS
jXtMJdVyF5PxBVZw9iDboUGPM5G6xCjDfQbp/W3mug1wtb/DAqJA6qws93Wevi+kBiSHZVdArE4Z
7dEU+ManEZen5MbjBJgTI/jiMKa3Pyc0k/svNZuaKvn2ovNHbZg0EnOSpbU2wO+sUMWpNK6JsDdB
oKdhZa17fAN3L9B+1fdixuogGsGwKAH9ayYmgSykOhHwJ9iO5yrG764Ya78UYk/jjf2QhrmA4lYQ
W2oR3jNcVcdQNs4idg5K7jcSxwRz+VWZxpNXbhC223/Ontum7K1cVmYQSOi6Ck0VgT0sjtGheZNV
ksbDS+k2gL+8uk0/K+mcuOa24KBmftcnbWKbtsXCoB2U9p4BYVVXWapMizwLwBNAZ9nxNCqmWxIH
EOUM78tv5g0dOSIWT4FOn+CGEKXcaZdoDoKZYhFt8CB9rNWX0gUSfnepOY820sFq5ABjEOEjh3R0
GhSjlZKMkNJC8/tfFRGa1MkPm486XISkvjgMhDHFhaNm23DKop2au0C1pJQ+lMFS2V6Nc0JduS9e
NnQ5+QTRx7jcDoiu2zo7YUwGivCmBFF7cc5lrhmvn3zMdePzczMFOmgkK7b4EUpyJy4kQArFHAtn
OYG59/451ES/RhUZACqx/yAeH2eXreiQf9FDHnsGBnr2qTzQPPbd0Y2Yh/zr0Zee2qMKNE24cNmJ
RZEMTcszpMnINRa2z5OmqeR7kv05Ooy+KE/sxQ5aZh5GZIo6jF+DwhrByxg92To0yM7S+xeTPJK6
E+P+NZQ6B5Z/fa8zCMJmWe3335qfYjNGuOOMP1pFxeO7UsctV+xgA1fnhIUYKyaFflcxrCvphGBh
gHWhj3rJzm3WcICOyzdWKCy3EO3XTfcSwQM+bvfEcDf1mxFmI+Y8sgkLCJTJd8luiphxSsUOXVPx
I5x/MXWIXfrO+xVfdG6xdeAoycPm8MWaQaeoe9GTE2XC2BOLNlx9olpblqoz7yMQiCcGshMQsWw6
3EK4mpXKguomojpKhpDPtCVobMV3HeViOk4t34CehX2d4QvumHTG/aJ5ceUw40uRQTxhBvSFyyIu
jScjgywoV1NRm+NG/gbCokhr/bnFsJwIoBqqVc4AeMdR8G26/9FzzaM2dM6oQzRFyGUa+oVzVdpm
tbpyn4iz1QC/bCrk5x/1A3DnYFPyVatOOqG1qL76lDn+BJM+GzRyFjWr0+x59n0nzzv4alqqvYrj
3Xpw5llDcMWkSFGUIU+b7vD/k0evo/0uk1qTa/y3tzf2QVjz1bJKj4Q9AOcwZbR7x+6TzFsmo9qS
nIm4L58Q9dG46nw6iwfVqXSgay6o+nJx4m8fVQk8Mdk9/ABlJ02FUP+OTS0JaJJdtWDDzIoRbRiS
QjJVrJO9a6DU3EFdXrWzn52mvgEl2SH1uCyz/Y0NTuMf1MZ3hCGaZztznua5Lds4M37KoSa9+aVX
h/0CWR89ztvwZsMtb7+f5j2o62YJEL11Wv+d1m5lptx2n4WZNh9fU0Tn45zAevTNa2YnsbMz73nw
ph/lAl7xITI24pUS2xXBhq1c8gKoDac21gXk0K9llMbY3J8z0vK73+d5Vq1J3MqZ7DxUCZqXlGWr
3wNbVk8NfJXgTch9K1Aqw9/qCEcHCxElsZa6TzIaYIdhLOttc0SaJJ+KSAbiHXmln7oMZLN7SC5G
frI8AJjPbnS7dOB76oDp1Cu5mRqQYzlT7E/t7ew1IiahXx8O1ABCyoRgtgaWrUzVHfu8BDIR4XdH
oOwi/3qV3KIZHv8HT4LLyqQKt0jStEnfGZWKlaScu/Tk+6PPjAVz21BN/kRam3rZdHlNe2jtW9Tp
DbxOZo9GyTQcm2EUycvI1yxgmobsInP7ZWiEAjIuvXXQfFKI/o4RHFb9yAGCGJx7bofn8Ehfc6Ua
oiAip40PhNcQxu5vdhcM4u7gd44dE3oAQI2gZwcaW/YdqSkeeRUII+OyenS2+kBN4XpAUcbrCRcP
EoMvGpKUc0sK7E9hPldOG2CSo/km9wsc7OU1BDWARbbzQAafF6M5xWxBzywiFXZf1BURq2M7EWt5
7TM424X1V1fa+X/p1DJdBA5O75T1I2F/W04E9l4mJIW7kcJMP3J4BkjBjFOtIHqXjTFFrn3laUlU
0BuT80IskIYC2Wv9KFPSEThhMhUNruQWCTntALa4e1f2a/DI0yQuLYY2W/WPzlsqmZOTVpkk4IE1
Veb11bWj2TW2J/VNSFDg78xrB00bPXZv4/VwHs+nYMF6uUMXRynLs6oXTmrI1IZEwAYd33ZruUsk
EM4dMgSo2DeuJaymuAbmNNUn8lpuxOdB5lmCGcCxTzXxzbjqBtfIggV1wbao9ehCtOJ2SGz60ZNY
JYM56GKvdSHSe+Ov5smQ1y9lq02cn2+NNvC94USsZ0LXEu1NP4g53Ng0BBJh+nAAfEnuC4WeYtrT
oC3pq8eH3UebCpq51Mu4AOX5O6czV0G6wf1MUREyB6Bl2n/EJz6zM0eUi3mE+H0LrNybmRVBGV1g
QKGhV52ZhFqo9CPWgeH+/kQ7Uu/j5zgAa5XqIUx003kYoDtXt8d1rOrjdFpag3eiL2YMkuvgNKDO
e92QrCJ2LsB2DKPIDvUx1EIbeSoOntHMtjaON0hg782+xLfTz8foDQEwrE0WbF2hY75l7tMMKdMp
uvTrCvV9GttQgeAgOW1con9jcCApJfkGFCsBPnrzrgM8TURG0bG+aGqPeb97T6S/5sqJSGNzF9G+
bJzvofTemHasK6Ha+KrA3ZifO8T3I0bTlu7ipEMRebEv3K4IKC+8sNzhQzbOH2QLe/FuuZVa+LRD
7L/KciGapz4c1dswnJDClpz0ngs/j6CtT1ejWORAFdHqELjCSFjMO4qQYhAB+EQF+IuSC8ieK52h
syzhhy5Eps8voAORDp+lu+6Yh8evl2PL0rRDqwYoMTTXpUQvZecneawdNb7hEaaGJzQHGhW/+KGP
Mn0sOWkpMUnoXPVVUDnycvRGaN9bPBDD5WLsyl9M6384NKk5W7CV2Afi689RL9xNAzroLqx0+d3y
RaWXLz8fV/H3HzdwzCpPvChcUdoVJBrjfY6qED4mZ/g54akNT9GnDWh3wc8LwGV6/PCj1Z3HFEpR
oDbE1XlVtQn89mAKJgHT9/krOU4R3RvAdJH/c1T710PbD+fT5gKK0LkSg4ye0wip2L78MQja5e0c
S8jIE0AkU6JlfUY+ckNC/agyj0jKiN9J+FwvWy882th/BMKP6ZFNgHxHMwAifMeiutdHyUIOjbzc
/Upv3awFDuW5LQSaF01y/a+5MP/N8qCBOduwYDtbvDGpsVI1690d+e7YfgZ7IaiDhaHY7at9WD3e
MekVeMoWChBLKm8AXwM13nM+nIGjl9380K5dyaq9AoCHLIE/4IsiZKK2vt/opnRuVFB3+OmBfSlT
4THR/WpKwDKf+qOFGV9gqRaCbtmXJZ6SJ2P0HI0z/GljulT1TSouEJOtVK5ivIkIZs1IdvJ7a4vK
Pm5CZkf3cI15VR5LH/ATyQoz5YQBYXX2K8B7Dd9rqE9MtcHlFyd3X3D/g0nLlWmj5XwAbVVXt5XR
drTqJ2iLcB5MjspRO7d6plonbjelfJMaGnacDKVGEHWmfRkmS8pp2mUIb9tTRpSKpYxulflMDgxO
Yyi29LJRexFAhhP3EFLQe3ojTcVwh8+UZ4aZ6Qww7ZDAN3NXlCd9hceb/aPCr5XARV0nVYiEODBp
0R21pxoD6Zo5FLTFWQjL9GwgTQZAGbQPkjIrFTNCRVBISJ+d23kNTYeFZI1AkBw0nU5XYxtNefb+
c3N8r9a+LstBxPpsZFZgu1J+qSztNDq8aoMTo1m7r1DbhLrIl3jx2835oFQEjXK5+XCF0PlOF1ED
M4/BRPP+XxLgi1vnx7ZzeUOVXT4QuJbltykMkdl8Fa3R3trduA7sE+nJPVBZMdW9aHc3grTJIuvB
WDNr+9AbdRUTPrR5Qj4u6MxABqLS8A3ny9RafaUpJW7fmxpKlxdhxHDFFceF2Gw4WTDCgw4+sSBS
j3ij87ZlEOEFlx3oRn2cF4hxy3pDGzaAgki6Ix25GFDfLGX9uX8OsRkRsLksBC2LxWguGvXxBfRa
fDgkGZ273QhGgOQ+TB83gwGA7hPZc26MqlVhmGmKPyTxAXYInzIOOhYoHt/gKGoJZP2F7QZXHkr3
t1TiaPgs0O1fsnTtAxmdg9rOFxcKDdjKC6pIpdwc4bX+9j9B9iyjz3lW+lGqAhmMby9sHuijW4Pm
aaNyTR+BjXi7FVeUibiMrAC/isUfoRcRTgXYRQNiYPj9snaJZBayYYxbyIKN5xQDXgkJomlBaBrN
qfG1B6yChlDVBCJGpyovY+GVDsDz3z1qIDvLErbLSMer9trqvWZYiYz2T94befh1HOiObrM6Sxi3
N96Zq5Imo9ABHLSOJ7r8ITKpSIvWTlBuyNF7KqbMhKUztBb3PhQ4ygfAUb1GuUYkPxIbH6Uu0Rod
obFtX5H+Zdt3LvqFewzjvtczhftE4tHA7PZ8Iq1KhJdgsr6FS8AXp/K+6wTEtE6ddEeE+oUjCzNj
0G7GlcKVuk2xOpKYHN2SgaE8O2sHUX8Ckx6JDIu/rxSOS6l8Y7tSLKIo+bYCLcpl1Bk1h+2FHDW7
aMBROO2cetrgPk8hmVBOZ8SNgPZjIOoVlZAY0iwBN3zzLoDAmdLSVWRpvyoDlSzwPOgrRi+/rAL/
xNftjElzuEgxv+EXmHzcmeRJZ1R+a97M+EtPtzV2yMXiP+uM3ypWDay8X8xJ1X0jIYP+QmyfWOxm
20zqhPWoRX5YuM7C+SfKhjPsc+qJeoClge6Zx6H+yY76e1wUAnz3ZnghzmWm8UrGQlhPsCRe+XWg
Va2/BqRyLKDGWwcqNgV+bh812X7+Ws7GHE1NM+X7x5OB82xQ4MB6Z3IxAoOg/1sRpfL6Cu+c1nlU
1sWB/z33uf3cjeW08CIQ3Bg7Ca9YphAhY4sK87wSrVBomC5E0eEC7AseH9tRkJQaE2wDB+vP4w3g
NktKa1b/mhMcK3bqNVIucnYscQbyK6rm+n4vaXbuuPumsY+9XBXsrxzESmud/33bE9SDeCaE4O3H
+gNIjB/d+SaIVfcWbrdVMOeQ38KrmWS6IyFkT+sq9YqkBzADMfuqEclph6x93zCNbr1Oo0f0pdGA
wQ3bBAOq/eWebrmaOpLZqoGp7M0+It8+Cwv0SpXFIZVwFXynBp3JyVO7VlRvzTCuyJFNquT/20sb
vuGDklk3T/xHAdDFx5e1U3wap5buj9xSdsfeGOSFfYnOxMI/cTAt5PLUnD2ywk0LjITCenCVIHs9
vW3CvxKTzpcKBmTQGnIHJSsBBTtKdOp2c2fuMBoqCGMPQ3Wq7NKmUi35ent5n4LQRM6JbNs24ZKj
jhmjvvkjcieotlBRIFwMv2qwamnixac+dqRf1x79MKnx8V7lrxQt3/vBhkJ5Z/oLLNKfGpX67wQS
8mWqxvm6RELnMbGej/bKUlPR9lnZk4pVyjn41kOm+ZYfdHHy44wdF2NbU/hsZua4FgN1BZrDQVfE
pTZqFapqiXbCbKbCPqkn63QtioB474eP2tJyKWkfJVlEaZNxbHuMzhVo6mzyW0YF9r3ty6Ofnp6u
xvTm2dLAeoSiEA+kOuk2LyShEsHvTVCwWS2iYYN7gJ3g7lbDjL6JZDCR7qgf9jDPKz8sHHlZP+jM
SxiBymmMmcLpoR+FZQe7TCI0phhMG+r5NwVPvfcwCWOo/7D9rg8+Vjn2AZHW7C50lBDl9PNAP8uD
hO2yP/MsPQZdOge9ftrGq1xQIHFoVwfzBybEtmEp6TK2dMhnZNKaPxKZgzTyC4T2b/WZNlbJ2fZt
EAEdnnfun7+Obg4wwhUp88TM+GcMP/clGOiC3uVQ1ZqIy/3kHhoSxV6uLnagwULUUhlsygIvht3J
qKJrJoUB4A5LF2qGtPWmxGxoN7ufRm/qNoAVIOxb44bMBZAyyTGs+CIkrBV6gJUgSUX9cizPiSKE
PmFA5xKhHenyscoOj99kW3ptbDY9ui9muwozEoPtAXwb1RpTcDXf229AINnFrwwB90mIG18z6VHS
Xe5W5VN7T1i1Ssd6BWlLOSL67JvDmPwUkmK8bbdFKtcgAcHd1IdCg7Fm+mAMu+rDH1n34sMCwQ5+
x7R4qAF+ET/Ytn+t6gJUUKMx54jS+qYZxXMxbfk4BrtBqwm0f/cKEk2LlClUQXUjab/nE0/Af5HR
R50a5tDrE44nn9B9ibP/atX68wwpvpM0+C32/y1RXLsYE2xNayiN3/Oz1C5A04cZ8UVcyfy/sgdA
LYMGU1MWEU2JmX4o2/xH6GVFU5L6+SIVt8z0R1ieHF8XKxmLy1zD4RPS86Cr6jfkj8RGEDAQkhJl
00/jRg3C8KAEGv+7ZBWwVnNNuoZ4dM+Pd6s5teBma46CBARn1wyUaxqOswfeIsxkYsIdkMvIhTUM
bAHCGpf2GUN1+vJJQPlT1QB0nSUeORbfWdOZdaBz3ruTcEWUaqEVBuO4ajL02EW+iJVzcs2SJSo3
lHbzZtvKfydFPNNmPqB844PDQREYNhQTMFiOyAaJ4acTnSMGEIXp5/IO4ATrRJY5drcj7lK9XenO
Jsdu4/b672NJpn0vuYsxwht9QJNrC/FvbKXMyjqELsME66r9nq7C5aylQyYgqo1xV4ARKpkEL9XU
SiWWc1exROyM3qZpQ420x4YBx3zQNrIuB5zg7+sqe20GP/LWzcMZMXerW6g0JIyNEWjKgIS4bLFc
Kiq+hw7LWov2+LnpMKdQz9e6EcW5ix7w1S5Tm8packdjku0VG7FKd9YJCPw/w0Os7gikzu7/i96+
VojvAn/rBLkTlanrUUBV/klp30xa+6vX94RA60WBCvA1nDb6xSTYdieZhjgZqWCQF6Gud+KBvPK+
ZM2nV5SrSt+6pcx+BqFIM8MgIkAMmXIo0Db6Y87/T/bawyT+Gx9Sx/N58Mff3CmBxAvpyAo5WIxe
NWcA/9Oql5kE2TReoRTAl6gK5Rm4/TxAe2yw9H4BYDekTC7z/ypsAmDunaSJNZKqIstBgZYrENUy
/ZRdysmskDQkIViwh5TB6MGO2sVajbZxDlvhkuRncv7PCMrr1PBxmUJmwD2tuW7I7xkCMpn68Kh/
lydtbjuzwEdf1UH8KU0+SJFspUyjcygwuQfvkUuBtGagweceKJPKYhu+cQ3Ro8KtzwGdX1HsNR5Q
vnJuBgL7K/kD6AN+rh9NYCNH9ZcMe7oc6UE1CCU0cH3X0bbNSROf9PP1CyVT+WRCc21lHgeXvDKC
tePKqjmKxmxf+TN799GOgH8OD/M8x+qWu3uG0ahukFvSYVP6AOIQjv2LItpDjRwtEl2SjublDVqR
992QLB6WjDijVkVYSz6SU9KCQD+hyjuS0+IihnzcudAdm/duWjkMPDy52JjguoM9CKnCD/NVwnPh
tM2/AfnO0uyC6ZKNWDBzm5xx7aMFR/UWWyE1MphxiRBXSno3pEH12E96YdjHX9VsH1Z29SnZ+XWQ
7wpcvfmC/nQrv3CRQm/j0bI5Mia5iZPX4QtTjXR5cr6OF/I9In+jFg8Q2gqtRyCqfhva1Pc/fhaN
A2wkopseKutgaXHuvxWXOHM2KZA2t2H3efoFrwPgvkHnp5Cf4FG+kghecVc+Yu7EbgUHncjcJA8e
dYU+dNZLvUzIuY74pqhLr6I2Tw4Gp8iofzTpbsXUW7J5y1NKfD1sbRheM41AWeC19zUvAAbRiaZp
EHFjemwAN8BXBgwTebLN27GUs/FwUPJkaADCWtB3+sIjseXv3JWsvD1iJCudPGeyKwhb1g+fLjej
vd+rZkw97iFtMq+/E8xpXBGxRa998sxHDYx8eIQHQTvc8g3GJt6Ofqt1Hg+9XMtj+kanW9ukETzY
kdvgnpflqwmOrxA3Tfsj0rQmbJ1Z9SaPXnkKiCtdilRxyIzhrGla0BMV4NNKuDaC2AsNGvyrZudN
AO7arlv9Skjepekix96w8tbDIqeHrfM1q9omEPIHuHTKDMxqhxQBYfJNjtGqObFgYJ6mLwjQ5I+R
SaMwKNSnWXSA57DbcVM3aQMzwZLc00xAk2sl73bFd0wAckLqC78lFVtOPnDnvjFsIAuVTfypv9cW
Jv+VLZjLjsDjkce6jGn+Ue00vR2NdSZapoqcvEiQr1BKcJN9yqATNVqH/Yq/llfY4sIpwhahSzz0
HGBwWKefEmXz7anDJTuj6bvg/li7paBwTVCkCQ708eA0fUcrPrZToXFwtHz6zCKFmk2QNh3m0RzY
ba2Nk/GRrpBJGesN0nBiuRZaUDIP9QEXntAZNC3bStQlBoB5AoXA7Ag7AtdZi2Asyc/66aLh0Kn6
i1aCBV7A4ddGa8/UL8U6lhOEODbx+zAgEfMQyqsTOmvRKxv2q+V6ltVSb3jxwasX1CNU7ne/Ynil
4xtNTuKcW9PMeWTyZJSM1mtOKWAKdctJnik01k8Bx2o7n+ZqcH4aqHib08I32O7C0dPnNVRz/0ll
yJZGoYKsN202iyYh6KmCb1WGVjgpobkuE9Ad2O15V723WT9ExlLeJ4EloIruHi57uMYzsicMUZzK
UBc/VHjgn3d3Uf8IyIoDpLvZ+TMSejU80/kIGkpLkJ2vH7pr6e3TVlSC6oqVvCBstRTjUOAvHdNW
DVXP89Ot0hZNNrGm50Zi58ya5kJgXI5vNP0EisqTL4Ynqcnvxfxf+Fr9sBw9gDsDBOikTqsk1lFU
QGCvA3R+klLCwcJymkO8S4Njbw9HXi2cef6h7hbQcdOS4vE4gSsPB9MIYM1alP5vnIsQvhGjJql1
PIMGj17vc40W5vgCmanTGNs7c37bIthGUkE8qFnf2lAn2R7lJroeHhJwv/RFCmWwKmVyQNMh3uWg
Ti9N1X8VkDqmysbinqNbN7S31hGxvseHO85w1yIesMABSr/K9xdOMQ3iwxIJM3ID1IIk4IPOWidW
VXtb20jEhREv90r4zcAUQ5mgSz3WO2votiU/lhf6CW4GqJO4VpbcPdSr0189C1GGKOZym9mWx6zM
rDrxg+zYhRyfCYEOVJk8DODYkoTSLyAK5AU5eoZNDE019sIjLY3Da03lNWwSqhob+au75sYwGnFV
rkp59DCej7y1JENEC2nYwP0pIxDCwwLgDI4irPj2o86a2f1VFq3HAwOAgVaQfG14MHRGAHVk7ZAE
O7Jk8pgmHYi4NjRQ0s/VIf5AXTGgJv9bttlphI5hhDANkYV9Cij26SrzDYcUn0/MmercNJENVQEa
+pEFFrerPanp19tQaVTboGezrtLgB+JyKPnjipTLF5jiLnQXvHRI8mIFY4UyTDHcxfz4RjNgUp8/
wlBkKPkQ+/9tuNv6tEWnJ1eLPGeRWSIrNuGokwH2j1LoItFEEA5VJQo01F82XOIrOwxOStyp2MES
p0JdeV/rB3xChAhNq6a5uwL/pm4GC6BF06qq4pF74tYjYhbLnRJ92t03C6mD5lRYvQXI8CwEIi3k
KXPlmnN7Eyz65DuoZdi0lG2wamvni9FTXhhJao8d2PsGBL5yd6VVX+TRgEl9JHksKMbtXpHonVjs
yVF+K5qGRcluqZONYv1VJxQNS+cvFoi3qoJ/BA3Iz326GqR/3xShVCZpN/DJXEyAqeqIwXdyJBaD
kbc92Hvr5hmQDeH+zeEK/IKvWySmOtGQYI+kYm5CWFTL1GWnQfBYAOjqv+b0uhl8zCawCyrNmxza
FiC3m3BgHNNj4IYWM0dafNYhjN9XtvatqC+v/q4/uoUx9UfLO8vKkpHiqf/H5Yz6eyjYMIBgBKM8
OfT2s85KpC73D2+uneTd3knQh/voXMj1iW+wT8I1fU+grzr3rFPzLzSfSetuvolxI2QmDUM/g7Vm
ecrxjujwzuglVJymFuuCFowmUk93PtP24nrN2+XLXFt8bgNRyZ80iP9ZcLB09riYkPuG1GfdH4it
b/bbkcY4ky/fmPdOUpjsUmDIh9dJfyEXH94j306CtYgmQ6GTT2NGJqlE+toYpx7CCSXPYlMfAZLC
NPUUcPo+GEOzja8C9IRyMSBLPpar9y5M7VTp3SFPUYVPXetAxptrzg6zH1WbaAnlJp6e0k/I2CXq
mWzBfrY54mJGViqk2a4nyMXXKrkDmgmcESg+pd2WwyXr7s69FQMtjysIOFXY90E0XFw2FDi9iZ9M
gBOmt6bwdBrdJ2yx66ccpPiscY71ys5mp2QYOkDe863GiGuCc5XSwSQV1qvbxBUAIEwr0EfbeU9I
AQ/Pe0ozd3IqSPbGwakgMOJ7Kj90znSRgok42BNJ0nwpS1hqZ96pSnQ1/srNsjYK1dWvGVTYiQoR
mf79qmIjw/U2UQ++QHDT1g1IM5yBk7RpyXH/C0SlysFhLFBqiLNLvSiE968XOnU0BGpK3Un6wO7Z
DwEKx0iDGpxe9u3XqEGeM9+MEuVgM+zqhnlcVSOPteRna7JVNhsGxEXtaLNCZDthx11EHnudn9un
NVpxxgC4p0nckjJHauD/HPoHGTl1L8PcWyNglxoBPcaIWUqMTyn5Xruc8hB9MwNiCIomwcyqOKy2
jvTRQVUjBLBoOh04eiizA6jEQafS5ELUeEiGNpyResC8HdxMa80YUBeRjzziq4tTs95V/39C/F7g
jYJtJzP7tRYYCMI7mfDIkEnI73RuJbb+q3i3d+kTdSJDTg8FF9tQ73/9bkPrCSE4Zx8Hm0NgYPVj
Lo/0tbGYrJ+qgK1v/mY4yjYoMq6L9gNC+WfEgJJlG7JMvSYzXDLLcswzIQAsu4FI91XdChxR8bqF
HCHhBpKiAZk9Wy2DG1im4OHLK+B1qhpPjj9dmBIsEqS1B+7yb0+eNVKnrQEbJRAbmQxHTRuRNb7m
NuSu5YpKfmkDAW8K72tyt1oX/rgVR2fMArsZ6di0HVBf8HzSzNacfseU4CPmHbv/xrPZSbMuEGb9
SRYWoYT8y+2yiyaGLxwOs7zzw7M1W0TXVrQPp3IU9oUC6JE9GK7ATmRomTmgl///rExQ7eBTirg9
rJ1Q2+VkY7AV5HbUgsbLCuTFmXiJwKlBSahBZXS0v578rRCoacOMXxxoL0W1RrZhorXbGDVBsltK
G5h63FZ0t7TZNhNIArqXG+JzECAxDcnFL/oKRrhBRj+Bq+zp3EMPyLkLXsXRQtkr2/72WCpNf+2J
v2/zz3uL7+zRqXnwGKf71tUH/KPnBWLrtTeMiMgNB2Pk7vMsUKXveN49/CJNr3VF8JJSRpylYmCQ
M4rvReIjPhJhJEpHl4qTRNnrhFlOzGI+bcrezSTlE4SVN48TdxKHbcHljFDd3DWyKQ4TERcA13Gu
nRyo0AcMl/U4Pm+8/30PL5Omdr0DsZ//K5temlUpj/SKcWPxGZc22RusYiDodMqNb5WhKF/wKG0k
aLYVo/zJ+29ryTX/CchIc97xF7L+/XgJD2tP+9v6Kd1JJ8DGdZoRi0ovSvzd8IFSD6ppBOHnCiLJ
OiLMFxkuxlpQFFAVECUkxOvMRN43PO6sejFRhRbFYu2l5gKa0fi2XW4c+dtieyUpX2AGedOEHyXw
WKsrks0fv3J/ifbeJDAOz+32nFUisw3+YDgoFFPg8yZ7phEMz/bg78b95HGukMxP7tpe/pCX7y5v
EwG0KB/cFocY3UYgpPO4HrUSRVlbxgUnPyRFzhE7abkkQe+6L4kh/24JzLZdUSlJcHkY+SR3le3i
gujbyUBpUM/8sHYujDXu0beJFWlSUb/lnln2klISSb9HLWaWQuaEymUM3OVL1Z+kbXfWtrC21yj6
yj5T9FFFBEXenCPKAB/rEHedOiYkFwmf6shR2V80/4KATvz2xKzORv5pZgD6lqQhDnGItAL8UAqb
wxEzTbetFbm2eJ2E5H60p0CjA0rXJ67Y5KAObZdejf6J24RwYXe8VFMuFTgYIfAf5FLShVX+XRCW
+tBFW6JYqCO1laTbxDJS3FvdzWzv+Qt/ac+HhkVXGpV+AFvKT2El1MeLeZP6DMjHGzDf3H3RCPur
b7cWI6VlXW3VQRMThaGkB6/Q4c32FO2gR2+xDiVHRDLI2gaEY2CWROwu1OgUwxTK+HEPhwKqQbXh
J1ABfisC+nipaBwtb8vdEcYUGlCqwQ0dhAXMBpT3FdOB7t+GqYldDKTHRyyI7xQ4fiF9Hu1nCOL1
+7Dtrqr2humLzwHaL5mYnPEJJBlNGdk227ApuWR383IyIji/MNZk6vBN9G7uFm1VWzUsUfNaCx8x
xEuvhd6jsrdtaaC3HjCJHdps5lwC4oKoy8JumAt27Ug7ndHU3sAr8CVVfVGb1GErqrD7aPL8MRrG
VZmkSUAKwpxeuA5aX5ocQOrk9qCfdcgXrq6Q/nOJ+GjxIQrosMPZiz3KyQ61HsF9+8LgO4Cl4DXO
qm5m8IMTyE5Ya49Fa2ZcXhTZzOvLs61e8EaZoStmO3TrRoJk1AdhywlIUf++7hppAjv41XUrwdQS
E6M202xCEBgXDl2TZk4ZBKGz5Y8GcPHoV/Kxu7eg5Z2FadG0MkBgEBdBEeeQKuLhf/kbzopoeZAd
YRUUiByCG9z0ygmRadUV0AivL5s7QcAkXWl+z7ioJPHgwZjClaH+3Px03UIcCLEykzh7BLlBBol/
HLEiI6Bq6zu5c02UILbZREtFGc/QMpiU+trZj9knh5peI+ILrIJ7Wbo1hgHTfKxPtOf4rcakauFe
62f4lIOXYtc1pQ4nc7Y+/KpKznSA18g4hwkT3UX9lZ2OruubiqhCGaaLkvjaV3UsKcD5AY9Nsn0j
ESkvGHtap8CBFd6bOUggaDdVNcYIv9QVqeubYY7Ey2/Zg0BWaLRp6uuT7ov+TM/lASzFD59vJkom
85K07XVmTP/R3jKKgVM5XO8k+o1/u4HLHuBfWH9mQBNoMutaoX2rcFZkeaE6gLqA46GhgGVH6KcV
z6FFW1DiXxbPa5LEkid6fJmdR7i/a6YE2UQvS2rwJ09mbSkP4XnGQdiOT2LKREBKJHVXzDn6208h
5nSlKSkQZ6NLc57/FMeCFEJPbHWmh1IQS0aWZOBpqzFEeMy9crlL8fnNN9Zoww1BZo9dGbLB0WFl
/AAlauiN9xk/rfzIjkTMGQG//uBw+G0Mezs3SprAFQx2tZe4lO+FyT30SalBYvxjYDHtFhnNvdRZ
LFAZEA7iLofqZtpRb6bFHbS48GZfrE8DVaDafWt1RPb93qnPaRkiB68i1RLCYuD01AQeqedwDPBF
cj38nP1GHrdeE3TS2kBgqJON7fKYRTCwui6CJUFwX4OdCvIlds2i2xNmbqqk11DGLqceH5gBUuBO
o8mZfLMWWCL3UC1W3wI6gf5xsZnGe8XBF7LrJj6K10LhrvV9dTGGSe9wNLOPhhiAulUUk7RnpoDa
GB4OmHp/MbAc/XXTeACXWAjfP1vicNWc0Cp+aArYXOXP8THhliCjVjVV6494A5aEBC4THZ1/zrsa
gElxHT7rqNPFfWBf7vBVhVh6BLnoHMenVj9tWaiyIxOGDtR2Ps66azmJrnhza2+cyIBlW/XKggCr
T/EH5+sYDD/DXkQQH/ZUHj8L3ztIoWD3C9mIR59mYbvOJ5SMvqTA8KHp9LxMWft/ZuXmtcLE1t+A
EL2SmrreieZk1ZEANvcbQ7wOfc2s3g87uxhI6VKmeaBpgsRX+WEiRwUM581cycVlp46JPmG5Vu7B
t7MPREl94RXaL5sxWIX0bi2sigf0icWf34HGisiFGCNUwGJmtaQ9bC3NZSQc3LtRSHesEhIsQIrJ
BsIELXyBuiOAq8D+tgGulnXhrdplYWjMmyVaL4jO5JV+qZiE4fNiTHY482gT8y/ufDegMRuZ5P14
us+JUIWA6sBPvh5qP/qb3ymjcblvKtmKF5zpLcg0dVM/AVGc05badBhiMsxRj7amFyrZ871sO0Zq
YBkn1XRF2z1YDGPf8Q7wgfqSBe5pdH+MEiu9Y+t+P3uUZRIqPVTLHs7/m74PwuMJR+zSBdY605Zf
Xzmj49jDyvt6v0HUja6GugmplnBuO2oSGMJgPx1aiFersdrYvR86cTnMBP6363tui2FS8832L4Gw
rPnS2PhnyBvdXare7A2Nzjne+KFdNKRAFwijoP+ZEQPsd3YQ2aRzVhRzK/rA0Ll6b5sLz9+3CfY4
QLMoa/+r3ITw/XF8hSfllhC3GFktTeDD/bkVGZsCgRIM3bP26G4ms5M/Q9/h83DACa0PrRpmK+Lz
trdidX8HQ6TAq7umLXhicB9MOR8C2uOT9gBdfIBZbCPAHb4pStDqDoC8G+JlqKD1dLNzYTlIpY9v
ppu8B5M4jBIYxT0FyV3KcKodh8x1KkwWpRq6qA7QDX5nlGRs76ylf7K9me262A0ydTskgUkq17OQ
QEcda/ZVwmLkxIhXntGKM3Wo+DzsXUVZHLffMmCTUBRge1crjzdJH2ViFEmYK9PO5dKCsZllOZTb
tdmFIQlr+HOomUAWwUJmHln6fmx/qtSuv/NKc80EgwZf4y4Nqs6KqQZcBHzQDpUncvZXxKnCuSAY
OfMZ4fB6/5S/4r4PM3KRQgGZcP/T2JjviTeVOZLAwRZ5Rz8The3jJQCuWTACPeXAS4vWqHknqCkk
5ItAd5nkCj3jhxW+rFnO5pfZ3OLXTSckOonUUTAAy/pSmTE3j2NvAsj+aPVRbpWH0cfbnfTfPBMU
XkU4PntuTLjJtupa7IccRgw7U8U9Z2C42ByF6fjnpDq2ZuCiiZLhtPQI4u1L4y5vq25+zkiF8lj0
R5+UPI9uIoRRGlVpjxaoUp9aS3mvJlic8IAny6CuhKdhpL8DYOkDKtByAZdYcOOluGgmHcMr+F/M
Jut+eNmc6DJU6Za4DsICf7xThjETY7y5JnRhSU0Qh5CiJSfF72qvUsEbdlj66NxpQuyfzy8Fzt1h
mNMw+82qtaDMai+zE/IUlvN7nfJ40Chj4D+vOSrDr17RYhmX1TDU99By+cTlKN60XoNMax10yjwk
eA0bfAe2HpMD/iy/Qm98MbfwdVDacvDre9qDxNALztJi6lR8KA/SPJ/vfXl8ANrUoqpUys7GNSpz
xHeskCEm4WDOpY0NrLugLhEsQ+0BfKAXpooFhUR0BAXRSroAF9l5oYYUqjjvLIKuOt3E+ZPDzxyp
gisUGiRzG6XkWOWN2+v4+AEFO81Oh8my+J4PLyfejvu2Inhpc/Iky2iKNHQ9gzdQRAYBlhjpVTh5
cW55+SuJIusAG+BdbfUMYuZprNJjSz938EMcOlOu11uzRYyR/tDvOQtw+mYOOH2zkMpOMnBQHghA
xxytmk+o2zmT3qf5jef+LMkmdaugxDUxDEdt3WPzIfZCUtnmbu95Y6YYx5VFr4Say0+PpfYpGF38
Q22/QcEZtB1XCh+Q+zlR0FZ87LPdBa5AbAKgcgrIQkJOhEEQw1lVZ9oziyPadDTUIxd0f8cKwh9p
JKFDyQRLizRUCuC5eYfMFYS3NZROIdNAAvBHKwXsAaSI1rCNkM/Au0gV1aq3MocntAtBHndJv8Vv
Xeh7nPJq2GEAHppLDwZxXafRERKOJyjaoLP9nrujYV9UqmtvwoY6jJX5ojxpYT7JBgoety9hkMcw
w6+lQNTaHDIZ6wzJo3riseQNQM7SuEvew7lzLhno6KWfzYoBzv6corVvr/ggQFU8rNBXw+8xd9tZ
lZ+fsKSXhYb5h4ABwZOJUzz10vVxZACdGbUCGfG5CvXNNkbqmF3e0KjJLJnCSFohU3GDMeLp1N4X
8jm2zjPQVaGBE/5JykIjV81r1SfeY5xjfYVsnFKGnh6nSQtrwq21OvQ3f8RXv5owEeXQYEYRfcWD
4fjX+qG3dhfQKrbinCnblm1A6tAfHLJx5jJm2a4yYIu+lWjk3q1UsANFrCOV9r7i9xkGkAzeEHlM
M9x/BbAaXbEkHTGZB5O/chnHWKCph6h8xy7B0jXqj6hz2DjAQqbsxNBCr3tGzAL11T27IUzmlIi5
GbSsRmEshFFWp42tvJJb2F9eeEFXWikbjWMr41i6mMK9dL1VGJEyWyxhLJWHMXmXa6BJxO7sPher
QNBrxWIJbVr3XRkNshvueWl8qilz0MC0GVDs7LkiCkkdH1Zh82oxK3Hx0BRvX5u/KZ8Odnv5K8Bb
Vnt7hXIsoGbE6d/GfSpfpV6AweFpiX+z2A77umfTZo7kI+YfnIDCD+PqY7gHD0d5oiT14XsT7Zcd
w/FmNfqULa/Z7niEhx/e4qKcAdT1s9uEyM0ejZtgx0WtKOYR/2sPCNuZVoUlHB0V3ngPmstm8yPY
o3RLm8galpM1c3LzSHxCKZAcsq/eE099pmLjs8WStReu/fK5IbXMEVXdP8Oa9aNnxvThLNEIoRu8
Q9YF0AGTCPpBeSE4Rvn7E9DkwU9n5nHT7VEn9XMI73MOGGqqAQPebyjOYen/+7b1wREhYJ96c2EJ
4zLtnCl+MXrwfT/78ry1UY+I89EZeO58kD/rLcrF5P5KYNbvFEd986PnzHdMhdjHioxCupF17PEN
BEVhpNaX92ExLBblE3v5aDnV1ezCcr7JpX4afY1CJTLE66Cyjt29w7dwAIYTXpXr5nfRHRI6LYM1
Y8QI5VK4T/BRzpSYWJFTxc2B1A+pt7g7rxKlI8UdMp3dn51/sUyBb9FBSVlIHMM0RVwCO1i1GUpS
fO8M1g3DSBFsgBT0gTj/bHFA0L1QKFj04Z/8mjJgqptF17RboJD3rDfy+0DbzXZcSBSyAyAJeYxL
EkD6cTaeSgYH6JlsrX4n2lF4WTG2JD5C7RGSnFDQMRqj9V2DLZNBv03KOKRPShiGslK6vB9HwiC1
YhGrd2e/KjAhefe9GFeVo9BmA/BytvRAuxM1DD0N4QJhxtY244Iev0AF1Pm5q7s514wMeP2YVHSF
KGy8IUAcGnbzKkMdEyw3VI2crOzCx8LWOrvoeDNO1n9ct9Oimnsqik2fxCBKoFdb5X9tibwOL9Kt
e3Ra2DN35tOGNt0ehwkvMM1hm3yPqhOp2XjkNgxGbldWbrDETHLVxbxgwZLDGo3ak7tMMzv2XXr2
aYMtb7NPylIry1hqouxe4dYPMATwK/tflGj5YBmLmkcOSF5kDWnsq20cOUzlo5z6AQWc/1dfS6f6
2qf/81dRJwklepDXnO65T3d6pqpDvUdYP1jFUmLU2XdwsufKOV6t3F8bd5Yv+g+Nu+CVmgr7NYJj
JDq5rZ9yuka586/7G2KRea8vMhwxZd5WVjVCbWzFCtZd2zwSZcM1Fc3vkn23m1RzxOkGWoqAsWcp
S4np/CndNPpixzPA642YHgXsxFDFd1t5Ig2gX0nWL/5U0GIbRmXSbGuQ1cwLarFpoWhRrWvLyReM
VxVS/s/EhwNrhGrAM7tgPSFRLj8i1uw5QD/4RSMQ0e1U/ZxS668L2k7tDvAK4ri+vPPG/+BlJkgs
fAZWAy63hquoyWWEcFVQG+STyq0oycIDDazd2SHwmASHrYZJ9c6u+nqJMPRG3mu3Nq+Yu0hhrHZ4
Olnj/TGZ3iOqcajVelks9S4gpcFUyCVy8skq5EC8Z9Rpds0rYEdwdZwLioYLCZ+O/GxR1qnZZQJE
k/QLS0AvxnWqS1fSWOTE4kYQKhRdXUq3yCKQDoiT7sHbGsY5jOmp0HXAK4ugnYTlfXjeL0Z7lwyz
s4n+R2fPInu5yqoZkvoxypOujWM9rctIF6YEUox0YTMiGhCRs+sOerFphhZmjOKAnmFXJlIlfBzU
fTO0r+bHXrmrf7I7dApua7KgCwUJhD/wfXTe/58tDkXE8VJymkmvDA07Oi6oe+JmSif56nxl2wlP
08gQn8fctj35KaBA586u5m7ziM8+Y+521JWQbLptYZMRwhu+jZABNs0eyhE+AGZ4GMNt3KeMF12O
ZaFeTc4HpH2hoGcaYEj5tmqQgnXOTzIgH4GxcOLphbT94o+J3BXGfdMz8EB3H0ujyR4Pi2gDE9Aa
NAfaZhf6pdmEG1v6MBfbBkSI/xuT3XqSPt0euA6D6lKZqWZ5zv1Hf0eDGAxj60EgJV14j5N9RhOW
zZub858J3jHnHKSeAJOk2v7auQxqNL91i7ECGjrlba0xBd6IMUaKWGM2n4Qa2orER1vEb8CA/sMu
rGifby6QyUuVslGoUeDE6hyyCg6ijm96vEyLW5Qke7zOMxC++FA1FFRM1IptuRbp5gbHAyrFpUV2
srvk08BsONUuMB/rgEc/o/peg9jp1Y3ke4ntGnfMmrNNqFASY3Iror2pyUFlCXEpjNBqkt8rzxTI
4dHLjFc6rCuYwks1SvryQssKAshztA+J8JqLGeJNavPvM9OQ5DyISkXMalVJCkse/wJQba8XWNSO
4HBIZ/+P5RHzFUXDKGekz6Safofxg+XTT2dwBd2hu6O5mdAq7MJP45ec4UeCEN5D2nBV2PUGrsqC
ViJgh4OTvlgC5uao1pXAx4YVzTc4p6vwA3/IUtKSlkqdEYd/IGH0Zvc7Y8rFcgtBXUjm1LM3kbsq
0ZrYPlZW2x017Fhgk+1K9TfXI3oGLlCyqsMeCMY+helrwy7KCXlEusxDkejwpbCMMROz9eT4je0N
TFaxQovJJGPgBGkmhdRYyaBiMsPAc87nhhb5fRjYVEzNJwmRBqEHp/bGzJNr4cjrZcOWinv90idO
yswb/1VhM+lTnJYu2sDNkNCzHBcfQKYUxNJG5iBm+oCYiPZXn0wzqjr6P8xswyg2UERSXdmQFGLg
z0Ku6kBAXT8merzOuq2sSDwrxSQCfoXbZ43rct7nRSemQkv65MaWxIYIhUnXWDBgGhPmFcNPGDY3
yR3qmZ4cu4oyDox18gxkZDJ0imaZejMUfj0VUns6raDRJ5aDvf//84MquaTpqUgXf39LvtyPyWf+
xaVv+2vwaHB6L1UB3SqLKsRfFixwPFuc75n7uaCbn1NpU7FYCfUoPf8T5KISGZq6As7pBwdoZHIz
guWAXx2becPZJSwAFzW+CYx7BU2/Ds1YvYP/9506D54XMJw7mH/QsR3rvnLhYDXFhZms7AJDMMas
BG5fBibI+N02/VggEmKbsgAHcnwb99OaoeLrjxBwE6nYgEGuBvEjmnt7AM2t+4GPSYbPii0uQlcF
OZdeJSKgC1YwsyoSPIQHUYBgoh8zXfRmtfKXn3wZGZzZ4EB3f3tw/WF12eKFnYPc17Bq5tsI/QJl
Eqf/7yHhQOJ/asJRx/3X7I2kJVfy/6sKXgKGV9IFfIrM5MFl14gv1ym/c6MSi062A8r05iCD34wm
drH38LCSfN9i8H3Ad3LEZDGO/jyh7JyfAh3u+bCtHS2iZyQ2PeDuefpGQgAdHZpTXVxKloFNnv1j
pMxc290mzscXYhaAWecwLdeAAdSQAyD+um2VMhI7QjzRrMTNJXZvcJuPcXvmDscxphNZlM9TNfS+
QKJ3zbO/OQ+cRcKQHlUcW8TXmzn8/S5YyK+PsB8IJBpjJI/5YiphxEjoEW3oByV3LzF6qpntgJYh
3MODqyNyNtNBqSMw1Q0NeDotiZuh8Rg6dWDek+HTZdSlFAB/vTFi8z0VbYGGrYeXh0JHXS4LLjbE
XlAuybU95pFy1Yn8i2KiT0jcYRO8+ev7VbjbsV+vWTkJTDeLsYosh8rBAVnHkHauxJkhFAFGon8X
DiJ+9ih9BASJf45TW6jKPr/HC/K8qXiPOUfpeoEaC4s9M9IeVC5HAk15ZWt0mDvWrBocdWWU3FIj
ZwaU9Bf9SgOj1ADKH6ztI25UUYGN2oBj3xCjBVsfHpAk0Ry/r8hd39CWeg4KWEP2l0a6bUaM6bFK
Y90V1QyIevTNEH+ID1/QLS1UAZuhfK1HL2q+MqYGsrwMbiBMg1dQywdE8FsQPD7rncoCVhfD0xX9
YB3NieJ13LGSCgMnRfEkVpy9o/spIK1dHUphExIdZ4M5V3IKwDZRKR72SQc3TfS4fTOdKk7c0wpw
XQYBawlTBH3TzDYejMef1gDnT8MVZ2bMg5tk4gOHMqbaZEXMQXQwzvlx3eyIkYoEnKjm8UHUMMvd
EFAxrcUPaf1gbVp7wOxsBno+g5M0AyR99V/WqQrVudPEpe8ZyXrp6y5vOIlIpoIhx39qOMfjI/yT
h5q2tcmRN5kbq59pWyWvDIwQRgu3M66XfyQtvUQEaLZjLIMeXF+vTVt6X76h6gXJWao7bU2T93HM
5YjwzcMYsqT1oQwB3lcYVt1XUnAYFPcsAJdYREJ4XEMZzhd3Bo2y7tEtNRk+bdEdr+bo0AmPYLTC
Gaom14tSjr8TIzZPdvGScX9bGbjbPhQ8T9H2O2XUbbllFxki6MP9ec0O417BrVAqp2PzqNuqp5gt
7OHRsHJhQa9zzpgKgsFqSErVc2ETx4LV3OUX4vphOqKG+gbfQbFnbtag3BHtedzxdBFCj4TlzXaF
JmOAn3RSJ8U+XHPrIEr9NPzGx5wBgSSty0rh3DAxWHRbEY0fEsTvzKp8yq2gP7+ULOhC8bTYht3c
yxUjA8dBAwovm0Rk/hsIw/gcT2wu3VYsutpG/NRvsANp0OY5agY2Q6JNzdHlcCAsDIEvW1HYGkAG
AXziauYMXzjBfwgy69vW2lW6p+9k0uhNtpcOFSlbKubg6niErrZjKyjVu3vrrdsNpTya2Wsro7aD
lfhzPBFfwQgZoe7Us5DPBPpktbc0wzdJZAXo8d7fTL/WGIDN4ShP/eujy0EziGjOrSmwN9RE79W6
VHoAuoGbYHxpo9PKfreCrxj6enOxRu8bR8vq+muJE3w965xhYzq5FMa864sBEydALoLOHzrAv9vw
gjtTraVD2pFcD237rTPHBUjBalzm5YEjR6dEOf5bY8dX7XrACBpWRhiYFZ0tmATX/ghj8I2LBpql
ji6UdYFSVj1ptOiRH8H5Uxn5DaF1JL7ue6URsIjy2+sR8IieK3MeknMmRbiyNgJL0NzxP+tFWlcv
jRtnuhs/jdiIsk/oa/LCPCsflGlp+fc5yZCqwmgAfXYYn7QLlaURMU9Hi61kZPeyV/A3pZ+2anZE
Znwab9q+3dnXjyeHDz6KzVnn4/+8UujuwfaIwLIJ8nKlgo78m+qo6onVwkqVgVmn4SgISXOUleMd
fqAgmlNip5l/No6iFJrL3U0WOPoZzrc/b78gaPDBQnycAQBmMi6eWiKwvyae9KqkJMshpNIIZxKM
hPutC4usfwajgnnUYMP5qfX7sJ6YTxWbtmBphCRrQ9l6LBaVfNCZCXDl1M1HeFMuM7/EXOcWZmXo
B03KbrjMMzNpubQgPtBu9cS+hciskUL3apBAVX1Z5k57E+EJHdlZ2UR3YOrlDK2LhET8t4Zj0Sl1
BUDn5nI+aQ36gKTdfCTNKPfcA1fIDV2O4BePOgSpFWKU6V6YPlwHYwEjy5WY2IjsYPQn475yYkLP
439ZtpI8iu3QKLUv3E6/FA8emjq3ZaM9Lr9sl6Hg4yrJ24+2S1WStlQfVJPxixdboWAaYeS6HYoG
gTjVmex6iVlC/Z+w4s8orOaZ6I/6h7/QURgGClV+KFF3Y/+K0Defgd3PmTmB6YMt2oLIRfCCd8QD
dmSUQBJv/ITjwF0AOZsddjQDyQbzGDPlEGrNhDL+Su6uBFKbsBN9mNpqOgYIHmGyz92zUernVxqx
qC3C+Ty2d4U5PaZdZ2SFHObd2IUUQ/CXkIYaq3Gt/WuR5J3lwNsyt1J2TXB1FuIwHoKJkR8aqUnN
b6O22JBGFpTsA71K+begTPbMKKnoawaO2svMG8ALGfBngZU5hJOT1M5gY3kEm9+0Kal6XDgoL1tY
564GBG3fktibtq23mbiTH/NGDHd4jzMcX0MXBpq4JdNkZDewrSUaKIg2XpD2GAewH2q9Qj+8+OEo
jws25TrJ8OwGx104rKqRrJHJI39+frYugSoqnb+c+EGgsgDEgtr3B4e6dRkRyRaOH19/nzxkO04H
CYDferM76xVaDgtz9ELuSHzBSwNQK+rbbz0xViir5tJ3piOczmYVqIn4BOTc4HpGIdMzdVKvupcx
sbWUT5HTVlQmJ/dA17CR0LXcP1AcEnew6nmFX/b/bjeL4gP8IGkEAuuGEqxe4fFMUV42o3ai5l7O
MnKhoD92KG0VKmMbguayI5ZHREIqR0ObIiWLHyXCM9omoVGoGm0BS52bIAFrgbH/aaaJL89cqK7B
RIhpxH1YbkYdPM9aQyikcKmpHG09LQWbJh+Gxb23TFM/W0vJqMQTDvCAkHvhxxD+bBkjZqTECDh0
efFY+CbEsMPa90G+D+wBhaGMeU75l0F+4Vv8ncQleNm8+COyebGwQ+gZDjJZgKyoLmQ5+2SJ1NTn
467uSfLetYIpxthXYIQCH1QyqialYogdCwnUFCe9kNXaobo4huX7slN+2HVJAM7IFvmBW0BvcY6X
VoKChIgFYnepQKAqjqF7gwYp5UNyjp850R+ckInL+qlZGnCJhpsHdHi5J/P9FbqQrEMpvfzx6n1p
q6P9Ukxz4B1AjDWr0w7t0Ndzp6wHKnDbzUqn+F+gRzvvZvYqazeBhlbOHIOG9hk/g3/GcA6wfJ8w
NpXtAogU40qevnNQWQsPGj4RebHVX9TSyToS4kWSEtX1r6ijPwiv1f0TFGd456EjQvuCfAUjjrnU
4Zd4G+EFlXfA497KAhs95qC10d2lJr94aRIb6Y0GGCi3pCzIS43Dag7xiPGJ6AMvvMM890CUESns
z08e9GvWBeRraqY2/uH3+tzRD/o+xCElxCpZSqMpDo0R7Gyr18e5wTFU5vZ4/OAnghOw3OTQ0dxG
lixTvipzU+07T8zFkWRaax8KUJCUokasvWUqX2LkMZb66kwFoh6UCASD+6mZTuBgzHVzMnfrlW4M
g1NTXd+pzSG+2DMrWeUsDIEjIPF2q0YY/eDUT2Qz71YUZBNjK/qvKcc7RkUBDL9q/v9v/gmxhljK
CowlGNkwAQhztLy1LYUWdR2LGsxA25KVm4w8oiP4hV07lZThB4KVv0sljGB/sXLO5WZcClWjOJZO
XxMG0tVHs/94Fuvont0X+WZbNGBmHeoe/BWQuswUxwVHpjWs7qjSjElKbWziSMiqCL2UTMjRk8JD
i3eZ6ij5hQlZEbIXOTPpylCoWoerHGUXw853fk4O4ecv+DWNZDxOMoI0gJH3EtbKNi4hiZwiTIJA
GHG8hyZa5udQ90nD0FNRzncDE57+3+WEVtNC1X2gQzyWfNRbJx5unMXwY67nVTZest63yWhAOSjs
oYjANdJaeTyegpt8B96I6b7aMJpbXs7GEdeVtYK+uWGu+P32PJvUvhbLRCO4Dcy7gwHdJi49Ppi0
F+hdrUNTy1kcWQRYjtVsCeK9SFEwSSgkHTvautzqwDpl1/d1yD21hObDqnte20NfxLP5GrqIV2CA
g+XkGAY/FGailGrFOAtKt9SDyMKNWoFjRvt2tzO2HEp4QH6GyYjK6QMrH6kmHC+RXY96KE16eo6B
yMT8EfZRSpw83vQY7mEbWIeDR939r/FczKhOOVUPR06qRs8zJBe0Y+psToXrdZpDeW/lqP0QIb9Q
Z+b0PCvLHrQ15B9n1BGTMevSUNLXNukyE46GRd5czBZ0alRURgnwZL13kcY2DpzzRctszqw+PsNi
FwAssD8/+MwlBVcRXPcel/OQNL/8RNuS8Pqt3iGgrAr/PatVzGLPw5ezexW3EG/GCF3fQsidP/Gv
nOty/pLGl78CmS8Oj6FbqvN1it+h0U6jnRIgoOspFoUXp/007iKfxsLvpv+s80ZoB4BXq8FCB86I
I94FPSsIe31KkB6OUmNL8Bnz4WGg5KDd94VwJ1y+XwtxF2JHL6fi26s5lIIAJHD+3KDeKrI8MAFA
i1LshIPUaAS5qaCPp03mJJnJJFfTjQP+pNEXvkC1Pz2aI54INOHdaYAmYQT3ws1pJ67n7Cd5h58s
YE39vXIs3O+DS5gTk6+uT4gh9F34BLQcXYxznOqSwp/LiIUe84SxjHqZpx55wAIx+b5GftJEkzMo
+Lcq2+0OukRuNYeLOLSuKdJrn3d+/nHQ3DRe+dT/Bz/fblFGJ/g2/WNB4K41cMzxhv6tOphjF+2B
+pMprSZPc0doStWp85WPX3Tr8MnQDzKN7UOuJiQLv/8ksqpLbotNrrdweJL6h1QJu+gMrHcCSyb1
BDfZIfUW2ZxIcK5emlfE9iyDPyVlLyrft9f8iHn1rlyEal4vE3GCFJLgk+uPtFnFbBWYvjMSpoJR
YFejoT+oEa8Bw+mtb58ez43FgFnV0xAXPhGARfZtsPtWhVpWi9hNlbWLdF4/1DUWH2iTpMcxpIDY
ne6VfdEAEcNtUzX1wK9qtX2WpXEYPJjuI+kFr3xN+3aCkhu6FLKcZdsq5j1x3Lv4RFJalB28ynJF
5pEPwofyimlQWKdl/ttSYg0HUGjjdOFcOd2btV2HoEKpzz9bxW2UWLuu0b1elaFGPgu66f+pXB+c
OZfreDtmo6IthPLYg0UM3tA9UBN12T1GSl/ZeViwkq4XKb9NHFC4Z8GRyLytUASyY7wGw/8NqfDO
stCfGhq7ax3OivmFEgzqm9DgCwK9aR+LENtZYG/2/If748FjCrNfs4K7Gzb1UuLwo4niEbKhMeSK
imUvzaEZqBPgNaRyKo+8GxrA7DCZEYt/fHY/fnhurVERKR4XZVXn91ceSOJKsKFO1mHN/SlNXxpQ
xusT2Mb1DdgYwrG7TIpMNj/iFWqQqb9GrUFx8eV6soUux0rYo57Q9Es1xwtGTJx3YC+PjiQQWN58
IuOcBy6mysX2n/CVzixMkOY0TrEW0xtTTp1IRjbcDd1kEZzP/Jyg5qsl3sbIx2hkiqbvXGqZ0kZg
PsiQoAqtqSgF07mO8AgtdBg9mxIC1uK1INqQdKxpCrVevHT2pAuRgBSybGaIB1f7JWobaS58fG0i
P8NpGYjIzFlOXqkwA4/vkdQM/D6K0s8oelJE0eDuKCOUescoZVjjSygyHTJKqPwkRO9LaHLANSIg
4WDncCekgVy8KWLEEYP/Tpym5RD7RUP5PvbcQPq+4QG0LbYniN+4aP4QxW5FqE9s9w4T3krWB1Nc
LWx54Gk0IIgPs8C3I9Dfk8487VmVsxdcPnDss4/JRDUax7Yasb1rZRQqWxLvlHHDXpkZy8pK/yU/
BFIK9B3EY/Xsxz24Bl7AYT9MCxki3MplbVibuGKwQsUzYHXV73yczTTFlS/M/om+CM8tExaqFiGQ
rQAwV0A/dsYJsw5po6iVSYvyX28b5wKKs4UpjdNvZfYDp+QfJhKtbnWhFl4pLb503hVJRsBdYKAe
Rg5TGPASZtaKfpZqlOGg5Ce/qaBhw46/nbD9t3XOqBdmd4m3Jm3YjtnZiPGv3fyUa7+7r26IF+xM
2BCeuQlDeChYc1dleoUOm9/15LuKzksbTeEgQE3zzd22ZOAF9UUM5RCtRhIGvQZ4+ICt6sQRpvLd
CpZpRiV9HWUooRpKSzxnn0But/k1RbLyVQ0eOmq2+hUgMNBB8y+T6HphC0q/OognN3k9xk/Xdjcd
3hKJ1KHoRuIvhVZh9GGN/78C8v7okYogIttOn6q0y2yTnOlx8Qan1vhvfD4KWshytOHlZIVHGRmy
6E+ZQJ/Yc7C02Wh87CmEVpP1oXdsx/dwuKkw7RD63bQwcRXC5qrayEnOYHknV6bVdeA272i8w4ui
kdOp9TdfEWqK7BF5KJWiG7JBOyMaxdBMV8IY2gX2O5JojnI3mhiCw2yllDWqnjF7vsicQKZvj9+c
amcBCfwpzb9diRYh07/WiSGe5ALvJNJY223PkQwIe4VLn66cE4y6TlpNidR6i2S/KdcWwRPYykaR
RLQzuMZP1DgENUgVeQG4ziDubu0HsUtPX7N/89afM5X4+Oa1te48iE+aq2D3WR97ATM6Fm7EC83t
e3PtFe1oZtFU3ZuXK0fIfmbL1KS6ECllipUqFNNruXDobmQrY04S+dhr1sjq4mI+BHCLPZzvbTCJ
ARzDxSTfeyu9UkVOt7dM8ZUI1dnUoNuhnBhA9JNyNfQI7Z/DjNO8b2V7Lbmzy/MVI7u54NsoqxTX
CAcxj24EzMMdMeYgb6ZcvA0h+NzIjOC2HBVfUNhG3jc5k++P9Sag+aPrqoTjHQTbjDNDMCFZE/6i
MrA4SH8OgVS5uoDV4UaK080iy+qLjfgkrLN0tK2wUwA5PKGHMEDKtVy3JwxeefpF4vyyZPqxZCBy
4faJeh+TeqTcUJsuSDiHxfPdh2ZerFW8fJIn3UEnXU9z2PaDSQci8352SIBEy9cozT0FqJLOcIem
MHxOijfuTGVSkoYOSiZYpyAlfUbMezB/3AHaDxcAfwPGVhS4F2lf5l9wm3gxn2QUb4L557blGR2j
Ht1rl7Mygq11u5RHMUbl2oSJSw3Vz/UCnls0l+XsUfFdZ1A50OLHH/T8P6Jls56fXqRUXrmXOeUH
adNez5fqcNZ1PdLZ8aDFfBKmmr2mPVXCYsvqVO5fnS/bQBkOArTB/vyOPITlu/e1eB8b9rC95GNr
MBubFUCJhvYczDyQjQpPaCdwc3JkudlJahom5a3UofC6N2CW/DHnPlP46gUNaSQLHU1TEQr7iCs3
RSvuabUW6wtsJ3re/58qEqokX5isAGz0vGKy+IgFhRQSux629D4d+qmhglka15ZqhkcGvTdc+jnL
ukKoI8ZTaQOAfeNR0VEZAaDMJ9E0AbDdl6Rt9on07rJ5NvcuZvQHcFGZavwpPIpGFwbcBay/qc7T
ocAUtLjWGBavhVsZW7HVkElynUSxi4yugYn08RTEcduePqs1abeCKZMydW9iuxdgeVn18VlbSfyV
nOdHKCSNwxz2Ql4w8DbG0m2cS3zp8ZotpPSlo8VWwkiaZ/LEUyhLAb+z+aUv9Y92S+EU5TKozao5
KO/lihqWDfMK+5DBLjO4wdWHJg2xp0GO4p8e3QZ49MZ9SJAzYySYYWK0TW5NNrq3HjdXLimtyNHx
BKr9CofXg+j9B8r2XKLgiYcaYYlA5tqvaJ/hqjiAbhKwEogJ022OOkO37qkM1wp+KxIgwOdhsJIM
788DkFUmJnUS/4CRWHtqavVHseTkaGniXrtQlKtOjKHCt+sfv5u9L4K6LEQsx+Uq+z5kbgLW/rSm
nSa5XMSK69YGZ1cKfrQjigqL5HWBtcRrXOBe2ThCjKXPXyGNKOJAAzqKhVUqySl8Jsp3aR4pgXNi
TppW5ab5xa2M6ynEFzsshgHdg2yomoGTl1uzU6KHe8MmZaR1KbGYy8Bts7fn0KSpMBWOPyjBhhhZ
I1Z5XnIef7W/KE9zCfioAdh6m332PVejJDvyT4VLCPbi5HdbRoFdDTptLMJ8nnKDf1Dvo6Hoqshf
MLmlL3MW816H/uZ1/ls+c1wRa4aaSxi3OKFasEhbdjb3Ur2P3MJ6DvXbRsNaTV83ARspTbxoSXf4
hwFJiZ91z/hrqUgE7uWzf2jTgtx2C1KshdpIwzj+fMPue0+kj++PMckankJ529umH7775FbedIW0
F2xuVnbsW/+uIRY0QUXHp8ZYKojhFW4JCZubNnd6O5BZmppbJ5faDk3lmLgPULxrdqR8gURwpbp6
UeJKJTEpg12p+CoFTmtqlgqkShsfgbO8wp0spNv4zMbH/nmPqDMgY2OtbG8MFHv3tzSb2O/u812H
ZybH6RS/ZoRWNR/JWAZqaWxJWsPClNfYKxtyDdOct715mCLUo8NBbVou/GB+y/bKiwoG/GbZqrkB
j7FOqwUY0LZd+UZQQCEhoZ8rEjnZZVfO0pM46Irmcr2OiRwMFWqRM9s+2Wmv3EwOtznKgf+R26hB
nxvG7Dfd2YRL4+PNE+db0gKI9cT33hVNlKxmK+LYC7gUQYM3i9TaqnT880EeMKdS2ijtzOVIcDL1
ZVvZi3YGE9ijYwHIoZ8E+Jsl6nj7ds8guiRO7lDzP61B/GgHx9RQLlnZXHAJ3dtWg4CqJUSuuVQ4
1VMWT/lH6JF96mYQP1o7KhibB1OEKJAEmUnLZCjGFYONDNuOjF9Ru7cp8bTzt6qngSop6oDEuaS3
OlH5LMioR7mbmRXJmYz12w3gZV3/x0mJ+jyKqZ1fyvDqfjj0Z/1uMg6gDBbDAS+mO6VsLfzI1U2T
u2qxuOm2zuugLaypdwyQraBKaTdXmez1iWXiCPD7GbG7RQsqtEMfoV2dt15CFllnbEz8dud/aFl9
HeUSGFYX20lHwUAwnEycNY2r3uAorh39SAwPjX1J8RBRtYozGd/3LegFc1CwjHRlyr0mFAKE2qPj
5XYESZHi1hZbCtYCLgpL0rZ3dJHIZCvRLSJ0AcR0X/UZNul7mKVb10NNFeD3Cjmma5+oK9H21BDg
B3anRnxrbIvJsgD78zGp10K8bg01CxrAXXlWiX/5+FQQ7NUVAe+fhpwCUk4uNTpQMmvzmmb42iEW
5gdlEZFyP1mpzYAe+MmZveRgQuP+f6JMu0fBJu7gZBNcvZq9KhCUt3WqhOZb2thMOtP4x6Yl4OFi
OtgE6o/LJ0LPQA0bNFK/flpSn1Am1lUvfEUChBy66ZeLsADWj1yfHnzrTCFuoI8s37jHSCCHCTGd
ZhCVm6bDxLt3L7/LtmzfQCRMB7CZaNC5w+N9A8Cqv3K0391I4jmzRUst3tVRoyHr3SmoaI8kZ6Rb
1xRsznTH26dLNh474Qq3qTlwpQgSr1d7Y/lyDYq1pCZiSUZnYIqYSGoDIJ+xHQVf+3w2SbhRkML/
4ZpKFn+54GD2zgYz8BxYGaQUOfGQ3oK2vvU+VOR54Rros+/5T7WUPq3xtZDu6kD+n4yRcTKwSeB/
KZvKOxsHMr7iE0D8ISCWx2yMauB+iX7ufBu9wKj1Vu2vgNTLGwviMNplWM7Bn9LrbPvEPvb1aM8W
sr8eC/bUfp423Z3XOPb3DZH4Y3aY1bh7uCQojup7ktUJNMQJP7EJkdgIaXfGVvEQa1uBlJgbp3lo
TjvKW2PzaO11TdD3z5rcdvKJZmlgPXwsbtzQN46WOUC0jPKfUtnyPvNiJIKB93ljT8aKNFG5e0VI
DP/QOpYVw0/2iIwmSwTzy+aZfThpiQZBf1OyaxKyNbyK2nBnsO1TS/qx/5+XDVRu0T8iVdmeyAn2
fPS6TxP/o3/IVzqDOwrFeMU7RFJX6OuFxGZOTiz771WVkfCqNa99L6RVPrx/BGyYAbN8wmu5fKHA
FsjjNFGYkTjk/qifVt0aCCqWbnetYnxfbV5AgkdZKsceCpxgRCakdq6Vtj47Cu5QENNkYqA4qn7Q
Wj2Fnk8xAjLCn8afRc6Hns9lOO7B+GDBmwdyWrmt4pt9Og9x5hk1ZEt9p6O8+q4cxI/zXQUGEp8k
Dma9AlXsxhXKhjzIwrGv8zhrV8X3gDN0RbCUeV/KsNDOb2XCxiOo/xNm2hpQxw3dAVGGtrL97N7C
4UMxS7hpAnSRK6D3AazR6XLQ+ENe78yGbUfrqzT7fVcQ4JqEMlDlxc01m3ZK953VySN8zsht5mzD
taryqhUnN2iAL748es87zFfVO8JzMi6SB8HXy4ojCKfGz88p3YjCcEXfdcOSuCkZLV9aVp+2nqD4
d7q0yPW6/B3twt49gouL5lOtYa1ceyVoD4pGQ5fTPpHMcJtbwH0YgXanK6wqB1paVRYeWFGpLTgx
GNArzs+BodSTQehio+JIc7XkFZjxCjazP1Aq4PnU1qHcWsrbRoNTnZ+aF4NV3tTWPQZClVg1ZOmw
Jo54Qlk9mnlPZKSOP8nhSzSZJ8XPA6ek8EWg3kO3Q0oJa+zPFLFHRBexkAcbmry35PJ6qNy1V1ok
vkjpoXq9xjZaBd1fctLRYivhMr3OsFzzz+aDiBHavUlmQmufRDb6cBqLH43fF1tTvFtIrAKWGK9M
wgvFrsb57xEbieIvt6+1Kj3fmJH1f8KjRcAK9geKNMzsZXmACTGBXzjnlMhQ3A2P+DwXomxjvf2n
s+iEQVqkMcP0hRYMOHemdBLfPgzKyP/j09LgvKcA4l2EvSWcPqpW04/1f4qXV1O+C9d/kaKK+Rkz
yY39nJPekpOOQDbkcgoD5SwUFmxqAYKpkIJ5MUQSPzxc+EqcXdyYOnL0FcGV8kc8fcusuAfu/+Jo
m/Kv7z1X3ODivOima6sjH0T1yBAwOIRPTIJCJ+X/2KXX0pUCOnNNBoKMdw9ClwV9CCP/dNiYpJtm
VWj8roT5Vtag/AYf+E++4QoZiSRQFbacWt9wVL0YJ2YkpRqp5TRz+D38pFaaSqubz9laIOjXqido
A2RuBGBjAKQ7WhWb3Ibgqqwx7ljUmM7tr0bjKHQJy+3sb7Ha4x808u5NLPu0dpkPUEVYnu1vv2XS
m6ocCIn3PqE8YosJiJjNWRyqUqvulsATfe2UqKiRoI2sXxKOVN2pX78jJ6mKDI8olMxPdmrurx1t
fp2KBFgrioCT7dIPDK2O52PHvaj3iot+uAchDLA2XZX7J4/GGBXvofENFDbHpbktL4a5/h7lYcAX
7tRxHOARvEMBEOCHaIs6MdAj/SPNCKM3KAeWQvDltNQSGTV30LRprzqU3/gqIjWs51njJUyFI+yS
PXA60B/p6dV+jylTyZsRX0XAyr6p4aeNIHh6ftggjGLxqE0OnuvThuIyPIlRVvLncPXBh8ouE/tZ
L4ISOBu0XwV3SN0zAcHY5+F14TqT8ipjYjFU7TZ7+HFvbSBy0hOfbCPD88M19J2PJdD6IVzHoF4K
4O06ZVj5A9juS44mge6nt+XZp4gR8RYMr8BucIPWNN3G7osODrxOhjzleCpJme9VyMFQngy9OSSk
rSeT++W4up1YQva0otjceKJOx6Z71hoOXiafkGLTi7YKP5Mn007TLEVQwLDzVTZBnomZohEIKg4h
Xtsmz6QAjyvCeoPu4OtU02fB67Yodwslemj0AWPGVOEK/y2OXHXdrHuiAkeXPIGGSR+IRsx02i0j
AAdY5V7X7XkgMWgBdL5p3cf5dCZ5VaAcCukdcpdKXy3PtrcMKS+dp0eybJl0k1CPOp5Tjre0M1lm
OHC3nCg7d7jhx/oQBEqzuZyleLsOwkMXKULoM6NPuGfcEk2DVUsZLF45XxHCcHpOp8uq4t115ZhA
HPmZn+WtIvpYK+5k97ox8C/fYx1CABVgyQt1ncloIFR3zfi3h8gsJqtfbPHODIPTv2AQzAwENfyg
Jxupyq8/3ToYGqswR6WEDR+N3pC0d5qmb2hkbtkWaPUX01VnmJkt6BOf5tV35fR5LdwCuBGp0sRh
+QZ/BSLlkuamo4QgMokPRzLFIjseYgavq4fK9stRanvMoWRxHprb3qhF2LXtEiShZ3UOJ/YUy6oI
aOWowGLRq/2pPs3/+FI6LfX3PilseAACFV4bg9iBX+7/gQ4PfHhCe34BXtplVtnrUvZCB1MQMBQz
UgLPz1i8WFkJETkXFplJA3AYPK15IWSv8eYp7eGJ40Che59zAWEzBNBDJK6LOtJKuJ7sJiEQ1B3l
E52eg/srqB1RKl3v85Vc92xuNTIxvwx0z5EUePjyZxHfWBeYqslEEFooIvQf87okr0/Vzi7BRU7C
5NIRJcz7rT35BheWSit5MhJz0Ia+FFJO8E3WGUN0+h+GZRyRQ/ZT9zlfbMofzKFg6FPbrgPaZV4R
MEM+K7ldH/kll7o79EG990tUX7QVGEY2usXUAQwHs/mcwodZbvQbbq9G6oFOEIb82J6/aNZ2ayzZ
oLiRKf5728Zzl/rlB/VuUaGJRMsggikqJmCv631eKzzRmlkGC61kU5OgZmBEO5EFW3BGHtJieS1n
Pkzpuh+EKGLGP9+QHHuVmnyPByGOKq0ppNwUjoiqSpNENYkd/bCDOpepaHMdJB4m260v43WYAkk7
v7Pld173hHCO4PEmjoP3OdgsrJgZNDqtG4RBiCq7pkfGBenXc7IFzJzsYTj/lZoImJQIFO90K7Tv
D21GsmLq3RlSu8f+pTdOKdUbzwtZfH97+08aZ9eSxBkGWPgZHv/L9P+fV+0DQwf92vd2OHJfgUaw
4eG3qmz+mnKd4io3ZnBGnaaBn9c3SexU4RZBb9STSi6dVL+AcDM8S0NMkctZzqaiG1ePHsTubWZ0
OqMfDCejUm6TnMKkp4ah4Fmic8u/5XaxCqbXD14kVPcIXp4dJBSONNvV0384ibEKRP5+oDNRlpKo
LHpb5wPjHtCFaJFOwZLznnfJv4H/XgRQ+Jevyql/iXoz3YrWAnttPzG9LJkoSxLRaLm1nE5AepFl
TjNPkJerK5jT0B6ryvTPv2DW3TV1+UIjPTJqumuTr6WIoPPAIY/VDOytGaAasgLjkIva2dI1lq+k
BgFk98egU3XnBVx+djbh8XxrDNg8K3U0x4R2SsIAlqlalv+3SKq9sVyp5G2stxeVrC/ihHpPYAMN
6N0N+lgyn7WBS5bl75u4U0vTGooBOICPK933K9l/ElCRGoRTm3pGDuj7CXagOAyNxzzzyV50n/J8
X6wR4gk6Hj4Tfu2yCbml0FOdfc45zw5n+GYs3r9E7dSB7mNPWLNj23+/2qBQTZb0B0cawtwP/sPq
p00UFXwH2W8uWMfkqz8kjNizYmQd5zH3YkZNQafMbEIP/Wsqvi+WLYDzwoaKA6a8WpPuP0TautcQ
HFxtKHCIKG3iHCEcdI9rmzoYNUz+mqhx+CIcbL7pQzDjHtdv9hgbpBrdaktbg4aCXiaJjcW4oY15
54gk++wCUzmc4K8i7QBme5AlUxt0syY4vCqlRdEtY3eQlcsUA5MCPXjHvxYu3PL51xbmXQWETmQk
uL5GIRMhwpOt0P6472ek5LeopcC/fmWh5nNuxZ44zm+/CgSa2RouRfRPSChy9NhutMnkMDbcgYKW
jSZT+vrvovT+rUNsnfZEeJ2iUuw5rycNEMnSm2CnBBkaUuE712gL/llac9ATlh7qNmeR5s3dac0W
I9frDM0NQPOmGntqWnrTxq0rQ444XTBLF4+UcAYQVMkR6OfO8re6hSFvFf0wnlQFM/wI9ylVozwy
5mDzzkkpBXsq3xYMaAPiIvmGozOpKSFPmi+pbHdjiY98zL0lK2n3uW+pER+RKOAw/95sW03opjzv
hUDeWthcY97x2Ub797SB2NBJVeErZyzDf96yAfB+7Xl9qcKPtSzB83REPGbBU5ddlmEhTyEeN/l+
hJIkxAxHmMrXuu/neCalT+lWauooS6jej7Ub1aG8v2Zf8E32dXqnMUE/D9L3+L8j8g64LZD4213W
N8Jk/Ug6R/fgHwJ4GDC506Sa6/OlL7XwwhrIUZOOhUNeAr5k/yfVBwdc8FQeeVvlhgBRhyVCojFh
/LvoAFpxplCprc8gaDdBy5Z+9IznaaIYpQkg1G8k2FPrIJhpzdaro6iLaOWuAE3NnV0VPT3J84fQ
xj0NwMzq1mkWqEHdIxvfGt+mQ78Jl4EStwJyPJLkWTEuE2SXud2FJZzwetZy5FXK+Cp5mKh7U88c
6YJUXgFbMD9iK7MMHCjCkeSOvLlHHifG+2blWQ7JL5ggfoqRJI9lQ45i/+hCaKFgxDzs+yeTpvad
YiKp3t9mH0lpPwOrdER3tC1oDF/om4LKDF1Dz2fs8JNGIQ1gO5z3KOEMIAfrUQJFVTSRM3j9VU1P
7upWnSDQWsJcx86BdypJGMjxnXqOByxc24bXNOSh5WgRlIxGMx0/HpBGD21X4KL2pWnK/WeKFgPv
5O9C6FgnuQOnOGc6+mBmQ8uDWpimeQUXoQCmEczlz6FeIYj6/22OMUUx9mpw1FZe2ykJpFiXsbrZ
xAqb6/lTny8xe6t5xU3/ygWZrb0O/irUH47bMkm9Al2pvrP0RSHCDai6mNRXXhCRkqN+vEyZ9Jvz
AZXzMLjeSVBPNLzl4WUP7kREiTpKJnXlzqKcCT5c09GV2hdYpoDqPgtWhxFWOzZP9L+HXIJUn33h
BX2j6J9jwx0aOVC9yCsMZfvGaPgy9rx3MQKCuG8vCMPWlrFCxPA/MS5Zsh01wNQl4Cqljd/D8AAa
hupvWLVF5A46f2ideyLTqwJO98nLrqHDi94TTHHD3lkMCBXWNsA3J4G3jL3c3ikv7jZGsAJtZvX1
2DTjB47LbZdOubqg9/iBQBkHb9guGw++9ltPbqSQLaOA2jNcL6C2qW9aA/3CukkJ7O9oHdMwp8IP
pxj0ezZHltExzh7Y8FMozng6E3udu1LoBEOMkLE1Gtb8muqrRelZ8gatdvn465YV6xl8i1hyTNZX
AYcX0vprCwS/YH95CqT7wVQUjPTBm7hC4qDMfIXqaphmsyPZdByWeOH9ZMLAsl/5uWZKAdo8amXP
93eap5j9zX0+FPOdZj05HRl3zW9TLpWrq5K26UmsRB3pZ4hvFULZbRtnBMLG7iD6jUTe6UNuaGGO
heQidAF7b2o7yZ+h96ttMStEnkCfGCPgKYNpFviqpWZ6W/+PZlo7Gum6Z/r0MssEVot6A+MlYUEd
SbKZ0OmrzFhQlzW22j1/0/4s0eWw+AW0rb/yJeESRPfbsjv4DMrMhkdjzCIf1KxtjsmoBFIdpL6N
iMzUYUK7r/k+iC6TLWVFRApRd/tFfGmX0j2ltLwgvjf1/kF6gUZcIS8TDYhwYaf6fHQbh9J0efx3
ydA9y5eIqv9pZI0efJPKKCS8sNJN1pAFhQWuE2GrrsES9+c+ZJEjq/yUAn/ZBVA6Vnn+oA57fuaB
68xihDv+RhRJxkIGhk9XxiT8bE4jECRw3wle7cxxzr2EXeEqtE981NjrD4y/ljDGp8sODMjz/hox
v53YTj9aZ1NyQ7fc/0jmueR0+c7nwJ7G6VipkOL+qndEgXL1a9ixIrX6aGJUZLvMgji5xCe+RcTS
yDBsdRkJ9NQ5oU4bxy3e0MSeMR76CtmCqtGVT1Au7KbJkRBWL4gM/9+HldwsJOxLbDAsfK+qfo5o
TpPt4ghJK9yVopRBe3lSXRUA+9DNhjXzKQyBTjSJi2yOomiqwUavp1mE3Ht5+E2ge0kgH1/2tREH
dhjia54OLsNJdYH6CKUHMsdfsdTh1FnLmQ7xoXTAz4zP/hNo7T6R9VCtj1B/Q+VqJRFY7jnD1ceI
2zeMNfD1zQwblOadvnadOYaf2YtPEBERVTsS3dbQFaMtr2+ZIbGVWzZjAhXSoVhlPYrGOPzPshtD
ur8z0f+bgpAlJLCLnzsz+0+/C7lTrcxZhxoRIE9jy4ygIIPepTJDkZqJoiFdcj3HF4Kp789uxamf
fLOPnRfQZ59RVyHtEMKvMwatAJmCgS5DsaVyup1+tx+5uyq4xpMQQkEXck0X7q3yyVlDUH07WskW
JgJqWymR/Ho4qx8jUs7rnHp/IIZcI4SECFIn2SC/QSRXgF0D2mxBVdA7NY6rHn1B137EOOMDeJJq
GlNl5sU81D/K2Wbf9tEyg7qQRXFMs5bHbUj2xiHeIDx3F/x97NdiwjAFczefWHTRmwfC1dYbdh1y
j4NgPDCV6GCX3DSQ282/vUCJZFxwLrOZVo0ojQvGCVVffd6+1EC+5JRuPwV9yWh0c/ECOA8fADL8
4EAeTKItygkVQ+Q/TkwyIX4UBHum0PGYy+YBQxpH4l+UmLG3mjv5HIRCSehWJ0g7rdFwRB8/Md8Q
akww99SLMr8DEuUm89G0joSa9L9Es9/Z5x1bQBGqhdFrqDAcycXvt6Vwk4tqmOUC9fdbJBMI+J3s
H9vX+FpJ6PXZ+otWw+CEabM1Hh3jqx3NZnurrGMw7NCLT+z0IkacSb4vBbKx/xBc/4GEzOaFOnln
CR5KTckAqaq8It6ijOIDc+vD4UvKFAN17TYPBclDenCDS+49Zo3FUV4x74MCp0HhrkPib76IuLf2
VfDr0blGjpC3WvzulYIBOUz037KhH64Jhup1Vp2+ICXrM9bL7r0wDwFw12yogQtPRCT6hMmyNc63
NpeZNV4fNt+wGDH4mrMuDv6YTmVEwIW0aULQWIcy15GcoVjQHtAw6PRAhUJHVMfpLFRR6ONkW1Od
ESSAG3Kw212Fg5TywjzwFER1Td9ukK1aYLC3GKz0z9EzZ73ZuEspUb5TmftRllbmG1kwS9SyS/Kt
M6iAN3WMV4EI+EA0kOmL10WTGhqC5y4gHrdBKTRf0hzs2ZXraeDb+At1RWnVYvIhshpt9RdF8HTk
7XrPYff+u2RkoYYtUUlbYhTr9nGYfmqouBNBlchOG8gJ2Z3JBGsJhY03TOpRUyotePF3cn2cpm+Y
76s8DvdF3euFkpPgXGbpZ09hYT/OJEWFLS4wZ1Y90I+UCdNxizoDqN/HIeKErMdvvOmCSzzPNJUN
0luzj4gj8d71+GIUPzD6s08a10uSwqYCPb+qz39sQ/7Ytb9Oo2rWlHfuBgc44t5FYEEM5vLwLXkB
PKg9zFUeld5ZBUrVd1gK5OBMsTaqkAIbkksYm78vQQWpBMXchUKhxgygkEUT6VcezzxuiKSL46ZN
84i2DSOtO5TeuXpVuAnX/5vfqbktK0ffxGRcslfXiQdRuu3lqcqcJu7ntxp9HwOvL86yJjpC53k/
Y3BqJm5d9plfD0TXIuaBjZ0GO8RZkZdTWJsqFfuKpawxr9XWcpWDyR7D6d032QX5glVaoUJMlC2U
JQOxtX3iIdVpYHUfYvA9YrTwLLgZVBH0VWP3Buv0EdIswM089pHZR+Sri9vbS9KIFW9hqYpnhVyR
2UJDkBW3lktGqjgeelVyM1pCspbN24mz7F9bPes4k/NcJgCEsqQ0VvD0PE9ZaUmjhhvksPF0WLWq
Ui9uE9Cd0T8aVN7plshez9r1xidGjNWIIlFF3eWvHvl277gRMf6ne6xvwzv+pnnRkmfHgxH6zYlQ
tVUhvUoyL+eLhjumontLCFUX1bjMG/UXr9vSiRsj5uABz3lgHKQSlMbhf0ATm7n3iAHsNuGasOlN
52Cy6zKyAh4Wp3eDo1KscjX8LskunGk/jC6P0EdLeFoEEQxQOe7Om25m6UjQ5Pws+J9JgWaG5A6U
S8d2j6bxOFUPe9A/SRkJosOOluiiI6villnzvDdxnviKLCempow0o9bLQODO4aafws5M255Nc7fv
aASK7y8XA6jCgNnksyfxrqhMIDfPKLX4+e/xRheFYJO7Aevjd2h45qrxAc/Yp2WNSbLimTwOZHhn
kEtxxO2dcolYDma3kSqXE5oFhi4DH32kV/zQanMOVWxsxmrWPJ7lCTCcKFc5f1GlRj4a1mc6CZMf
31T6WbR7vlmjFMbnZ29anu6OtMbU68IFa19CoM/X/SNW3k9sDvuIIjTpnCfOCJTZzZK60VWxAlZr
rYcGZDXCvst//RMQvWTGr9ZOG2bVIjSxvpMQyt7u4uVf8xziOQwOoATmOOjh+WEpcl4+k2vP4wb7
rU99RUZ6T4VKcrhcAScfSMDOI4QSkx0IiuYsVun0frN3yf9ex5MmyLiBK4B//Cq0ths246wp8/JC
Akpbtj0mST3B0AYD2AjQlcC5Shfdaa+VIUNi5OxXHwwq5cb4rSSSaUcfIn9hHhZa2BVH0Uxr5Tkt
w3iv03QatUbxGdejj6VrUbDHIiY45XfdGeMEQaxeJuJWNT8sMBd9OVcSFkx7RQt4zsfQh86KUs4X
9huUx+momiw2LE9cqkjzfiJYVnKcb+1fc4BsH7Xi4AJu7Oa/Ek6EvNxlEp8AxOrA4p0a/O/ZymfH
sPFIW/iyR4dTzL4GUOppgJRySMC1+T5Xptg8Kzao89sGgh0VAiC8Q0o3Hwad1+ibewWAWODm3LCu
yAlLvVoW5Wc7u6wRkUe5DiiGpGO/aN8MsKTxNprdkFpbSbY2RPL8NvVC7ktCCCq4jnPgDOhmT4GJ
tEoiy35k9Y2p7F7tbTvYfqhJL1h76bdVKEK0HCh4Ry7fOdQLwMhAJTCnN4OQNGTBITM1nHOfNYbp
Hhxz4Jbf6E1XiFQN1yydYnGr7RZB7FUeTER5wBTDsprs9SMURai7xiYK0Bcxy1o8N97L0vXNZHY1
teHX5EewMTQnEpExuRJf/eS2C3wgZYUjEQFeBR9M8gkDsecuer/E+yRRtiNSBHOWxBpHtB+hBXCf
pWzcIJ4r9nwrLD0uD/28B2Y7S+RPBFZmKSbt3qH/LQ11npP8UGFhHl2Q3SDhkk48tyTnLty8ap2w
fiNM3EFhZI5MAgB6SQisuJyqTrtR3uEQRLgHyJUTzazijaZ/kN2tZYh631p/cRgQnt3VBPkRSIvv
rUNMfpPXPpFEwqJWBg8sHzwTBG+acpYZ9sthUsqdbMM62vu0+MRneJ/0C/FquJ41ft8ijtzRGcAZ
iKN041ySRhUy29tU6EUZGExKqSs+tg7X5nKdXtS3H5d/6NGLGdurUJYgkb3EHdd7yVbcSPiIAyMU
olK3X1qOrHFstqsbLLdF0h/z/ag6N7+kkmbsOUMxBKWZddkAIKpGd2pgYuxJmkgN7NDJFCTncfgc
jSkdxHWJZGTHP5TtdJCqMCh7FBJRFRESEjoGRBqKSdgWmEpySkRAS79fBo+g4xiu/W3tltvsZrMN
3UjvZHfCDa4erR1n7/7/OOdKw+zJodT8X2vGTPYUKD0AnkXVMsxC0WldCxGwAy6P3qJ0QFk/AMH+
jLNvcy/d6uFzYCKezhieVTZd2MKwhMknApP10rdBifFQiLGQkA9tpbf/rvxAUDUzaws14IXxupoE
BiM47ujB66vpccyw5WnlJttWt7XulJoLDLLXr7uJ2+7wAn/KrXsEtItC4HOQ74f/r0wUZnJBoSXL
ABiLnKhO7iG0PFhrQ7YiL9OocI0Y1pF7nsvy/DQVNj2iuJtqBzQ1kufUq6rNa139oJguFJKmq9ac
J7DwO3Z6fb3VRuXkQNE2BubhnSoRe1vrupptmfISpYX1PdlBxTSOe460FGnkUGDrIK6UanhubRPQ
L0Ot9Rrg2qTxNxGaBNHHQUfF1L05IzrxMuzmtRH3osTJX5hw4NR/0bED+t00LdPECk6tKZZIjweN
/wGHSdWFZI9BO1YvHywLOIA3v2485YVnEPB21PPmV4I4SauvjGVBo3v5zKBnPhLNOPPn1FiN1b+z
i7M5SrdKeVohKAB3TVLq3GSCRBYRtjWAGluYii7aV1cdsf+Muxxour5C5yJCqBVQVupESfKEBsM8
fpwAuXKS13cEt983ZGStVYaLxbk985IrsqM9NQC4j0NbIr2a/9aKJblD8aTw0+SCzDHC0sIZNKeD
Vz4o7Mm8d2dXjTUqce76fxZjExy9HRKFwbPlf4LGTjl3Txs2A6sXH5bRcZo/jUK/0yvxSHmOgCBX
Nsx7ctXVCHUCaHoKECZUD7nO5A4ERmBb8Jwb2fOPF8eVq0l4GaZxVzlIONlsMxhuY4fXgAOMjoFT
ER8p0/QV46HKeZljQqWKjTeUPNWSby5eqMIyXG7JN9l1kU3sQBS5u2jiO2uS1h4iL4lQc2e/aVZy
L+8hffXpbUoljw3RuHXr1m+rH07KENEzP2UovrItUOtAxAmDQkLkI1RGb7hnW6OoM9+41l6OuKsU
fMocOYxu5eS1kTCmYdpDtzy/LC/IxAphJhzLXZUCSelUZnYZMgP3X0TS+SHc/Nz32xvcB7/iPemk
mVbwhyQNxjPdej47TT5EAuIEgcOP5r4PRGoYZ6ZdqErldViqr7RO8ftZKWR8BlJ3PX9JjyIKUI+c
Jsf92z2VD4Z6PxVueLpkaiaWvM503XNTOpsjEoVy8ZFkFFDneBThrWGZ2p3BwvpA9dNK810rW+ln
5whRqlKKobs1KODdcSx3cPGIdgCaykvCyUbn1sYiVHXgEkJ5PhOgEsLVJ8i7oa8q+DEzLQUYHcIr
pQwVZMDjWsmaKL2bP6g4z7uYPGCcLxL9nRaz1pPzOuePcxIiyRN1ar6kCyqBb+CdBVT0rZQOC8hf
4gmwoEybN8lLg9M2QkTe5iy5P+nXDtx3O9uWm9oIxE+2Rqe+xWffv5XlqZpC5nF6ckBUMRdx2Fod
v/PUmoiwV4VU+GhjwvTpzt7SfabN/VLSGxmCykY2SY9k4v2FkbIYokP4SUZxvru+HNmDg1RhPeLq
05AEw/2vkAAnA3JnFBo4g3qLfl2do6aQth5nXKuzQkTW6S638TL3zKSOtaKpg9FoxYQwMOuQiCc1
ftQKwr1y649HozXcSlcrNOVyAdObgiRy3TER2s0OvigllezjwiOWKYe+v65Lpul1cIWUuA8LJksE
cYuOQbHuHtT8CGN8qa+iNwwMElpBZsTFFaP1CCEePae7b4EaxBU4mq2tCC1exYQL9g4vx0L2T7x9
j66AxU7uiUIoSo5oSNA6fiklyN6LIEpt9diWWHccosAq9B3GKzDa+qDu2ptp3RqxXDuDbgpT1UAm
BHfyj3ptBvUkTfy4IhQGApDSULuuesVAC7cT+5a/3tHydex6YOOZhNK768mgKwsafc2v/zR+177Y
yir5GcyciPnJObKM3JXTOqNOjajpPeFryJWCeENL47xsHstaYgvJimb4WhwaJGArOu6GJrUKyG2V
Zy3k2lU8/9bkEu3uZutVPYMlqOYvrxyB1u1NmIjGWAXX2Y7chMJdVdZpKioJFKkmHMuHGHXJb+IV
UuGsPLrWG2LWBIsRcuEHg1BaCHQ8/k+kjiSYEiyV7+xKRpjbli7HeLxBtQJGW+jMMYCQFrI55kdg
TVrP/PUKsHBPFPJ2qqGoQ74Lm3h9V6so+inZIZlxKFxjtBvO3YMTWcr6zJzDtrVWlBPMr5SD2j6j
qNbUYBO5ciXfVCUj5P2uB4oJFVNkaUBnoHZE4n6G8pxmLVxyiVTkQ1lgEZRLgvNoY5usJz2/4K0C
v4KFDZxZ9B/omU1mVAOQgMcUNY36M04a37i/cSNIpMTQL2ZUl94o0I5e/KuEl8CL/Mo+UVZQIoCG
97c/VcRSeczfPbjvgFxsvhOEA1G5om5XMlKQ0nuN2hfhTBXIPjm5Jl+qs7VSXMinWMXoK2gzJWwV
fVM0Ad8sH2WHWrpYM4q/YSCsybkF7nTwIolqe8wU0MUNJETeYj9ZKPCuO+p1qfTvUx3OEBMRFnqI
R+CqF3Fd2gxbhG8BCgtaLOiWopNG2rsdTYrykkVQVEMpJvKDv5Ka6kzPNY2NeIq82ohWlaT540LJ
76+25kEuW7ijOSPrsP3eOzyj0NuOMwNjlwQdhtD9e4TwGEvyS032u3NegcVIBFZmBSWcr3CAE8bH
JPxvKFFJLL+nBQDBGY6NOmDApci+LLXB8kV1m75il1jVkmtaJe1SmywiLFTvAVRuMCSKG3xgjAYH
ntSK1d6NOs60y8eD5LbSvZNTuCPLSxfpZnkBMy7EoClhzYsbJ71JeeJSTbBpUviIl1voFR2maIXR
8PYLSDKJ4/Qz/98HwLlN8k0nStEp0gQ+0gSk+llHUlnrzm8F7EGY35VyZkXuUpiGAJcIJvKXB1nI
VeS70yLnpvzv9Sm+1aR6PzI9ORou7OONjUuj6OMmK68wefd90nm47DrRirK1qGFfPslULhOZOMoF
FunqV6ZmytPqNpwqwgOHJSdUwDZrcvUs+Yx6UZEJxkbdUlMtm8MmFXMx5jZJs6/MfKegK1WxOCyK
xdrQKGeFeeVgFXVQ8aiLc7w9y9ZC3ai/qrQjPFlh1Czwk0hDT0jFgv4WDBszBOrUV7P63B2jEvm6
JwrdZweRnObqFddanZtKnvcyzSWeqFjs4US2psJDzkPDSREUjTLDZwY/br682hiOVx5LGgG3AUoI
v2utz07fUT4CzGvORxrPDf8T1nPzVwh6KdNvtcvh6exZ4X4pZ/D/1MEOWb1pXadtbGSJPDHjyn2D
91eykpLe4yA8e6+CEmjNtrhrDnVopXoSEJWzdzyuAoxl55tesVk0aWMK2+82eKGvOXnyIeDgApsj
CJJ6tpP6Ei0uNro5E0vwKCzujnDxlZXNp28VHgw2BKA3y8IWbChs8s1+nbrs6LUQANMwrQaqnuvw
IvrJ4Ox+xxqn9uqPha7nlBod7BwAhSBSDxECZj8yAh2E/gtdslLGvYK06yynD4R/zunVCWtdk75O
DOM+5B/QftqNSM1jo5PUFMQezLHezegj+yy3GkRW58LH94iTqXZwe4lbWCSCYBG6Zq9vHhqRb3JD
DklG6DN1K4zH1CFhsOgHZGPbHzPABsYZoKzrclx7Phene8rheF3+7IFFj0gQThG9s0BsWMG0WT0e
0tMNaWeAcHMAI1W+32mpwUMhxcd0szR8s7OEHyoKISlZhy1LsUc9dhyxpVx9WYlyiXdkdxeEbGTV
ux8TCiEI6QvarMAkxNGMcMl0vbPePRcMuLw9uaUj9b0HUTwSwz2AKY9iEt9zLi4mrn6Stm6h2HoZ
OJohcnL9HKlOECFak3wjkvNLnqwSWGWRUaW4h8NEJ+ZOXZNEoDWGbwKvJVofh4eoXLP++u/NP/TK
zQmax16+zwtR0fwSgQkevJDH5jFTDAcZ28VvpAoky3jjHjrnhTyIDZDNTlbYGVISQgcuGLOEbONh
0oXYqs1t9brOS2haSO8WO/Iup4LQK0jTY3TmBaaAy21IE9+F/PCREWgI33d+bq5n6gzMe6mngMoP
/NNTgo/1dnSd3xzjCiMlwfxwLCyGVuL2SQvolu12kwo+jYYWGI5TgyRmtXeAkVhUW6Ixl+5KwdoH
k2k7aUkMhvvNJxUxUfA0UZtsukLzB30Yo4BQj6dJWfIBg2r55iIao6PIngdUQO9jOhCoi34R9ROo
zfA7FG6Oyo66cGEPZJ9bhJ0rAVbaEFu6rphH2SiCfSPDQdpUiima4cscwpzzVimt/WrI43eT/hPV
SlhnLP7a5/JhaxO5XaX17lczxcejrKp5qe8bcLlLV+4PtzN4ruVKxOm7ObRfku5u8c4YTUsk0ett
blnhD+KSaXy5x9dnoNkWooL/EAyQJYrWBDLz/1kgqdwkD0qsmtxn2IgfyXTdyR6NjhPUxvzF7TfD
1Iv0cCndVcAQAFoYBbyCuLgmOlsmb/VSsNcKtivZsF41/l3a5qlscy0jSvOlowp5qsiJmICLj+5v
ce0HP1pkgxt482TSzODVE5HN8dd8VvTnySR+nmvnruLA0Vh6S78iHEV0375J4D9qQTcamj22zPrk
/Y7xf8sTSJ08X3PIVHs1M+Lyln2RTiUPlHOMQY8FtzpZCR0KsgoLJp2JHyX6qwTISdS1QV6gvwAK
QSTe5Ir8vuyXgYILAa52CC3IZVwy/XDxGzj01eUugVV/90BdEdYR8WhWrQuUqtIvNdLsAyj2NDIx
AwEG40YqD/leANZ/JPSNN9L7KaHxxQl+vK0IGlFdTsI2G8KjokN5/lJ7ORFnZtfF0KL1FVPBQ7Hu
3OfRPt7BoDKQZOyE7M7Y2bY9yFNlkro/zedZevZ55wDLu/Vv6gg5aq+sgS97O75wv/bkZJMQyQr6
q/g3e6x14vn0iIm4zMJbX1yblpeONdrm1xRbUuHPqdcKgoUw09BoTHOlmcmzVqKUdIC1aXwa1yMG
qCITwcMY32KJllDgIR1XOhD0UlVUQRyP2upTGiyvTymmiCPYa4s5piVeUkjROJAPFhUC8LXcULBz
BFElGX6B9nX20mmBLqHkbxAhITtOUiH1Qf94LjTE4AFGmTxPU16GAAN1fVJmchGFpHvycMtFfZb+
3FGkHp39D/itES6aiw991ACz/us/szuBUX6jlWS7cDyUyOm1FelldhlRvOwoE4yjEGStXTXjZbUA
MyCJ+P8IBLxmWhZoUv8ezeEqvhDpt4Puoqn5PlmcIWCyHYUcSOdvnDZiIRLWatLHKFyCTarCICsi
ZCjd7Ha+f6JnrdDTzxSpo1Xc3t7Z0llD2UZ4KaV45mW19yj3BuY0/m3KFN/xZh4OuBkNTEheG4gK
kGVxmn/gcyHqPwniyfdrmcUWCdgrQicf7iSMKzPL0Y5StDoKcC2EzDqiENfWc24h2B3D+fhKFc+j
a+QVDbMsZNLpAn8c4GXMHz+VUF1wL6B0LrpKyJG7jL8hb2LoP6hgB75EyWnnOkcUZY+kkzUsk+JL
5iWaf1iqAOXLFiK1aZv5qTcEl5pAs5VfsbXyb4EC+clJk4ZkDrOmNp3/uDMDMjGSG4Udjq2zNza/
bZBy3NS0KqTzLGkXbIWH6OcuwS73Q5yqLlxK3MAz4RS7g1VImLGYQWoqoSKvGyoVOdMTb/EWQkcU
x0vmJBJkli2cA8SZZGWdglW6xTsmBuk6btaA5uiuMOv+zHfBhbqKrHG0lx8uuftBua+/B89C+6lj
VGL9I+Aq64M8bx4Rl2YMcOUa49aSojudKl0Q7oRzM7MiYROqjBXeGUUIEaiS+2WvxfqkyEqIigbJ
jXZaNVluC095jHf45MPL1zh1ubgGEArEl5H3Cdd7W2uocGHmRm8Ym4hVIwahjtw0EPTh5oLhIIh1
ID9RGg74ykmFpmXfpZueZ6SAURlr6yLpPoCA/YJAULPhXeC97TAd7/6hpMzWqco5BTg3MzX894mo
7AbIQrkQfsHoOnd6iAhU711KTCVRiYX+9hSRz3koIktKpd7uxO9QkcbkZ28Z0xuFt20HvT+rJ+7I
HNr+bufIzhnOAb0VlHkiwiD6KiAIz9bl0k4xWXx1BefxMPb/PKHrG7sEtZqHIqIiCTCeKzpkfm+0
U1doMZ0qharv6BYTUVPlf/Y7IVJ5psn6XbsBGd0Jo8AmIBb9tTbizF+JdPyZ5vYAmPLNnTkleu4o
oGPEgKRUJ8Af9Z7Z5QfbzZfoysDAiMGKd+N2YETJSay3sr3o4bA7V2m/XWlgm4HeK70e4WbLj2ko
/jfdDT4y7wXYW+sjUu1VzVpnWXknKhYBaNa4vJv8jTSjZQaTxN0558TsQ+ywvQkCOx/44Vd2lh7q
bh8JsQMV48cezRPrEvIrQjaQe6+lHfXZBufI3iMD6xAoz5KBICMiajU/ipo3aySxxm+gqixsfITd
f2eSwv99UPvL54N5VScX0fBCjpKkwyxJz2Xv41bipjO8GmfHzXOcaJBDvsglQInMimBUa9+jTrZr
jlqy/KjK864W2Ly7LJGh6JGb5J/jfZFe76zi3G36/mtuaAZGiJXIomVt7xu8joidZPE0hWY/eXvU
khw2QlDXJV7AQRsIWDVfBKMFAviuOtgQbn5TynNLjTOiN7x1tnqlDvpk8vV5Fqvb9WB1Fv9Y+cL+
VhT3PK/UbOuMoC4RZYa5ETRfLnTC1DdHA0PWzE/5eQAurA0PD0YxSP5t51TRi1ldgu+miYT0j7X6
euiUyhGNYIc3v8MKYaZitp1zcv+ZxNKx/6IRsoLTEi2bJ8S/4ss22tpdGGcDfx7AFBJ2u9ofhxAu
pyHKFJN7fbxkXi45XMo9q57+zICRObMZLme7lmxsTszWxHouwQaRc2nb5MLioIiptclZ6S+uOBGT
9xLVLoGs6w+2ZV81J8N/GdOgYaFuG0p9mB5nttR2Rz+48ZRBe+jV8SaePLvpDdwnHPxkR+yoeEh3
VX/LFutxn/hN86MhKWqxxRihfvDjFTzRqL2rHhWypQynhp46JSiGMqJ97fxpnT9laXMrW2GZiK13
VvV/I7sQJjQRhhRroRtf5KS6+NANscBVqxzwOcCLQwr8qXC/Jrb3h9EY34Dmpp5xeY1HGLbBATQg
W8R2YcQS/J7jXb2f3OD4tszW3NeVvcTRmL2n8F9cpDrl8zdQTqYL89CXuMMn54+Xm2XNAhoNCIbJ
7FY4WWF4GFvVxQeh5bFPe0e6YJAqu6NTZgMZ2zzXHvspv3ciwc9M36StPFSZmCwXbv08a5B4mtm8
EkWY7YPNw3vEhid8b6v/cqiXILvg9pVPMByKRDpZhubrLSo7a8Fg4aVPVixaTb72xvuluR/krKH9
Z3pu3wjUhY6aEFbDeyWadokQiL/P24LQ8St3E8TeqWlFG9FYanPFZYnvUAS51u1P2scrIGdklhwt
1VyyIuVps5lAQMn+oP+Tms4wafyzUTVdKQ3twjLP6dgUJ0y3HtN9mRAlw4qHD9IGdwWwNK2Gd98l
2dypu82aLLKUK0MnhXnoHMQAEjxGyCsDmwxHYX/V3auLN1FTsK7YAFcCX4odKAgdZvIGgHjDCnB8
NBK1doNsHC7gNltDLFUp2lW4yUkyVX4jBabzr7gtstFm762PzP+ILvfbA36Sd6se1NXZdMZja/xg
+yzCLVumhBzsyTdS9UGUUX1vhJW7/TaYV7432ZYyFVN/dXWv9OffvghBbpucA1At9bNgtnIR7IIH
NHiryhUiIB0FliMEYlqr4W/ZdXY8ZHqluUR2F3vTRAEyTJhO/wdvFsJPbegFMvzdKdTr01mSJjMl
jxpw71YDtJlvx7P9Bgzl5vzUdpucDv/M9K57hGgXxi81r+LYCI7BBh8Oe1ztsCQTscj7Z/eEqIG4
lYMBRGrJ0W7Q1Be37ikgpFd7ZRf3o4wpGtYrCn03HtutXSE+6VEg+mcUZuv3J9fhy3MJYodJamNS
+oG7LsQJx0GplJ6iG1oqQ2GjL6zrKYrv1dii6hU++Na94hZ1EV+g1ElXjt/jJBJ+WoDqF5kx7fd0
pHgKrs8Msa2NTTrSLfGJmogwd4oPmFxsP+9s+m2K7bOmcZVbi+sN8rkjSxbDfvXFyJzKgcR0A4vu
uJ9hbsDteSJjTZTaP16dY/63HbeQS1pRMST1oFkQAUxbP28wv3DHu3hKRoXCs5WLo7obpF5YOTMK
N3LXH53ePEp8MQXgQ5nERlrE+6KKRVnwgwwIhJeBGR1sAHjFBnFvIFsUsqwa292hu4GFlXwVXhrb
exLrOmp4Qzp//vB3lIb1uygkrJJelEgEUN6rfESVLcvG3z0XzMoMS/h82og0/h4eNVdzzH/5bJp+
WouXPQyTUXxO32ZnXzI/nDypz3heL8y7h+iO/1jRK9xAY9CKGjkZUfBdy86V6oyUzlyAAas1KWyv
+2tDac17DQNM43XZxZHYm45e09QuZn1A43iZK/CH4M2J5EuBl77vrMJzFb1tDth3WvUd1Vhjga1B
1edSYC8pbcw//Uwtyf73bq3Q2biQ9LUSaqxc0MczsYPAhX7z3IxdxYT5ey5mSdiexKO+pQWzlV9M
absjOeH0Dm56VAEU1AaHprI+Mi5hyHqJFiVhfsN/SpGEEgxQebdPt1US1stn8GfjgPYWiJWjAqds
iWsTQEaP1N0PyXVHqIIpsUOpo3rPg66Yew6Oqa6h887hvIL5HdcMIip66Pi/JrFRRB5ZFwndzHSs
JNAUNbPKZ5boJOIdIEPYDBpWDJ3aHLzKRyW8T/cdPVuUJ7qelqWpVZYEHl1HCmK5N6lkPCCA4mim
tSC01e6p9oPIq4kuA1qknFdBeJzGXdNos5yUEMCBU4VO9lJI06tNpd3/mXzzLKkRJUOJhsuL9MJB
886MIfjQNViGlxaDAoOmiDueNmaLBg6sEGjqsPl8S0dsHgWHP6YJn0ZVkLe27g2WDa36T1iXeU9W
Vyc4Yz5zzKK+sq+uxD8G7E/6n59l9KX6qdThnmguQUlnpUGnpGM9s85QJuUGnuoB7cw/R/TzEt4n
xT7gm8NtLL5dhgyQ872cqTP8WzEpKdWLol1FldEulIwfs6tj2vDHZ8pZeiBvVSlDMhrDXzAVgb6W
NoT3DxFg2+v4MJPjLrm1kHc2vU+XJlhl/pfNuV5IkThgclaLE0igK7iuoVYKd4i5ze05dujgeNm+
bkTWYrNeCMjwDuGs2Q49s4RyOY7OH5HuCWf2OWD+s212iO9JJHY8IgrJHbm3lXBjoK1Kfr6mlLMY
MpfUuizmipCSrI8phIZJgGnEK1moTiO1RiI7Aq1mh3Qy9lTvGYGmaZqBsj8QRALNfadoqZvsuRzw
Bw32ESrH/Z1IIhjtT48YPSkZCmw+bzcSFaP/JfNsc7/KTHxKDhV1Mt1x6wa+lD5trUHKbZDIUrfT
zxzwfbNWUwJmjxdQskUXX6GmTvPGK0RY60eB6MSRdTD19XOL7wcgpDkiYImcx0H2x+3m3OCVw9I9
YPxV2FiofCYKbGr2TcJhjFTTHiqKJyKaO5N/mYYJsAvGk+LvG5FlmqUuAxgztGsIMLO50CPTDjxe
g7OhNnmrLhWTR1701aEXJhjGQOb3pxYhyZYWw8gZ9O59KVchf1RwkSiQBvy30QuMnl55eXP1Z9cm
5eFbpbJ0S7aO7FU+ArMWDeO4OosiPDQmxW35uhqUdZ5dZS8AO1Vp3DGafmy6qFlR5q0y1lAyDZJ8
pzSq61eFnEny3yyWGU8wy39U7w0MLy0LN4CZkN9lDSigsaEEe4igDVttNTu2RhOl4nC8li6tqdVO
9f/slR4HJSkBfRJ4+K4xG7V5Npmri5muHpHHTMhOqXXmC48d0isgd7ooSIfvTSF9f51CsIuKLOfl
iGcQsvtXocLUiaMgHDfA0Wr6ySVbhOdKKz9P9P9cVFWgFxe1UqJbDFSZGml35tLfH4fTSE9LOL6j
3RWydX1j6uRpL7Uw6pp0qsNkDf0t+8dFoZ9dFH3Uj+fD99khnlTEBV0wZtJCtpak83pFs+NLcao9
LZL2veeikFjfgo4gA7oouY93kX0slYfYw+SKW7W3nreiujePJt+XHOKdSdeaSOCesSZjrkQGSncE
QvzZ7/YATDr9z+2a+4yP7nNJXv0o091WfFz65kTaBkJQ9TZW3YtasJGlMCOXVxQWwBHaoM5861BN
G+j8pEq90CTdB1dB/C3Pg0IXf25Dq8NQbf/zbcOtxLgKATpBLOVh7V/nTHLR8vVVK/sGR+KGFYD5
1tG6q3mgxY8spfPSP8Y7fPk3G/EI/JveqS5vwu/aWyPA23hCYmbvfzELIcbrKtEGrnVSwROUad4M
ZIaN5DvTiwOcU9fOi5CdKHFeyjr+xeQGarMtif1ahgpacOWMzkq6/sJyTAHdRGwSM6WSEtIYO/x8
6PLqA9PrOTsjNltz6xSnIWBwSnSdAsgRYopBdkaDARKxweiKf79PrOZpMNhQayyxASJpIFc2bnBm
AzAx1BU2U+7PpR+G0xAbqShihlNBk2fTI05MnzPxHIy+sTD9vHZQnJ/4wo9tYUZP8y2ghrv6UIFL
qhWdmwlXwuJr9wJOt0bVuqEjHjKFcLjoeuQORfpk279GgNIMHEuedDs+fEWw9vfMUGCdSs+jzc88
miluxkO9AI91I0+Ew9dkOy4BBXFYxQipJ+fBc9/DaakJ7KmIqX8RAXuDe3lKZ3DQlOLildMiRe8F
wIQ76R2GFUBJRzIDL7CLjrhjOkki47KIJO5czSHokZyjNs/pjJSS4k9ZgmIIvYwYOt7xVbfO2noT
o8pjWqwttLo5z4PTaJaabbcpNdm0Zb1mDfRv39+lefBnaxGQNfeK4Lg/QeInDYxH5LU3hC3zXrz1
G5q9HBB89gXaedvdX0DbuR0iFYg3XxK4dBT9TkJ7GoI3tUzYV3u30bg4iwAJJFtMVOIXjjKoDDGh
fIxod+FK+kQc39l6VOasTokCTyjtxpJ4fYe/CvY85fIg7f6LWfafTjphlrCYGaZB0jgBFhTEvirb
lUs980an9DIkBFF6O/Oz9TdZezbvsJXxuTas6dBRRrzLwow0xZ/wTdVkDWPGXrE9NVfts8EYuI49
08wkk+XSDD+iUGbTXowvHp9GdQ6gDKPAvhPM6wgDk4C9zeaxGgmk9hSAS/D0kkbSJKCG9aW1P6mp
5Z0icngl6FfRUiKeoq4BfsfYCNOLKEsXH8i8pXQmt2j3yanFnpzo8QmrGt1lSA4SGhvwgrNQ2p2i
IuY9ToidCrOZDnNz1KC5t6F0/N+eooZ6WSlASMXxw4ttAh4ylw1njVF9nscJNczfJ5tQ8wx4oBRA
9+4qtEmP0iaA+VMLnHowtKO4h4QWhHixDTbL6D94s9W4Q2CHaZvjBwvlqKU2dER8Hm29NVxrvSed
KyobANeW1fMUEwU40c8tExd+TlIjWA5Hseik5dSIPjbMX+yhw+tUcHQCHL9TCaQc4jpMhanmBQeM
lQgYaQSbQkMO3O0yPT6uPJDm38zgQaxmQf7LcKT8aERXpUwVu+7s1RQnHXAe5Xo5PNfsYd3BE/0j
KVZcV/+f07bI0bwqGV/Lw2siIXjHfujTlLKyuAp/jcdVOpV4cgmmU/l0Mw+JJbvJ0p6AjAq5bTOb
6GMl9rCCXOTomhJ5EHuQ1GXrbPGHdSbFoPTsNrS4yxynWlLg5Vj1CGPx8x/P2GPc7tKS+ceEkfYG
ZWO9qtHh1JErGcNV/YEx8DBfmCxdfpg90TeNqNfHcAkd/+ngkYyE4u1imD74PCoijMgV64mTAdbe
hpoiUN2+3+JDV81vZ3ADYqKVSFobBzFl/UoGc2Q7QlKhpfz5vKjUifmXh8LS3/3plkG2VrVDb9ud
W9EqQxjmee1f31pv/+sWbOwa4jHzehWOuqssdVblXxfxjn508WbtTk3zFDNa4t8uwyRvMh2gy08G
UTrl/rrQ6qGWjMyGZc+8Y6euJKyO2wSrcam/Thms+qhzgtVZ2ZducxduJb3vqJgL34Mr2JSvpUZ9
3FeX8ruaaBrGS8PMcCxvvZZzZGhMNsaHmPh+uEOQf9I714VpvTkXdkjF8WE+yR/GZfCvCUw2/Dgi
Sb5Ov/DqWHxKVX5nzfJlxKeL4hzuw7/7rJ7MjYQnG6PprodFOtD2LPyAjGE936NmrLiWJV3XekW7
P+OgoJM8/6wVoYGAaI/7NtwTBNmK89Lh3cX1MERXkp16Jc1Vmc+zlXoem+VXRmxsWxw+yRSfg7UW
PfW5cTMqyumw9fn81OIGolfy4dIVuLuaa6MAtX63EAmdGOGvtpHHmzf0S7PM4r49/GjRAnO1zbtE
kiffjNWoGEgW1DavniaG/M51KrhvRiTWxluraXRQvbUXut24TZ3oVzx3MqBMdGrfWVUDJPtIOllq
B8YT5XhnW4hcOsnmJRG3FvWsKBg5E5O4gZe0iYipe4cs1sGjD41mSabS9yw0b4kqXXpNpnKHTqa9
kF7idQ34F25fSr/JOd4wwTzFBNeVtSUIqc7ccNBWHDW6q9osjjlqWdZGRickq1AG+f8w5FlfrIuE
1q4x9ln+0sGJ58G1W934s+RiE47fS+Gc3TfKC33IGe05ouXe78cAn/p6KkUY2gBkcridxYnmwwkM
myYfiW7TU3yloOFdHb0MmklUjblvgWXxD1BZRpjCycvBMxM+UrNgVfAu4irmzsiY7Hxws0HW1aVm
9x9/EQ4Bh3uKOB+FlIkqYiKCBzRmICDWDnshPcV9L16y09prvhtAkeDeFU/Z8d40N6GSGTlPoNnX
rYCeOart1YVVbBJv0oF8o9qvt6HG61XtiQsLUBKCmYSH+yFEJxqb3bmr96lvZ1Z1h4jEqbWENnoe
Y8CDpM/RKadqhadgcti0OdlyPQGWrJMop557KRXCcAicCUBU/9r32r9AWaEI8XVY3NqG8MjpbuII
3Y3fvPlOICFgf3J+cxOSSaE+qPOInOiYHm/9JksAPgGEaXn4XnuQHhMT+7MfAnwfBAS2Ay76J+oy
HqtNZyx9wMZi9/CpvkOUfClh3035MSmcQfdviPOnhYPCEAh9ArlXmVpEHAw9EUKeP1kaXlBSFQtj
TMLF4Iv+L4csGJUB7eoEmR+Xy+CpNzeNi6u7YtYgW5SbnxTnYmLd/GLtNJgEOM6P/rwEdfZZ12hL
vqONz2K9hOZntwSG7qePBN81TSWWYx3215pzAtKDjFPG7T2er3O9P2d3GNXWCWPNRtbq12/gfG5j
Ujwe9qgRVLSGhRiLRGYoyGaMI5UAc50VPPRb8+ux1TCoy69/sVmfltTFfRPPDrsMzYsFhgmgtEOZ
od/hTpwgWF8D2MmjFa/UoamFup4qWSwSfQQQpg+pPvh2ZfFFTjWWeZsWd/jiZOVg31lh14FK5sRq
XHC/0WLEy8MrPx6S3MS+4cLkiCs4kukndLtGf6m/o6MLA4EifFvPlgdBuqq6UKIo0+QtR+iH7fVU
T4d3JIYGP0DhIychGO+StkjiO4+3AzoS7T74Bv+Jlog7qKfP+L50K6+vhHpWZqjimCNl+nkhHXFi
5wrK66+zZG7ts/7h+bZh2A+gTF8Q2RZ8BAt5KpIIxsTTYHXXe2r9EzagnI4GX3RvgwKQKkQU0AUy
/KN+f8fYnhmVmIZfmDK+u3mS7FJf6F8z0BnkQanqBXExN7+1LQEAyKbvEpofcUvcI8w+H6QZLpET
hQEo25TL0urtnsmsEV9JDlN2F5M5ZKJl91n6eqI99w3X1Cwq1rRqndjqtULZFbTOrBWKwiY4B3Zo
JoiqHymvNBSGSCHlIgseJbHwW5DgkletS2RPf6CJ16KOXcEp0Bk0Q2IRIitMy+YdG7t0Pu6MuPaw
mQSKeu0nOcTvFLFWcPtJZ78Gy0Tw8LTB9fqZMgqRptHRazHPEmvGNnnJoC5u+pnXHcDiuwaFVgYC
/jqjuBx6tMn5Y8qzaJ05cXkUa1R21dA/sgPXXPpbQC8pyxPoFT1aah2u+sLl4cZsbSZ7QjSpmfsx
q+4MFxd34NBCXx3fGiClG0uyb86vd/4oRaz8KAmj5oxWiQyBbUMvnVf+J9ecvWLOS+ofzG8F6i02
Z+OTXWU8MLKZEGfo1mwg3Do9IasUer17IzQhLXRbAtzbgM4DjCRNGONMBeesoZQ8uX9rm9f0Dk93
5LSgKXP0twslbqS9Tg7DdHTN3QTz9rXUJClED0qt2gCldH4tZIWRcBHQerr77q5+VVdgJXzPI+Hw
OJvXW6AW5PaDlNAHR7cRVHXiiriLqPWL0zJhSvdwfZDuHF3se3Bp6Bi+WXkePMiEOQO+7yYaGyw7
3mhj7QVx05Gug2AhWaSHtQdgrVIvtFNMrkutFvQ97KGuWbzfN9TGkOW3Doqoebsy4AK0KraSI1Sr
VL7Yhk4LQsoj9RBUfN//GM+lO6GRu7zaidd0GXI15krwQzvWgiBrL+6+tHbD8Otr+V3Oh1Lh8RII
ZkX6PVjOvx08IZefEa8LcBTyJnfmQ5QZKn95MSAAY1PQh5CXX+YsS86Heg17EXXDmKLDcDfbZsgf
QRyF//XgqUtDJf2c0T75I4/AwFWMVbJOjpFfzDuGkvrFNZLxSbQiCJjdTayXTUtMyPX3dNTJFQwd
L/bgFM58Nps7iFpD1l4bw5CAhNmFXde20P6x0dczT0G4/XVJh1jaXUQ5CXSljCtVFmgsE2Y7kkkL
SfqG14gwB+zm1AghhENXWJjzYXBck4hO4jCbDvSlmy5l2QBVYRlZ8f1MpkxCefyICZLdYh0u3VEY
h0pKfd1QDMgfI8iXsQHhxDP04QJqYBK91EpaO6EiM+Hi7G/jocQmUqSCjiBlWjx5KGgBh+hAqilL
QTVwK9yHuqigooHBzLEjnmHahugZIkdWvuSp4dy+BLMWqCMd98iSRB+zLozV/Wx04gXWnVPhMpM3
UOnDlgfEQcjzzwZwLWfeAFpQ9PsGQbQ3ypObdFDx7n7lBtCabRtHHwINTkwAaLQ/eBPuqpOOcGBr
eVgAJeE3hLp+V7jBjD8HKO3hFpeLAC0J1JntPZUBvNqIKj52C14hpt2vv2h957dUx71nNxUyx0cY
yz2kObEMXzBp8WtAm5/7YypuWGjs5M4/ISVhM3nxiFIC/cYTfmhd0iet1YydPF7AE0VpYAxt8pEN
mKp9IJqmKpX5nZtOzNSjmyhJD+hnAUZf/8joecmFfdyp3DhD+yhqJHndUZQekwvN+UNPDFRM0+eQ
X0JEY+VnHa371wU2TjIpcrSCiE9ruVQc5WKe/jvzvkcpgiuJa3+ETxQNMtKSxbR20irDQ7kNp5z9
a1Pc3jK8rPQzKC1InPzdKgOJkfWjdejP3WTQRC8f5FVIhwU5kpEfKJ5pJp36F171nIhGq01t6hmp
IXws1SSI2ejJHBueuCikjQo0OyzoThcQixgu3ZKOQLI9USI0pDYsQQPVuCXuVqnv5/yHYB//8PpX
1dVnmZZzKGGn3m0exr8FTtBYODEvZaNfn0n1Gr0QK8+VXHyUh34uCZs4ZTSwmwTovvBkvG7JUnaY
4FAQlHNgVzfaNkA6RnKDDcPKdyjR8BtDLII9Iui9uaoNMIoBZEvR7q7hzpO4uR69Ba3yoc3rikjq
q7posflkWE9nCi4HeMunJFeL5MP5S2WweyEGtlc36vRced1zYtY27DkRSNTh1YBXykcvPjKKLqNz
hnu/MhMp64F3ZDSZJ9M69ieevdOtOidPaL7HlEkOvGlzCQ4MCT81WdcJDkgeMx6+3AS2KPltVh9e
YDaJsd2UE7MEExG/9JuDa+MqcWt4CkBWNS/WPQ2G0/mQqY7ocU0JoOtvXSYf2+awTW6Z2h5kicW4
tupyrowCjKD+2zCMGKbBX69rwf1dUXTn9SxIH8Pr0iE6mt+Xvs9aDgupZxlb2hdQoc5xwd/5J84B
qaQ4gDxiyddrvyrTjsxUSPvnxJpRZY00SnvlG7+Zv0S4sTej7gWOrgKBeXQMVC9DW8FzCeGadtbs
Y9EH3RwZOxyGEwJ3LqXIXF/kYrDZFX5AXNx05kiIWUwvwhtahd3bmnec2HN2hlRI3vLPsyWiHbRf
fqrFUJyPAEt8jNYyWMXW15/6tJSr4iNPRaSVXkfEfY/amsKk8ws4Y5DV5LHSMCENxEGtlkccxvmK
gMxjQIROK9GNYrKg0oPfQSpUsaMHUaAWVS8zwJbKg+kZ02RsujhMbZXsz277LiCV+/d6+musF4FM
RGiXOJ8/FjTQf4UCRPXSBG7JsSNSJIO4ITS3ZO+R9uAI2iUCamqZsvJywUeUCUYahnebo3P+D+Lc
8cz2IP3wPaxSzD2aKNttQ9J5s8mFVIah/wBWgqAoU7OqtqnGN9JjL8sg6v5vslxvDvHWlAX9kHo1
v18BVs7gd55s/yz5bkpIsxQoRz/+uVTcCYw1D8koXYEJ34QyYk5Uf1ojjwzPF6ZqmIAR59ktZBu6
hpVNmuo5bw64RN0uVA9bm6xCx6eXhHyXm2u7gsvqevqBQjIv2ezwGGg0l+sjAGClTpR0YnGCid47
n3b2OHRSC9tVgOSX5esktXDnblZT5I/CqxqtDbwNeDXvWrTksUcC3BdyvXI2YhvBJdgy4goO1uiJ
Z2jucjhMW5wy80KFBGckhSqoeiA9tMWcraSfxb4In45cfgxqI5e++PXHzc98kmL+qvEyHfjdnFIv
03KmSfzbctbtjmkavQDOXPy3bVju/7VG5CtVrHPl84jwYj81dduABgk4/ucfj8F6axnQ6ok4hwgj
NShp6abfwBJLGqqjXBmDApyIRY7SRWzm2AGB9XpEYWV3rIrL4wTZ0l4+JdGER/BuXSJTs8E5uCGu
bqx7nXehsd6DV0OeHx/P05VfgQ3s1aLXDwFCgcmpYSbtv5lVqjqGrKOzVr/ROgO0z9/GBWbkziDG
f/CI93LPcbCWCp9rmCEl6zjUCXjYITQ/tBX4PPp/x4EQc4O0zbd+ETfxwE6LVZgPmiTZO3cdiBuV
e3p4+A6/hVM9GxO4m9ctdj2ve899U+wJ7P1RtBPkQs6WDQ+uLBxTb1RcatMpQV2uJ2AAlcBlP3hb
5d3wkwGC+YA0HdT6d4aUAYeD8h9j+pl9DGCVwyfcin9RR427XLlRPaBSijOlWNaVPYdBHaWlnkgc
v2b5d07jKEtbkPa2moAg7lp1j4PUlpXyUq3aSfe7wcf0XmvDy9d0xfCn/mAub8KEqaDBYz/YR2xf
llA9MNuBO9c4PGaTMTwGU3i0dzEKs4Kjss/QBh9Gl702ltlA1Hh08jXw81ymYJfMBuZib0vMnCxV
Mvo8cxb48xLLVI3JJ7hYQG8XlHkt9kmfN8AeRmKOujoqIVXf+6ixD2EIi/jOJbRMDbpI1N4tP8fh
6YFYaIHKngsdCbKzBdBxGX8mB8bdvhaZX1JSZYW2Bz6Qq2oGTSuezVSm7aaY7a2kGFfbFC0rMCyR
2AbZS+lqVCk1pUVAhyaqPcrlzsYLSEWTAMq2W1gcNSs0mS3dd05yVouq2y1/XWzRbOeEeT5PGehk
HVsMh9yqjca92PHz87gWLVTGBSEyQZOmGcaKLTegK9ZcAHU2ScgkAhuQrcyNQ8wJsJEyZB/AUv2D
mHZxCzuEfj3nDNTq/8POqJ26RMyPKeYplzpFo+bfoJWDhV2ne/lGCZQ6VDHYcrMMeUGBx+G8rZk2
bY4z2Rfsb9Wde0XobGyA5aDTpHAkMCIlK8iYVpG50cqkjpDAGuoEJi7+aY9TlYHSFRdvDFbobSnR
jiNZNVU3pj6HGyGW4+pRI8Ou3SYuz5K2f2LDq2Q/vn/hwDN91z+TudiiNhooQxpCf+0yONz7C1Am
SoaBOAms0iW6YMaV3oL+lFpM9qVZV/dm+6K65JpV1kG/BkaSlQcxk0kPn/7Dh/rMhdenjf06CmfK
u+rJZFukJt+rWjNEcS42sGgKQT0MUMPoXN7CGTAjd5kcYYVRAsKR8L/eiLp3Zjf1DYEw/AexPtLB
EcTrIBR/QO03d+xNTZwIRFYdP318S+XMuiHGg2Hz1Lbti0wMJPBhwTVQD0Et46OsODkniy5SfyxZ
Q+pm9fUCvpvALsGrSFaMSAjii0unqOex44vQ2kp3F2Rf9AbWIgd0RcL9H354Pamd/fFD0wGXrJ36
XgDuvAtufSo5BpHsi1ufjbbgLujnxHfvOSpHuI/40HePP/DwQHtcMOWDqXFHJirstOOaxHGa6R56
5axy4fpiMjjv0Lz00yITpbD1SRkX/Y9YA6qiTljDaSEpvyAgluclC/zSWBYLz05jSuooq5h0M7w/
OI5Tv2PAyk+2FDw8EzND2IIQ8eP8kxfkgCAl29C64p6snWpKYGF99IaqDrrPNpu7eK99A0eMesqL
9heatDpQjupGXVJm92bHT5ha77SFtdVVEWBRfsyGDpej5p9zGj4vARoEzeVtWG5/a9n5+YHl1fxp
+u+gMKqbt+B2wrmyVXKWH8adTPDvTJrECpM3cLouqE/YVmolgWeXJU57CV/64C9dfmeCZorfizee
QewnH54jXWF+BEK1tFb6DWjyN4uwtZX0spUAFPUC53SgYTzSOrDnoN9TfHs+ejfxewz/ND1QRO6H
tkMGc7s/hlTIcUqzt3NwXS+5WchtZ/OO5nCY/UmDnQMsbWL0EPBmVlE8ePWRhQkTjrhMC1nSW2ek
Gz8XkXW79E+4LwUZ/Xh8XWoRAIPRUZqZSiiItZYok/gOi5qDz8bt3JXbi+5x24hT66JZar9a3y39
Sz3win35jLHeH6UUkAy2p7HdPm6OZBDNit2pWtSP63a1Q9jV/GR2WKKQVzQVseldoWYPUo2CFjUn
RwHKCFpJ8d/VhlUDeJFme9liIvns9LmvVMfK7e378eQ9P6tFfOQh9BuyoOmbaeliNv+Dj5QI4dKw
N3K96pfFb90s/lQ9MGQAZ5yB2BmCczYv4Qg74DZSDfO0orndTpMqn34+aXw8KeTDqb6zpSEtC/Ea
LCaJp+Qpsanj+XGjalo7qJNhq5fHziIPoh3nHz/3fDXYzfrHZXh+sLfegTXckpAuZIfpyN+VA0eW
Xcnxr8oKc6O6Jdahl0DA1IYBqxcuEZWP0TUhxVCnTJHnQXJTLO2i826iMloyYmIdbxgV5REOohcs
URTMmBvo8FsD9GcbvFaDLzg7Sa4xy6dscDyEo5rZKDhVVQQu2It/0vdbSUedAyCQ51ONqIBEzgDH
/94Lp7SEHu2AVE8h0vz1Iq5fTaY+/SjIhkuUQwsRaJvis5L3ijuhuD5GuvpNYRslxf9qZBGe+BeK
HOzqmfk/G18Zpiv/RPgq3SXT7wHQkFO+eOfd5H1h3SP0Ek1uMqAgcnNlNQUBKqhGOwjtlYnMW3EC
80ZUKRMDRstO7opP3xpCJ8wffvz5222QZ3F6Z2/jDi/NZ1RTl5LBMZ/PgNJZo11L/tSYuMNKpFT1
lagWLFIbKS+6FSGgMEQCZfFV7O/9wCEQbhlfpaxksIe/5cFeRGU1SMG6+I2nG1du8TsMiXlyQ9bQ
CCM1KoWgP7gSUW3icyrKLRI9FTzDyio53uyXfQtvP1Pk7bU2LFW2NhRfdIIp+ucL+UdEBmW2H6/N
gQHPq/24bRol35qFslU4vIaLYjl7tXeU//hZ31oNkgisGhOeUjUXsGvqJS4qZeaLJ2zKtKwujWjj
hCyxBB622IqgwhxCXl8rtuz7PrCEZSLCodXdD9Vo+9+jj3FXamMWzst3f7pKCdzeTM6KB3D6MGZR
EX3Q58U/FnmCyd1knkGYBBbR8n3SVjKBB789s50s8l0BNBjgOS1VWwZUA/bSMC1qWO8RRAZmtwHT
fQra8jklm5Fm6LuBxDrNYn0surnJG/aOQVuW/fwAIFib2M9kB4DN7H83jsQVHtKplyoHOCzy2cNZ
kHjp8Q+Xc2Mv1ll8xcg5MHssx3AdPiiHGyA6a4rVRIZQsxD9oG1XGEk4mO0RiJaoBPh7FoVezwCF
MvllK0M50yGfOu9PsnKFYklzVkNfeysX576vXLCOWm/FrUbYjbwXDXOt+8V5tYKc6tkd1wm7YPKk
RPtcKtirQvjutmCbssKEgzt/9Ba2Rgfni/BKP4QhUtpzi/x5Hh0wvwdr1LeR7H25Jyw8ehszzAdD
IucZWAXOs5PJ7xdsGpn3ZiqpAwU382Ny7t20uUvmrrvJTbrtlFrsYlBo3Zq1Yxo5ry1qoIUcvn5Y
szSWziu+lEMVdsxoUlMp23L9GEehQ+ffB23Ju8JYy/8GTVHF2hquTnx0nZv+97ED8pRPA/Z0qH+/
260/jY550zGWrssxqgR1a43xKgRdab3o/RZp1W1NX5zSj8dVAJT2zcCga4K0xdEQz3inUvEYXzVT
QtyGSij7x7g90Qbg9lkjMnU4pLQ9KKzymA524PjEEzEiWDM7RnWMjTuk3UHsNiyEEg1paMFgLUy6
/aBoeJEvmEQDfhKDkaseTifuKShOER8HfUEamEo7MICg1BG3VTeZj+0N4lV61ypjeLzAKyWjqAHJ
sNOhc+qcot+q+Kcqfr+Hgei8s3HQFikIsz8kG0khJgCOvpM2XZq9TNEjvJ/moaDRNE1KK4O/sLMx
qImMKN1wXxZW3EVoYAReRkRty+lUp22lTkVXC2SiPyEZ4417ySMiloW9gYOPRi+YPd4L4Myo9DXN
a9P3Gl4zsxpuxFh5wqYtgKqnU6mluRHR4U9vjTbXOC6V6bitV0rnUhRcDA0eCegYiSop5xWnXtTx
XwFSVpeUjd6C9Q0qy3EmDKaEtC+zvHZAfniZEg3akoCTcdWb+f4vnfQ+BEX7ZUzl+65MZAPBqO6b
KydQiyCdmTNa3No/sDxEdfxOi8KQU6adeFQSvc1gGu6nm159kZb0UbMBbsAbLRohPLl7YCCcxiAC
7w6Bb9pYuAc3McyMf8CnFOFTA1ZfbkU+IS0vCVK+B5/241pL2Fv2KsQJ/dGRCl9TD3fCaPl8J7hY
hTsVyh2Z//JLyuJaoma4ibmojM0u1ozEM3tKXsskNu9A7+o0EjN4R3WOIAG1CLov7NwFpJTzv1sx
3RXG3hcpN8b+wUK2p2HKHLtM/ixOQ5HDqR8fgsf3gQbzeKowEx6xc7h0J3IHHyM+HKN6idIb1H8b
TBoTOM2uVcaSQRAeI5/J5UwVLwd3vNdbaLnPFUXB9qtq4MIqQvWbwntru4rXH7npErdRjL83ifSQ
QzHNh/fRfZvy+236zWTPKfO3HWX2RaibDkR3GL9jkT3S7529Pduze2NhqJ5ngmXR8stvww9yYQar
YTuOXSVhqe/z9DTm1uH1yVaQ4LBYzZAMLNGVWoQRQZbVAiPt6AnzAZuMYezaUv5cQXXi+Ta37r+V
LkF53Z1WIuwuGdsZjoF6/8BGSn3oxhhTCNnpm50gRg9YE/EnUV3cholgQmHzjA9T2vrMYKA/H6Sr
/INawXQ9d+LgIXg9CuUwl6mDTzqyv/xpzrxX2y/vnIazfoeETpMti01m7blmPKZrFbyGlVi/DBMs
3X+cz24OVt+dd4/vGg7uZkr/8fNo+x9BXW3WRms24OfvQmJlCvP+qnN/UfhLQ3ATkQOk7HqVbcqi
97GJiKZBGkjYRb9WR9hF/AzYcfaoOBlbTKcmUr3pQpHpw0HFyeNJplmaEamezJdvPhhgVNbcR8r6
i8iupvyx77cPCCZNtixVoDojB8yQN2cBXQ+bE5pF8x7U1NV8D35lf9yeSlDJKWw5spMhh84Qm2s4
2yerhLIsGdBzY5AjCZvCvvxRSRL9WogJE9FK9ZdC280qiPqRtYYbEVpSKps3OoC6x8AzrLcJB3Q1
lBwcSa7G0KLLtxCHG3I65mGim4/cwUf3IKTg1avzEQO0CvuSKWAAElhu4HA3tXIwGob8HCaa4Ccl
n5gMh0Cg8Py1sfRCp25n4APzUFjuI5TONtv6MDSdfTZdomYMt1RseClNfuTRBIPU+pr7VavCNRoI
hAflzLOgUHdDDGPczZakxlESGCnRyHJ0bLajrfcDYW2Nfk8+HxyftSaqwbescPgPgdSU9U2GEein
X5h0Qxm5gucvePdxN3TzCS3sRyMMbQUIqnNlXXdV4bK7DU8IhYbQIYy8pfiw2wFe2YR3WKc+zXWO
KIpJIsUBoFpzGp1lwBzDMpxPBLamDckrClqEVTbNql/mdoyylVYTDN2Vjo8/T7DH6NxEBnVSSdzI
mmxTVZeNkltsJMdtdlcrjz/Rq43sMlt1xplLhnrCL9JmPkL9BQKQlZiEnuDXtCYK983uhLUnYSE8
uIVjMBgh1Pp3yvyt0awL0fEwlwn8BcK/LeQJOoydxceKJNK+WrAdHIqX7iMyj3gPwSyNLGyekEr+
vfxZ++ZtySjHzqoufZUyJ4zXObJM1W2ccpVf3mRYkAnO/b3Qu6heO6UWxLvt83ZlS6E8Emli7y5k
hP8zcnW/JL0t2x7GIAgWj2bWt9Y9okLo7VXvJZp5Yt1GGDpZ+5rModtLaz44e4wKcCKtX9p/Nmbu
1vJ4lXngMds45AhViRHg15ezUg15i/3fZUdsLPWL+RD5uuWBk4+JjnV+X/UieA9bQQ0V0UUmBose
ONcnyFJ1Huj+6WD4I868pfdGJnDICEM8Q25SWCOik12ZvX+8GnVl3RwVG+j0Upxk/EOeJ+SQ1bKA
WStfdl9642v9pntPBXFY9YwnBbxfqvXvFxgj4lybFF+XQObvyGOnz+R+vrpojJhleTwV3SQyvTgl
do69NgxUk/yM04Z0XiwCSDwSbqZkUgtihWFSKG54SztRAyr4uCAIanazpf69fTg1fP+vV99LLqy4
DoqcpPsNfb9BNFgzyhARgshrsQhssL6QcrTu4h7/PgrJmlrs5hdIgaJt8FeGBvuAjSTh8113eN6m
HGaFhIZF088cSIfvv045zH+XtFwlhIvkeTIpLcjk7i4thAsIMD/O4/xSyqKARbDey0lCpOVEf8Kn
sxozXpENlMTDbsvOz9of/FqMmT7kZWVB4BjtljZMCo65puRUmNXYHBfkfgOh5wSu0wov6aveCUYp
A0m6AVTgtFoVSSI1Wyc8FdcsXwUMNZ7rMfKZv7JKKx6TpASLYgftO5iyiRXwzE5bHNguaiBLnGXc
M7rjY+hevW8wvMIp3v4Q1E/GFbVuagQIWzT6JbyBZB0U+oAcuYiwI2I0S6p9Yjb4rfGUXFaJqApT
+wS+dr0tNLXmhQdQ+icY5ZKv0Usa5ZFlFWIUsrqOtQGvIzFWnDteksytnbXC95IQ6teBPtF9jsWM
xbvOHVaYg/Dk4x6pArcfCen2uFBdU3TYQKo6rvBqFuwjpoU31MZZ/VZw0OazqJmO8ijfPvVaU6VP
Hxrwoeha8pJ4M+9D9mKC3VdfEu63Vjb9gIh5oV5vCh6NdSg0bq75HWJANd35T7W0oKD96e98+ED/
8XUAXrORxKHBHPrYpkyDFHTPWV97tbVpfkpsgHuFEKCOuZC7APC4RcXMS36WUv9Y/LUQlQW6AK7y
o6q/Ym9lyjY0Ny8Wm1SkAvdAveNwovX7VkODRFqU+1+vZH4cZ+tChzoFYuiRG1L7PsxZk6knA7/A
CgqIvCrkntL3ZOCBQ3woFtLz0vmmCC+B6ZepsspyeVZuyj1QSiTXCyJmPb/40z+ukcof4t9JeYJ/
shNODHqczDxRaFAjIWXmv/DUpesexWEgEtf0mHDK4it4VYnaOpV4UvCr3amK6aKuZawlQYAKPZcq
X9dWeCGvufhm/v2CzYSU6R/F7D9wQXQI9ziCXJ/Ak54smP3Tt31SIn/KB/cUkQpZJ3PiiVPWCeC4
LEeljmilWY/m9N/0Dqlc9DjTAv0DyLhS3B8+INDrhyPNA9y7vbZNcNii973+nbeOaOFCI9hWEYye
jwgPbmFJ6N5xNM9jPEex1OUsYDU/kxyIGAblxJe0iAwPl1mbr3dZgYeQSnHwNBLDf4nKYeV27AaN
QiR0bTKZK5Q+lYXApWbGqMwItBtWwZyOGSO2NhKz5IZMnxnpXkh7DlfOxI/CyoUfFkzN0N2sIju8
5aeBYWrEDzVzf8Iqiir0VHthqc7xSHUehM7ObVNXJNro1Gv1h0g1IoMsJ5BzNzSfKVDL4WYccX1X
BkBfq1gu0JZFkY/1Jx61An+1GSo0toR61FptEfHVxKzklyfykfQqGkt7ly8ZOtU3jJiHqSzp/F4x
1BATa4LeCSz0s4jGI2hQinhnPzQVzgQYSkqzDNIVutyvSlmH/QZn95jluvN9h0KJjWzsO9xQJ4Ec
UigR13xJwHgUqjq3FPnX9A6Jad1kUCvIdHiO4I4wkxDe698QIlHP9H7a8MAokLqj4n0WHMqM1ig2
jdl4XrQ/ikSpWS9Gq7d78a0L6ppSSd16zAYWytI8svnLpYqq0ZfLZ3Iah0Am3KdESbqWpuKqDk9D
nDQdhSJ03y/fh4wXrkuWjV9WcrnqI1OcuRnYakVxunQAXRmSdjAwn6md31lHDQz6CXxH450et4Nu
JXMJ7yoJt5FKG+RbiEJqOFXn178rxRL+zcLj/20MnKSvf+ymPrFq1YU4PWlll4QKhZH581ZEQgPJ
VEWH1LX1aPv5oOke2EbWr1gVVUZzZqk/ITvpGqaOvikVVTn4Xbj3ljw1FyXMQ1a7fr7oamqGwk3c
sSuRVQXgG/cHBk4I3W+EeoBuHeCfhOpUUmPXlRROpsP1xdtOkJv+lTJeSkvLolLR47XZb/wxIjg8
r8Q9qxf2j2Kp4vGrUuJggm2bSd8VGTk+p3Iug5J/i1UQjUn50sb/HRMb75kkumdNeVxRcpKn51ei
73hOtmUn+s+VSBl4cJu/jxiWsIjt6yoA9+6ZNW9F9lGeX+GHV1jYriR0aWw4kBRuWn3Ze+HK/IuD
qlOg7xrNTazS4jCj+NYFpFio1FihGcAvwOIQkiD3SXivvL6N14QcODP6B74F9h/vLFalV+iDHL2U
9xjdc5TWQbTAGF/pRP1RC6DNGsqGLIWlWmS68l5f8RGfuKgVe3dqEq3J39s/MhG3taf/lOUDnEkr
9ATCu9m+CxRTVjMMX+qKJFEHDHM0eR4/dEz7JyqcEiN3Tamby4/bezUehQbjJJep4u0UW/Z+hWK3
gBeXvuIRIcCGSEdu7dlHPmxmUg19n1C2nGzFAJgoif5BAGFm14EfHPj3rcOgiolpg6ahFMgCFUre
JYaN7X5WVLV3K+s2eOfGZANeTBOsjR4gCZ7fhtrOavbn5KMjFmaySIl5JZWMpsePNFS1NZkSXA1/
O09wXpoyXaFIzM+xztlw90BwSID9xX+4exEYSO+5ieNf7jXwf6G4zGXgEenw+jl0A4h8gmOqSAL6
WkiJZtA17Vd3E4/OgkcByiMac/MFuQJRbxH70Q+gAwp3rbZS13ChXd8f7y7f7ySTFbDb3JsRkOEo
1jmaqV/CrLquJJ+F/8JZVCS+r6VfAJiLN2BjNYtQ3u1NEqbRp4VkGXquA9GxdsdP4vzzhc/wGBAC
CSh2eZfT7Fg6RgD6vxJm5PjazRKrcMb2nDTTV2iqn9Ke64kCi+AdqFF7Eie4WrgjivUSp0DuPcyt
bUlk/xTUaACCYMKvl1IHIlnorUlPucRuEQpO4ANhWYsFfdoowtc6sx2GnuUU83uWy5gHeB/CVwPp
IDeURONUFbc9vSChi8Zhu2U4Wvyh7fUsmImQQp6Wd58SyVU/e01vcvFuxZoVzA0Fs4CCIxg5/FiG
7BNQQx4RqGTj+Isjl4VBvH/iOTwfS73qOc2TgCtMzT0tiYXUvlUe6CfDxW+0rPFlHISJ7k/JlkHB
HUKZuvaXamTyuDZaEk6tE7/LjuI+y6d7NoLjj1F8/MnOm+FIbTXepfdGn4NQrVZ8WJ6p4s0qUeI5
ArSYUBDXED2jbonWNXBEbQaAgUV7iqKv/JlHROJC0uYU6DauaG3jagpGfmvhf1W51G+PIq+L/CqX
GLVw3UDRSlTWVQCUgQaZHys+uv0+NUSlATyuL7yNtUdD+EbRxL/EMWa+e8tLEliJf5yv726IdUoO
tWXSAQChNmp8DwYPDWCAgoafWrff/pTBr44saf1vem66vd1nZ6P2tVTm6IKKC6cS/KnQuQDNWx1i
c26W6AGjJMnutOIwIkCtiHlJI/UTWBEcRgidQAxkeaxE7al0tVZJeEb7oDMlLp84XgGV6FqDsKRK
Zegcygf2kcnc0PVx56UfrUT695L961chUJRYs6hYkH6RvrTqiKEyuDJcLe0XSvKTsuBDyXUEgQT5
k4FnixvghIxtleEmj6Z61Plk/jXFszr0i82D7Z0b2hWUjA1H4jFkyuF6MVXUkEj1OmnDKzEydY07
Mp/k+8aa6iQVIoKTEf2iB0lX6/zRn1b2G+UpZqQUctVMPPWMb15oSdT6ZBQ9Gym0fHT8KEYdRCTr
gjw0wdm5AJcedisqMu72zu6O4bec9lLp32llw1oKm5WknWrkWEC+ZhXdpJfX21GibwMS2qm4phtn
yUWqPJHrT7J8mEla/L8QaDt2KXMkNrYOF8aTfZJgphrN8yFnA5GP/XI2e2gGSBheZReG9ZwN0z+n
GFS/7TpIFNkrvgqmwqSC/pIL669B4H22t1LAcrdMcywkl4nogibBNKPZaXRIKFOfG58kFvDlVQRw
Lq05b1dNryoksg57gQ80BBrBZ2VY5NR0iQQeIW36seSnqlC9qg+ARam1ygiVsYFRJf8qblVXwHDx
eis9rR1+I5xt+JTQH/dHMh6DvXxdm91sNdauh4b+h98BLY/fwMjNUIpdVAm9bNrkbqVKMu83cYbQ
IEborHL3Y53WNHG0sayV+Bb7kMdjUixb5DG7z5w0iGbTKPToXD+NpR4x8UGmq76hdve1zRhqgdyB
Yd32icNM0cFBN6tfg/qPySUNvMrP3IlcDh+BcF8lumuUKb5GGCuggjeVt1iACSZA/uvBuOBrAxEE
TmBp8d3KgzAcdIpiWbuUyIX1GrjwKGE7U/5Un8/zQV9t4qvTrs63Eptn1/iMVZaKkykMKVssvWt0
JJsUlxRCt+ipf2lXrX4JaSJTkHC70xzzDI3q7JtOJ2/bpW0FZ78+QdWWKqM+7VosTNy+DTWNSdou
yP/LsMGdT7pDZB41XOyioxdj+P4av5rvj6TfPhLIkgVfClsJU5eNaDgHHps0v6Lv5NMyvIYKWsAu
zVsOpiDNiMxHh1xwNyaez945NdOhen4Her/48YBeJozspAhp3yFC4XH3XGPVxp6gHjzFZTPf+aOi
irtUNObGioyRDsnQqZnNojNTnNdBllm3+JE53rRJee2/YsntofVPca2mHkve7hZSRqX8jym+g/+2
1oAOpEi3uara8pKOa4amNJHvjokPhe44MA/tkdMcEygLogMY4UozUkHutOV1tUrltlMPv3+NU4rU
RzrnC3uyflGAi0fGJKHMNnvHXTjyx7cOQ3r3ZQmCoBCgTw6lJj53fKNRacSPc03+NHP37kTC4Xdo
u02zZF5mLYmxSvsSh4eB4Km7qpIl0upttb1RP1RUn/WueXrkpg8t89GYEIsNE78Gg2hpy8WwqW47
HU/vSoCsWRgi4wxPPpKvhUJmjb/mU4VSGERlR7HC0av7Ws0V41VsKNF7UTj2GqZhCQDimHj2lt2I
U35H25zP/NAnRKhlJU/c1pBaiFpemp04+QKDSV5bTiDsX4sIOoY1mywo5wEDlYyfGprHXyhN6Q2q
7vQAbQOFXHKfdrflKIvvPKJfH5DX2t91RkkuLRS4oQo8e4BK167g/PSHE1EchwHKAQj1WSTaZNa0
h7VXEDGKI309A4Rk3/TCIkoK1JCgN48PIUZP6Uh2AEqTn6NFaCzaI8OGjC3iGwxOdBXv4JkpzR2O
g5v3jaZog402d3MhDzDPbqLFEU/5DIi4E0H08L7W2rmdDyTXoaGOVvSyZO2UVsaxL6izPJnj9qE7
2m3+8LR9a1ifJHN5qqXMh5xnVzHMPfM9Tf6tYBAfmOqL9rdRCFQhRp+PJoQdwqqQi/DewpTnV7M8
OKpX24e/w+zV/qcQlojlgjmHmM/wgV3WuVfhUCfo0YUKUvGWTxYF669D7RxOsMZkmr5jjryWAMz4
uoYPBATTKMcmW8cKusieYW4eSv9a4rRlkFIy59OuHHKueJbPrtnzlP9paNoqmMier2vDInDCFrtY
ANw9H90YXTx6uNtOYpDTsqFLzh3345CUWvC2mKBYLZxpkY9Tqv4yRxFB7r+kGvn5AzOnMtUSpQpI
QmyygsPlNj6mNOoVA73qVLJ4kaWhdRvCUnt/htcwvSiPS1hxMX0cwNm1h21BtAcuc1mYBvdNaXBJ
HBjPvb9DjlQRQarlGUdXlonnj8Pa/OOEKlda3DT/zobAQwH15qUqgo1NAMqxnyS0U44nyo6PPow5
RzMwSo/8UZ9O7tEX41FJtvo9cFDidBEjJ6+G8mf1FS/8HwAXHJht4a6gEncJ637Zj+u9MfT8cv4Z
+hqVBoAZ23Zx2w4SLJVq1lbOQBmp8S7CnvTesYEguss53QLWgYdHCR2GGayzLBODfas5eeg5DZfG
0e7kgQ8clx/3YOcHnaw8Y+Z2md8MOml9ibtR/aWBTkB3fHN2gfSntX9vjP5ZMDmAH2uCOF9rvJe4
7dY7zkEm/9UOJdjY/6G6BehRIg8USI2wPr7jqjzw6yiqPvPatXH3Q1N+sR8L6s/fBTD9lvSHBnBB
za5/yyo7Zh6+Fw+JZpYZImG4YnaX40gVPQyeRQ5QIfoM90rqKnNO8+kB28v7txOJHYBfNvollIO4
tPPWvgAnkoSMOZ8Cztpri6ReEKh65Q3f/DQJwgEgBVliJH2WieD2mL1eH8sPH/tTf93pXaLf+Hw8
YBmCtbgXgWFqSaLKjM8v7JDcNECUTRyP7DVZjpFzpr4JtsKcBx9YULC58JlIE+bvRS02OWaZNLzU
zyKASg1r4MMMH0I/FJ+s2ehaYOSWkRt17H/j7hORn1Ipl4hq4imSYBgzSB7dVCyucJ1XeuE7tkZB
6ezE+PmbfkNlupRKcGtYWcsWRJx9UfiAz0NJjc1VTaYmNBEoqijEYnQHr7vRQ12a69NSf9BpZ1aJ
OH6+vi/rsRyOm5NevGoDZ9Amls+1Q75Tokg+Se4eZiJrvFKYe4UB6/6DjhSXqnw3SElodmESpu3F
aItIED8fkF2mHwv5WJ+wVkqGjCIJAodhvIxqCHOpmH4i4FBjJI+ZzucIcjJ8/4hpaSj6k0+B+1rb
VzOi9qQud8XIh9DVRBXxDWqI5RecmCBuheFhaCn+ZzcC/uwq5S/dfIZ6KfYxbOrZa8+3qQsCVEFG
45whhDS419ck3qvPXpCgJcB3skj4Y+gPgTBwtzIsk4RpyqfX15wSrDU27QmNUcyebcLAHG4ZClkN
BcDsDTMlgeVT0UBZuzwbIeDSYyFQQ5eJ+tSIGkZ3E1J5i0ywFYgBOHP1THrLp2iKzOs5VPbZNjyC
4/2K73PK3SGoF7TZcB7ebAhL8JyxZoj5qCTbztS9F7CcDMdLzxX+KvBl9TAWxntKyKlxxetIA4AX
iCb0TFY3v/CoepHRhTWUEWajpefe2CO4gZilOPg+OUpvEvRiouA7Yk5JPXDfUKSkOasoa/iCfdnl
Gs5YUKXTk0os5UqbLfpB+sEU8uYYX5tW2r77JzI17Gdb3w2D6slyINJiXpj+HH5N4rP3OrmUc9Ff
s9kArYIPVVcR+TaiJF11bgTTJ2MBAZeK8eAnRCNxlYCShB58eSmMoV0/RUdo4DlGRLTm6lk+5aKE
d7loHCAg5N9sWUDXaGPxCHL+nE0CdPcbYRaJMt41y9z6uJokrrkAv75nlpN5m/y5T0FqdiHf3kKg
BRj+Q8tRdeiaY9amZaxfVRHMj94kDy2EwRiuR+LJK7RuQ6vd9GG5sT9Kv92bggSzv031dk8hwBxB
6U78YtLd3dBO4vgb68C/roryrqgUur7A6X/Nt31V02RpawqsTvc8gS/84gAQGGu/5rLL51svAbB4
ASoWITfgoCSKy1CHxnpK8Rm+eqq3ulIIFR/wG/k55ZEw8qTythB1XzCcyVxFF7RILZrCpuejYSmM
GQV5jdcRd5M0YRKFiovakGODA+Ky6zsLvKbSbuxPHgyzPlJxUSCg35M67ne6+wpM+vkjK5JZZzBM
BUk7IHHPhHQIVnColqVfow3bsNpSkvniAH6jB9ULzgr52JwM0ycXKmFJKEn+WYpe318BPwvT4brl
eMoRgJ8do7paoV/HyfQ11aYOsDPlsD6CnORvDjxKbeHvHio55k1WK1CWMrnFxRh5rYHFXnZUClZ8
SsOGLn0kSg7TZP2hIn1h4LQcBhrjyDIChvTMmceKXs/kCXWiV5okB5YXgbv80wDg9YH5r8PokFMF
XRHQHO72Ai0jXy4Z1n0OSls3t9+kCo4inqUiP7P9j3nzHyFwuwHl/fytxo7ute0ZVyVE773voASR
EUbUBO8GDfe1qFye8kImhlErgI7L/IwyC7W9hAET3yPFUox/53ab5KQ8odmyw8M3t/nX1ED0zK9c
RA8jQ4m0tQ6wtmFdJJWatm1uG57ymjtKCFW6znZ3AoNzxf/nzJeaQpakhdff0FwnAJfzq8qx0e4c
L8iUppc3YuJVVKUFl05f6v8yAk08U/HJLnDThnbh+PNlwzrHVmauWE2GMRk3echhvD7LQK+W/yWo
bbfXxasbc5Nypntjq5jkBm6vZtKu/XPa+9mjlqdolXQj/FNluCKu2ObsfZZHJYiuyTH/6kPMBkyC
nyqDfRbaAa1iB1evh3ugTtwasMM6LzHkiiDsct7tDd1K5YjeRyclVlbOHted/bCcPVZ8hE0uZVB8
fnAL3wYxdGS9rTbHiOjSJDY3pJhHKr5OQ4dyxmd+kAdzzQDZRx3EWnc148uzPzRZorOuV+z4EqfK
58roJh5NQE3lpKnGYFb6JQj1rRPnICENr54DyPJqfJ63kNMfwLBUXZrFD4tL9hH9CZy/G5CNemHH
YPOfo9r20Bs3J945r/picNAL8hvUWX0r5oWqw4AE8fXv9vHWmWTqVCW2qGWaEyWIKThPol/rzvTg
s8h1aWrQsTmveNCKG+YFnE4YE0Ku7t/nvVlfjI2uu6Bon6AIhxweV/b7y9dpeSyhAZSXfdWgj2Ep
962mUCz/FwpXpj9tIhhFeRTwWSu4b+IaE5d41z/v1iRFak59L4prbpud3tx0BkJJgm2+MF/b/qZV
DzmiHwfza8EPuIrjB4BPNbHpJi+eCPEtvNBO1J1Qqim3qQq7WA0/dK130Vxh1w4F2injk1yUFDxE
2p7JFlavzXWtlsiaKumiPZKoWMpIm88OZGWokXCYQ6mVP70W85pbzGQeyqwwA9nWPWTkqhQQ4NZ5
K647zeejn5aLoaD9U3xp5L0RvnYj+CIR2TmMGYpASIDpQa8rzjOvmsxsWKR21/6Ws46yTbHNDgFr
OMh6GUWAowxJncHPW7VOos34hILk+maF/m9jglSsA3eNyI4N8X18fo9botBQ1fkh1D/PYUMRcr2c
KoJM1dM/Zuf1c+8ns/1VcVMpGTMQoVrj2CzwqlJ45UQdkrE4Of2dR4J4M0m8yW0cDJFlP37yOIoX
koHjGXfxIPjxqyuRrdNUN1UWW/CgehQXOeI3BjXofBureP7osZyUzyzEzZaKcuzt9NketuU6WKLd
9QJ0uWkbST373CFdcRk0X3+XeT6JQGKDGq9WqGY/+M9ygfwCuCNNiP3kIju+pT3c8N5uLUdZPpx3
yOuVMXIyrGHpZWyFklE+/BHsrF8u7HccaScNiDw5D/XEisFWFH8v+xYp72oh/emp5znGv5dRK3Lc
UeQqm8ustKXEg25a27wwJ3oZkdzIQyuTnCP57Vmb9Lg93o3a8D3Nwanh7D/kAdtI2Ij/oKXk875V
mWG7Nnluo127xY4Y/qlcFtpSSoaEcf+eTCc/JHztb5smP3zJnuq/yJBKllOth8aaeEuBt05fRlxc
LAYH0EfZzC9eiplmmCgAHOK2+DMJnQpp5qO2lFmT2JtrNBo2FvEsw+Sbun1ZRbgQTX8vnzy2CCW3
EZNV1R26E9TMipBpj6enYE9HgY0bTTWFQjzKjIzHfO8GhzMzEP9tQLnDWegYLtvSFPtZgq+xzztN
kRh/veZnDqtv8YT02eizNkSpDlzrWlddt8pzqZSkpfoN23SrWkOnA7z1/6hgem1erZgnkmQpAm0Q
Woc7cYFhJ3yuc/lfTnKhNGvXXqD/0AW2y//NjKN5bH9vqDnPKWjPWI8x/9rlWaXM5vEdpw6kOM2J
+2v4xCZ5l/XNm9FOQgbrvqX4eRE6C048anvKs+uMOr+fqynk290QwF5y/wNRukeVoT3s8rNK7qcH
ER3AuuIbll8MXBzdayb9X81QoO2MCaj5GNiXzpfernN56OTX9E860Y3FDbMrL/4SbWYyn184j4cw
Q7ehmu0HUPV4/dl81Wcvbtc6vO9LpjCd0XVZ5BM4J0Blc0oiJekeSEzZJPNISXj9NK8HS+xUy0Yk
lrPs3f08smtkfn13YPNStsq/o4PLusPdbajNocg49Ih4gZgbxju7FKkURJdjsW8qMjxZ2fv8Kp7t
GiZ5Qryxx0q8dduk8fFPrv4K7akV/tF6JND/77aC0GKY9MD8VHUVA1Sar7Oz6tBF30PSyHBC6/vo
E1BjJOsrtEeH7kD6hvT2SRcidDztDpsQ5cTOS74AZwpQZFl+yOLLgHRze7YkJq66lydwP2ytOwfA
Ge0o09HiaBpYkCiYk/rps+gFTZP7SxxBg+zAeQgNakOAmo3sbipi/YLlBW+rJa3vhOkEAatCaT2M
D3PulIMkAf+Du6b9qb5qcjLeoiYJdVaelaq3XIpa0sQfZ79G0AMfDjii+gXf622QjPpan10MvXJP
7aGg2CwqFRZ8yKn9+zkrGaUA9NiGc2bxYFNhEiFfipvuJo3S7o/eFZ0sDg0yh7xbwhrTANdOMnNs
5gtSiO0JqD6C2q3YbjjDyF6ON2MUyXfvFkXdmF8jyFNC9AbrevsKQtNvrjAL6uH5MFBBTEMmukdc
JDhsPOg05MGJob17exZbFrlxbRN/s0pW1bueRUXC6lZ31GZdss3HoyZT/Bbi5jwXgqChDqpR+pFa
1ZLU3HkIXJxAMt0Vlc8SgVaFuBh3o960H4ivHRj/4Ibdd7lWBmzYdcOpq3c0+sf9bqVEW3tRLVQ0
6zSWHhR0SP0IDFyhsvGjKVFfecpQcp0cEwEpW33Wgw2E4lWa2DXcdfGUkE1SBj0p2ounCYMeO4ZQ
HN9c1PRgeZaBUSV4S04AvGl4THxPGZjSgZRXgCpHHtLgDHbiNMZnHDNjtFKhr4wNMu6w4/WosSqJ
15NhFKgd55+NVPmGGWgTqj28OupN9LhKeOMjz+s881ZQuYe0L8pDx6blvYkH1B+w+/+xn36p1pa6
qXn1IPoJePddr77whs5452m4GmmseI9BWDExW2u25+luALnvXgWODbN3scQM3OCmbquZ39NUr9xd
rM56c4BAlam32UVgNz+XXn1t71cwD1h3p1gGxun3VuWnobxRW7SIh7BLCqQLlMjtog58Lw0VxGTP
NmQ4H4pDq9/Hv2hZDhhxTuKIMSR2/E4RJDSLQzmpBpmvuowoheC2+CYnslucoPT1KHOoVbXXRZQE
HqYtzS1ciWLRG9nhVbmRFzn04tGyk1rMwPvyy+XIgYuZ+qOhDphHZQCP+TITkEFYavNYGyGPvsJM
pZnrL7MtYuc/d1ALGmZaoSDmUgmumP9TGtv2bokQrCxEuUbNe10j6S27HDBdjPGMW/22TAVWwwTm
XTp6SLX09C0ps0GulZfgoqsumx/rhdVJpB5u+rHqZHaFYj+T7ea1m7Dpvq8DCAy+QPL+eKsY/TxA
jVgW/q/6DlKCEQ6LU6p5eSrhQtuL6xY55jpc+2VdDCk95K7xyzc8JqOiO0htyLHWV4BBYp/4OxTS
DCKdybMEmZUWJFZEINtSEDaBJVTNkXkM7mPSfVQ3jhDDz7BprBeRNtfnkkHaIvpQpBfMY7b9pcB8
K7sZtvSbXsNR0p2d+U44XCG6rYURb4Yi4c4GBazmfvjglp1acCpY5uNwk4Z2fLWgmoi0Cq1OSXGw
tOfXTJ+NZKzg1HiVZp9FzBHFTaOcaHEUOdbjnSyjv0gy7n7QtHcAGEIJEVzkMNDJrM2IyEuS+SP4
4lCyXQie0bDQ/baX7HzK09ajI+wQtZ5SaaZyGeJ7BhVqBchXpDaCo5IKbuEtkCvgOsf525N9vkvl
ZWuPUatqiTw8NjxjE4X5agvOvo10j1HYj63aVMiIrXhmrReQRuJ4pk838SXGBfBy4JJWqeIxYX1p
w+nkY1E6EIVn++0reijg9YvVQBR8nwxy0if/aemroNc9u++cIOn8y5oujb5ON/NFI/TV0hCFppEY
xFWIdAR2+zXiBc/RhyuLqSd306S99moj0LPHZSLTGEbAo3cESwLc+rTa5wfDZfLeeFtXuJp6Nz4s
e6Yh5/CcXIpgOS1Td1W0d3f/UGYMN/suskQn284UVNZ3fLykeCuEMG1zi/boTcc3qsTXAOFnxhZ/
aPMu+6Il3YmZXRjT34E3sAsFoEaGs54rjzfS8E5EJKYhSOqD1ZL5ZD241Hyhizi2XntGSs1+5LXf
s4eH777R8VxbauiZyj3R/rJ3EJ8WsUocP34BqbsUDoe0E8smLgHnmizfVTm70ikdJkj01gka6KIU
XwFoGGjbQHLbBE7Uvg7K7wxxyswUTeRdEqQLm6W50k+JFdTRzHgsXKi9p5XiDetM5icgXm0PhFb3
Cr7Kz+uEeXKHELvDY8gtE8qG3XW74v3IiRy56Hogb2zXXaLUIYZUfcrVsDXnAQoNBbSNVKMcUy36
jBzlTFgY1nR8qVo9e/5rvb6FFa+z6IXtJPluz43zPXFqfbNfCCpZ7ht7m14BrZnyEOBlORW4pnef
yjmC8G0is6Y20a2rqQo9yiJ/kA2j01RzV+sqhv1ATvckr6PCoe84eUaIZDkVEWGw035mkZU352YU
OxOHLIm1/5Lj9vQ6Ks4ExMqVsG++NQVqbTsZz5mrFVOe77BdN1qKK/KFRvtyaJYmXj8C9y27UUT/
Hwwtz4TK87nkyIm9agynHB5JOOCM2FMTwiAu1Xaq5Eq0r9x1jitTQusb6kkZcOfLCT6csNIk1iyu
5fiHBnmCvkFXo7o4TVPuUEDCXobp1ISS17eFEu3ZNvJZhq+DEBlkkqfJix+NOjERz74JrWa9oI37
3Lb0Vp5ugZZa1BG0e8e2QfaibROf+7VqIocmZngZeZEsXMcL/XhbzEBi3A9ezxVnffB6CV4vJFPi
NLuEwGdOWytQi5NuTbR0cRbnm0b2IBsOuTZqgAOjGTx7aCwXboolUBQJhnMHas1rnJtnNbM9lP7d
SO4xfI6LzDFoYBNfuGqEoyMZwiykqjIq8u9Ia6AgLTFwORruoji8l/H5Fog8lKpu42N3N0Nkr+7b
1B2kELWo3c9ST78PytlNdiBSKgbbbI9KT/6HNoiKVfUAYExYzyTvMLL2UduMzPoNKr0CXwKWou8K
jKDJs7ww+MGR6fFoKJFZGGFuiS0tM3g4vBBuFh7aszdKhX1ZA4ZrKdWrtxgXASyczigaLX0YqrFg
t77gPUaOhERwT0zJYf1/aqJLot9vOBhTQY+6AwFuU1E3XdukN1QGEKPHOxQx2cNROheRBHYse8pr
qvU20SmECzQKK1tGjglPzdiVQ69onxXz8GOAfZGLKqF41jOY6BeFyMbXG81QnBElzIrXex83R3fW
/cfhWeBITwpDWbF2AOpT3jaJt2DsUCnCaFyl5PJKn33KgU5yj67jXDOtfAD1BiElqt6qq2bFDQTo
fBOoPuN9NlW8UsVyChgEfKV0Bx4b0Td/8bJ4ZSRD6CV3kqNmQRLQGOJlgHnnSCX4Tvro7XkBW63c
dXwDfseq6lKGjBHroISpm5ADhkuCwxr1iCCHje+tNea5T95U+zCzzcumdmPNwmUVaZgb4IK74F6B
ZgXuppGkCpQEiawZleVNyDv+NNNhsGlb+r6z1FGVvqxKodXSb4o0ciIx28vdr0KQXNXA8pshXJ/e
ri1s9d0ebQkQNHJaYAqQ62hOk9LJ2HUFMb2DLh9U1Kd1mzdvMHWIXlXEiThMywmW1C21QdaDWhhh
kya/22KsBs1Q+XqhazJkENKWbZ6xkI4hG36BTa/Mqhu25yHwA0+wcz4+Xx8Mo4GNSIx3h3SZK59t
aDFA9uxBkwr8VWbb11OPKVAy0LfniYIeFI9DzsKNORD1COx/ydvf4XxHBnO76N13BryhcD4/edKi
/0XDotJDaLUtpWmuM1zZzlH+MP5oWSdd1/4s6ulemaK/NzSk12IC6Ye42LsWU/VW6SH4yAF3PSiV
fEn56IaqA33BvkjZ7BF9EuNhXA9xQsN4fcjL8jOmmCG3vmqaBrDi4rHj5PoSTKDmrbKPhIeUcwX7
8rrX4diZwU2Cuko+dm7HY9CjwoFTPH4depZcvvD5daIiZrv7O/C2GBJEDn/fj7pX5Vth5KrKcS9B
Zg/xP+uNqSIrGGJzN4w6z2bFnubnopBCqHdlKDZyfzZ5jcOG8NQ5CVZ/NluUPsyvC/9otRm8lVha
MJG02GE5E/sl9Kzu7TwKtlvoSRAbyTIHLmzKzyn+qFU21+/VSMyi64AHuHOT3cku21vKwAtHCNiP
Nk9VqrkEhsAggeu2DVf1j06ryu84RRnBvxnbJKgXAWtTtMNrDNeu1MoL97SvBeKDinf0dIBqGuKm
H/kYqn3qczheVZ7Qwbpa6Wja9g/Nn48hX+b/Xo5ocvFhEWlaT2jXAEncSO75dcD2MNGTS9wAvZdW
TbU6C5MjT3C8htOMNIHRok4WThTFBNNffvJOAk2Dk/qmZNxvcUzWK9McbRIuoqTrYedzOT7lHdY5
nAhsmsqzvKqgm6Qlu6mfmMhcVF1i7Ab8q2boH31BGHc7mKN/S0yJDlLUbqfl+lS51/My47l0eiHS
aNh47Zsx+SJgAsGJ8TGc4qU4oy82MVZKkGV0YxOz3B/bJdQWK7BUhdVYQAQo045dbrTF6p+t9Jrs
kCiXrdyd1oowPUHBIAQWi7DZ/T4XaKc2fMZun6yr2ZHDpXZWs53R15ebu1qh867sR0A6fboEJ2wB
h18c2El7Gnn2fGAELjuivRLs79K+jq0Y2juAt1W+14CMHTot1A38jXhbfhdPpgxrrU5TjD5Sy5dC
zVqhTnOKTmNFdBDOct98FNMOSkX631PpgWBwMoJuQDTsNIVbONGL6nvcY+4hpiVlX4vVBcGeXuK2
y2oQjsws+ETdCuXRTX8zo2OLM9eOwB8Z3bAAjPtcx3UIxLUeXqc5/2/28aVSP+eoD2nLmq+RgnjN
UHLUzXbrZoTBNarMtzTYt6T8nXxDQR/8sFj2uKJoNSFh3SKwuyyvbidpeesnS8VXhIGkq+PKm0mJ
8ozCIdDcVUFNnhK5MMbYjV3pCkETQbxwYt/6OmyiSNPy0aoW4PkL6MYP+U6Hxt3SdbxWaEPEtr+3
Nk6rcdWHEkwx0AYvHBZxDE3zDwIeN3JVH9hG6fY+JE273qpqLDJNPGZgcaVE/C95UlhF4g/Kw2dd
ydHqKpIqL9jc2s8aNybG/lqF6zlM5yTnYVc04F7g9bKZubf95pMvjMZLwmiOxc6wFo3Nlgg4Zt9e
Xg+Gf6rxuQTrPhxHQ+LWNungLalbpgasj9AyVV7Gh/OKxYE7GxoxkzlNhbIPf0s3XgCMGcAl1VjA
bF9q66t7ERbPIII3NIrxvHqvZ+UmHp+34y33825cFx7dWcyTI8H1NcqzU8ge+Vo9mSFNMNEv5I4G
nnLseLcLIfClMd8fPekobg/T/c6gr9vhHejkxT8ij1v8Z6ftpuqVRj5VtIaVx+hZLZeCwQoumU9X
L1jZW9hRoerF4msL4uufuoo7fkxyZAcV+5B7wq8MEmI/CjG/6uMUEMr35mpOD8arZWisL7a6i/SN
O4uSfzYv3zJnzlvk/qa0c+NO/ejDPZi0WyTuNJ+Qe3poELoCVJxyE7RlODRzlc/IXBeg8fXFSI09
6Y9iAVfegkCTp1Yx27mpvPpoAovrWinc8qD/qDH70YIZQQ/jyFRyAL9hbdK8nwwPUbMKbJwsoXfB
8UzHTYljEiLnmHLDmaZvT1Nm+a/Sv3nWAToWMd2eWendVib0QfPjupKEpxDVHYKNYlOU2IZlWNTl
PTlIUZynvhfGEcijuQAeiZPWfOpaI2zhBdqGalHVfQkFfBdh9a5HF0QsLrDL/8FOvum099zcewxM
xrKGMAJf9Ry8tDUyj6ugvu6D2RUuarR671j+temPcwIefmYT1Q6mYYsuw3H8rdwGNoxg9NfuD7rV
5cmYRAuRgQp9OIB9f1duE6gjof015eJFZ42Davy11ZbOvHR7IPvXGQMmn2oQkkQmgUhmh0FejlFc
idsOuVaVpBoWl4GlfhUXoTZnzqbdEs8g2Zyg5bn8nZ9qAq0V7KIcnelDAIDRBI0wpabFTwS1fUg2
IKjDanad2Ed7rij+MmyNqzAKzUO/651HVreCrbmQsoN4VK/i6PgXeabKEhgUKMwTlij+JnUECbbe
qUHqKGRtZnRQFYJJfRDLnE/fLG0oFkUkh8dY1dnapOk12bAKpJ1sS7rdT773T1mGH1h+TCYCIRMf
HU+U9HMuC7GOb2KBkZEWM+fj4lM8ftExaI5rKAUCn4ruXriA2bXYaXtzIdfd3Y4pC5FWo0rzkiwP
bZ7R1fi2RJCR3CglENws09OznHAx7gYyGerAL9rgtJDFEbKHi/lpVFZoW3iKpnkowh8ZV1i9/UM0
322TvA4BMm3Q/jxdW7LCHTB5aEq5cMSzGRASmYet+gtrGo1e20o0Jku2y2wdxucaynaNCVEFsuG9
odKjNjv00zMwPFAWTCwnpVFAjhN5mqqto5dEpmdIHAcGzw9SwoOuIavFE80rMr6LyA1kn3+iOyyP
I+fpgvMA0jxM6FYuhIPBW+UVPlY8aDtW3vMZGhMg/lTFDo+ogWT9KwId7tBozdBnX80r5JVV9lVA
zMoF6YCF6G2skaN9G/uqsTdWALcwffOKhfaaEUCl2loS33AsyLhOY0rAe+CzYcbBkL/Y/YFfXL9z
+qFA7MsumLUEDe+DxJKG7Dr/5T5RnlruhhAjy+zbeP3S8zP5YVDR4EXmST+PZXMFhDm/6jLUf7XZ
mGI0FBVv4sRFU0OJB/BvlRZJ9+1X/gZl0TNc+Fu2iE5r+FAQObajW32+R4IQKo4iHIXv2JvhfMIa
tTRxhVRuObch41Gek5EN/zuw/3UhvejiaKK2vmgXMeSyein7ajRfYUd1xLA8WW4f3gWiZOpQwyPG
JVfkre8/KHJs+aDFYQSnfNt/Y0DQiXI+DyKT7oqmwCxQ35f5iscplMcVQCSKJQ+KOs747Gv6F7SX
z3FOy+QMKQLtEzAynvIe0D9GblpoM+uZtTIQV185OA0tW3tjY9R6fclBSIkTfkz/ZtrvjqaPDpzc
CX+Yx5WFSUgZ6oRXXKtoXWNK7Et72/5hrn/47ETSedSwNsCfrlkQlW2q7H/qClLc11/9D+tXM4Hx
59M+uBTu7rI06vLcJTsn/oNUwvNNGUQHTUs7i2vklmXX7lsG1sPxrI7qgC85THwfVrEn9rah5DVT
/UUD0r8cPONsiNFkhueylGEqlnoF3wxbuQtvyYNO3I4YsEAA9c3ZUuercutxb4wuW1WxvwucFp/N
H5H2HDPzjbvhppbpDputjo8KyqKr8xOrZho2+x/WvXgjFoplnJAs5q/WXX1Jzu8LDkR1pPYiVm4e
defo2n2NEoJgt6SX3eRyHYAk5GecuL/fbhc58scj3QRoHqP20gSU6pwc/PMdI9aSekenysuy1f7B
C+XLy9sheemBlyFUDlkZMrr8Eh5KzQyBTNu4Qw/ZaHpi9506nFFtR9tYVG6xjg/MQMsllbPAUGnQ
qDYah28Wooo1IgaZf4G9QdAnzIvdJF9yFTLk2IWTtlydfsxG1es1W3kg+487Kp+uKFx/nXO/ps1z
rUdPzVsaWCaCec+Ef+CPPIqqG2eQJFiAwwJJrGXU/a6sadGlm4HijOYm8SuFMyfEshpdW7Lak7w2
4arRykSy90feLZfdLFALTpmqsazAtJYkJNk9GmgIuI20je41BTPCexJXaA0LG2gprxRSKw2ep4SF
+jH6VPLPmShbMzN4z2Z2kX1R8rSOryuM3HGJ/Y54eTH2xHITG4u0QanuPSpFX718yzt5WaOaWjEG
cvHzokjgPDvCmDsBR42z0Q8NuHyfIapCkR9/Fro43i2150TBRcdXg1hRr1qPkSg7SGCzHI3aQCnF
IETZTnzz89LgxoYVZ/tsrpkUXXGxo8W6+ZLaXtKurLPcKHnuryacVHilC9J967FzFuLmlc4oHEDO
emBjgmWivncKDDKbKgMq9QxTzP5cQVbn6gaauCprsc0M7ogJkEZT/9DSHNWfL8vlZCNGTx+g28KE
LSrN+pxEOeI5yzDFore4OKKWD1xHouwNh6qumN3GWXvBtvaaTabWEirlZpUh+oIDbbcBejCFV2u4
U4L1vn66ps349tywO8G4QQbKFnIV228itvxMzXtLenOtPzdkyog3DILFQxSTvyaaafoDURPvCgT1
xOvzi+ycJUVfAkE5r9i+TgKyk/a9P2kuxJrhn94yj2Ms7QUoIQ8g8RbPEUYmhi4bp2ib9rHCBRjj
wzDaycQEtUXJ6GwOolJ71+nQ7cjyTv9xw+DUf+8RA1dG1+T/NNgWYotEFZbGIyU1LNe4tWd57Bvt
V2hF4cVKTAfTLwPTMG5djN+vHSCazJL8hO/8v1ZZDj7yvGn1o3AtCRCjHLFOHUmkL2xO4EllB13q
QYw9w0jtrrITD3P8o+n704IRrNtLZQHKhmX3CUdg5RbzN8ofnf9gjAd3Og7shVxkHtRMT0eDfa4e
LrhT1IMcUBrAXEyZyyrEdGMdlapJtio807nmfkKgfTIT2iw89RaZAZtFRgsmOF4JWAggAk+BhjPI
ra0DjBYD5K2dQYLsWcvTuvfc6zNu8pk7AFu/NI8dQCLhkDX9MbWh98q/ukoo8HFTXpjUAhD89/j5
/bWoqEa/1le1y8eFRWuxjnTw1yW7FLU3yoCaavO3InQlK6V4y5ul7DjcvHrlKQlX5EfEfhlA+z2s
1lt5wT3hAuozLDd4np6pY+2Cv5/bPAKgg0xvpBV4FgNDZJ9K70P8uRDTBj+m4pq03Id1WAB7c3NX
kDgfRqeD6iWWjxHr0LLNxhHwrhxd6egSBN44f91pDl+F2p9/gzS3YNkTRpK36b5NexFEOh0fApuR
ZGoHZlGUSRXuX+38CmNMhmHd3gXfl//nce+fhzzShqEPLBR29szri6JZDCTq+l9EvX22GYC7/xYu
iSgRI7bOrgT6G6JhDg1QluAjCsWQyRsr76UESbwtznQe5ytJ5MZxqFVDWRjIYbzD9oJ7EZZNl5wK
eJVHXNj2uphD+mSVrE1Y8vSn5TPpG7fVwLBjYqL0DQ42d2uVx+0h+1zadfzQ4BVRYOxuoAFjLJeH
/W96in3g/b5IEEnzX/DStPkRBc5DzYpFyR6AvPlSXoLqmGXL5NiMyNErsuv2cH3eokelbUkpodL/
ehsEs1144+vfksMqtifFpxOgC9gitvM1HoMYPRXf/QiEe06d5c8s1XNKlSQ9Eu/M/ctgJ5uYCHh7
aBsV1Lzvyd2KbT3aoKdQxoRt3HBamOOBy0EUpZOoIS7CUQvfG3tVrsyFF+TscO86S8t+rHPrhqfb
yiDwVF2tLVF39tJ5hb0XTQmV+gJN/BQEws76Ud1HH1Y4IudngwHF0a0WZJte8/H77UtaaLT227Me
hzL1+7zfouDgJVJCi83Ug+PYbuMPMUz9G5QNmWfkWNnS3Ii5sJOuHVUQs8aCWzMTg5UlW3wcDlk/
Jf2ruLYcvVX5S9h8USdlNqdu1R6UCrB7iIcye1887VXPJ40hyMLNzcomkzRsBhjoRD23QTGrz7zX
3Gw1s8Cb7aFgUPI3uw4K4QgVM+zohyg3YBBo+nJnGKMJZOFUOhsXEWSUuHabJs2qTp+Uh8JFaCX/
0YkRWApapqjl137l9QYd2gHdoPEOReOrJu8G/Uab5cK6H2nfgAuPxcpkeJqaHyBiSFh4etJOHD9n
QFO1l0MCdboetaubA4tyFYo0tGftvMYyVAvMxnwN/F6DnFtTEz3e0OF7jMoST+VdsNAumwThRG9g
Rwpc285YUXW4r6PpwB4ybhuwJDln7lEnkOroPkoNkLejCk2hnjOjG/YK/gdMkaKo35MNUfdTpP7h
S1MQm4eyDqG/LWHkppwVeJ07J9VqlmyRnAJLoBkep4DMvwhOy2SVpUTTF2njXCF6/ao8dnOxnJgp
F7Lw/AhofVZBRK0ryn8rOtqpWgaWoGPML4XEJNyyUW0AJ0f367hxNkhKoxFD8h81/nRSZAFgeADf
xKGQ4Ks0sVLkIdjWCOEJIImPVn2eNX71pUrUckwQRrGovh0KToGs39dR6vaVXOkThjrHNWj6tLdy
epw39golu23voTFiZg6Cf9iy6QVvbvAy6dJ2FHtNBC1zEwRHBbCBpyaQhiuLAaKhVjAWNGvzvRAb
V+SqbjhcodPjGpkzEISLshEQsfqxBhgS8ny5pLLUmD4i17WWnq9ZhUao9EJswc6uARqTs8JHs2y4
X3LkgX53aWGT13t4MDyhNoEmQWjx5Gprn1oQhI+Yx8MbD6r9gTQ1+ZHlRQMHcLRDEh40Un2dJ5Wd
W/fabr/4OEWstcBjm8JOpEHpcRzmjZbsBpSEsf1dZ9aequ9J68iRZy1rZu6YfO4l9Buo/EYwLLhp
978JhPdJ4Do/FM0V1URasXnVs4hptlQtPI+uig6o7WK/KD642CKseVu5IaJdHcaT5/VNf+YqzIq9
dDxOTpnaJQ9FLQAEPlw15+3EUK8mrCymAuJ2kvIxzype6G9O3uQ9UwU4UR5xgR9ZQYir8O5CCZdw
q8yAyQYvF5C3Fb/pINeQSvRvI3Ab5qEp40HHvmysT7lOaPnUPZ6YCpiGQ8KY81SBFFgAHRSznZCA
iRGlz2JteCc7aOAxV3iNsR44iRu60PtQ9u+nbHwnMuPqx2QZvYC9R1nCYy/iZ9i8f2Uva8QVRg+O
99LevDP2rik9j+dWWdtdI4+cySpQ0hqyZ7FyrHVQKHRrOE+J6m3NY/IAs9HtvvvC3XXbB8bzvaxj
UPEbe7P8siZdneW53s9ok9+iF3gZXB5PqN05k/2N6+uLxWhKGYyXM6sE184+kDYZ5BXRBM/kaY65
pT8CPeS/4Wo6uA8IYouT9TIqlAVL7j5QHDegEctUrin8ZwpZzsC+rHznFtCq6MXwZQv4g1xuJwtw
q8J/vUqmJ/3mesEi5CrexDi+begr/J2t/XJZHnVA18cvVgjKWQem+/1Ykr5tRDjNULFkabN0R7/B
sjeI4GSGOmczbMv4/bu89MrRfoY2Jel6NDLl+CTbHgBblhLJ+A7481AhqsTctPm+bs9wvypG3yrO
TxFaiPT+Zqkykdv7jx6LRVY3RP+519acp2V4/GdXxOberVzHqOoj5ERU+/TbbEKoOgB06KN/Ts6l
AW7xDqE/HPSWI8KS81V9vQGTdJgXMx/QsaPnNfQfkQ39oVa37y+0S9agh04Qr0kVXeAByb0kauMN
DvqRLbWaEIxd7KCx5yV2UachzC89VQKkcQJ+RZbDnVvpoWZu0cX6qFm1h6TT/V9UTkzJ2NU+TwIi
xTGNTHZb7BxV6ykS8ST5kL87y0Bh623O4a3RYhNR22h08iqBss1jybZM/KwbA1N5BB7LfKoHpFfd
3h3+u3PIkniA+o0xa0H13Lx0IdjcWJfNBeEDnIVdt4+3c/nZLQ+AlJeVitV9lzyvB2qgtg2CDDIn
IokUJPED7I+XObOHYdowl0lAoJQ2Yt7PIKH9ofsC4MU+GbDPEN4rvUA6JYKz+2H7lqzh01Cn5h/d
KBGDpzUsEWrM9yZNgi4Z324Dh6scd1Gxy+3jnUHTS4fd95Ro3ScnU14amG5He8J7U/L61dsE5As7
wfosjpQ/pwCWBqcCs9cf2WfQbnxTf3BqvqjJPPIKMlCUldOi1fy2oU1rXYORXMGElfe/CBiWMbZP
NUu8eR8/WYk0x8HwdJajMSGqrkAB6EvdLt+401FMskqpL4VWVt8fsBBGeQxIY+ATtQHdXCp4+Lbj
mEQYkhFDtOvDgqcdirAE8ETl8Z1rvzYaJulgtOxduyt+miF8D9jP549BlcTVagDH9kxzrzjfcrb5
qSk1IVvZyGij3LQuk3AblgbauaXPdX1cmBBdxv/Zx8zBDg35R0p6F7wm8Drns6eFj5T69VRraDzm
1Iim3YeupTizzu6sH8XndnnH4kBTZTetxZq5EymLEgKFh2/K7hyB5RcXYqj3KC8h0T0vBzzthhkM
25qAkXvBbqc6vVHxM/5+UQmgyTgZx0X2ZgrVpBlO2mDm4EjkMLU50rohA7rj667Nl6BdwjgmBFHP
FppaKT+mCO3lxY5mbgGyXJmq8EFEOlna2DdlUUdc1pNQpfAIrSXjMEpif9NqiOlv8froVMkHNuqh
4dZbB4P1ZuqlLT8WkLppEqw77+pqPsxAyvW4leValqfhDhmjQF+3Z0X52JOW2VFo6+pdLZsM0QJO
UdJP/praY98VAEZbJcCQXzIgez/N7MBFLxQd5ReH2v5lI7/TZud9DZ5z0CRd0KfYtSQI4Cs/Bm4/
7IzsxIKivdKfoRGZ6PIkZhYf4eeX8qXtRFAM6UTCRz2Zqxm9o7obJw96Yfbo+HaND2o7T6vwhkNy
uaEAWCooC2kDMmC3ghgPmO15H3jwrgdoE/86eIQCbiP+bqWNTJnXM6lsrCkx9fhPn9BgVjQbnVAe
TiKhR5MewnXkcjms1PdYs0cLFOqODVqlADHJOUcN7E4OCMsLj//jq7OK7VUzrFJcpL0vT5HUvOFX
LwbWRHQVP4BzPMi9EMX6FwYMRBgPoZd4UJ1xx8n0pUzmAuxc4L+1d+fz4WQLtogLFxECQlqC1lXS
9kZ4B0uoLSOQPxTQt53uKLJrwPAZG6QRj0iqpQ7O2xT0fIDpib6DUq7T1oaLDvU4ID4YT9q54oBW
zUyhA63Y0u12wL419HZcQ87Q5dDzHOviqPVDN4ljLwS9nGp3waCSsvuu3FJFY+XQSia2qLcYu9kt
NvA0qw6JvWOP9Z/tCUzGRigUuOq/sNSpfSA4Y7v/PHrGE1Kh+Knk8caByPNClZqyeujnOYv+6jrk
H2QQuC1qfUc/LzCDVJGonh8KcMrgl7TsWMAgctMRGN5GNDmLX+Vslo4Sc3bXPgsT0a9DtYXYAINZ
oIo/k9t2iixVLvXklfIXec1OaQ5nfLZ0GLkwhetBkg5alWABQgddYjptxaFUSOgPtlLIt0p5hgcr
mV2ObuwT9QiQ+N/VvVqjOgRhnvdi+l+lu9OYUlk7ZCRkKyYcCjpOaUVfoHHcCYl/bvxtSnXc4PYo
TOz+JCzuByU3OSiZGXKjSGLh0EqVMXq810unJprWwZ0OcGnJp6j5xJSmgbzfkYpT44D5dYYS6on5
mGdFkumsG7LR+G/t86yYHulkRlh2TLcX0D8iew7k9EDJaqoqstpYZgjDEBt0VT24flubOr56sB+J
m9FP7v5f+eD4oI4zjcPVleSb1AG50vWcb/zGyVTxJs5g8h9YPJHP6lzA6ZDgr4C0p8T4EwB9NSvj
nWvzll9/WbcerMjrhVNqmFZWB6JTisqLFaUCFjOZqQjdLsDexU/wR5l0n83vcOh6KpEJXQXwAWl5
QY1FwK+F9cBqkQ/2XGLO4eGjifguw7tcMkeTlHulnOnd9oo/QgLPyg8awatgpUHfj84becN7Kdk+
vm8dm0ipHr4bd5OifMa7Qw4WCVv/hqsJ6+MVzI74iIYPvBKU9t7hakQxQH8+Hdt16eSJ93nt2eDO
KSy0T4qxNtjA8XWMJ7snFB7Yio2iGJZKxAka4XYmHzMP5vrBRupf0OSxIEYyDRE74pR2ZYL5zUtb
D34KRU8VsJLip3CTwTLhlHWM5vceq/tAU/vhm6y8zCqeqkn2+ovDupPyq0fobETpypTS3DSf1R88
Bg08EekraQqcOpQ50gVe/nOz6W6focMdZ6lRSedz49YTRsft4gV7pDhBxDFLfOL4TwOeSNhlgtE9
Re/LGPQ5to0TIWIdwDz9RfigPYK9IfWraqUDaSuCNO1YRULgsqVsnLLx0zD82M1xMpfjA1w1EjXa
++Cu23pwUZ9Tdy0uwGkelRzXoi4neHFRSoD+tqJQA9YC30sM8KrhFqP5dcVZzpY9heEeVpEtKt5K
1KQGYOZk2VcWM9kwEyWZEmPACCieahTabAbGc4cSK827cWifDMQfSqPUKcQJnk/eiWZoJ7T8O20P
k6d1HOR6Z7x3oPn550g7XZSXcsscR65M4f5+TpHmlvQdpPC3aiKwijqLTEee2P0HfrI659CFc15j
HUEVp4ApUQQyHBG1j+i2zK/xGx2KKV5oJsXCvF4lcYKY36VnoueVMrwp8OPpo8XMTsijriRPHMP3
dHspfXCV75XeN5qU5zvdMIXK9xKnpjyh3Gy7XS/LBq25jVNw2ZdaCZMbS0MCektHQ5813hssP9Mn
SZc1IMcLNx6AyNfzYNNYXrwO8fO9ErYdoQAKOcGe9OF24tFdEJlOfSMtgP5pY9sA/EhtEXUeZik7
frG83bu0OHB+ajL3pt26eLe7FWxG2m9Z765xlyl3d3Gw5hQYBSk/YMne94K9JAukjnGvNRK3cDKC
9RqGUQ3g6p7Tzx8KDmGdYyktk71G+nU1tQyIOLbT4F72Jsv9q2NCMnXwZfKc4EuIfJ6UWNN0VNis
yZ2UaTEredJi+dam6Ma/tvF5pmNu67+hJSee0/jdu9rAF5x7/JKXYl1EYbKCejNzEZ2Ug1zAAQ9e
NPRh9Zhtm9PMkMv4Q5S/kc6xI1mlkIJvFbw9WY35SdYLkPOLH4/xbcpQfCgKktM5PXUH8KHmbb5p
cUZ6VbEhNgTpSFUvTWwU1k+34uX5KN9g737Y262HYVcJOIT66luzDVRe5gyNhsro3ek+0yNIzrHx
idli/Z3Y3oV0F3oWtery5l3NFwB6LpACIJgqkpA4eSQS21hazPWA68/MmB2+nQJYsXHSMigrORCM
6wMNN4B22APnUOgzrLEtwmYFMbE72wM5kuOcVxRl6NvwbHZ7Di4gAfNurgjOMgaBx3RkJRbHMl8r
8Jxeoz2Cay8xYgu/HFDGyHdHR2VMzyY+gerr99x1vYiwyhDm/WatZIxK1hGCo1+gBSSLBxtEJ+xA
eOS7UCQ2+652XhXImrvrWG0AuwcwkuLEGVQ+E8IhRnlMpJpSjD49yuKI5QPc9z0nN25dLaPICrIe
2Qb9ZGK6B9Nmw3vq73Bc0CCI+a90+Oy/N2gkXw9DI0zRZLfNfnyXYtg81bRRjvpklkCQnwqc9UUm
tqFiV/Wutn7s2fmZ4i/ahaZJeD1d1DThdmauKwn09HUijSCWQT5HplYDcN1Ug7ySJUG6EPoR+M58
tdTyFr5Sbt3lCCECJGj5e7GDayll4WVgotEC07Ulv29bDp//wTmWREmSXlltRjfpcL9aTTtAqz4R
mI7z5LDDca2hY0gHe1U5WTnO9oq+euwBvDOqxVeghGUiEa9xbkCiayJOMsEg4cvOSWnE4brTEq7u
c+yEFdRbCJJ63mWMvQ14dbilD9lJTnujEOfNcFWb7Klp489AJB6o6AqEuDZIhWXCTUs+yJv21vtN
YjXFbA/U6cjw2MOvGK4mOgguki2VqW9P6RaR88l+XPiS3KCdMogGjqN+RXuGlbl389uqfUGiZCtw
iaNcfnAsOnltApq3wvRXjQ9K9kAI3AHZ/wsPiJalhMzeecGrSLI2uGGd3R+NxRnwl4cYVwkm2BUe
DTGMa48dphJT/qr6ElleXmeSK8JwBqWew0cpTm9o/HkedvsuK8/vdF2PeFKA1eAWLQHAGE0WMl60
TwBLPH5jz+u9N9L0u4r4+eNazo0YMxIDgmhWj9AtmMbsKjF15RW4cMma47TXE+pJs6wsfWFlTVXP
1NCyHIlOBdUs2FE58YDzn+kROWUHqEXuDKwlkNkg9A2bJ6DetVxjnfn2GzDps8ZGoU8uWcFAR6Jq
b+aNI26w03xzQ5VTR2Qjm5d1J7xFUg9826QSWKZEQ4BPs7qYA3vlTMrzhnGF72kWaCTMmTSk8fZP
ABFFAxXEYPDzV5jF8QP7AEutC6kaOHcPgrpG7RMufNiXdjMv6z4nTeZ/YVozKS8W97FM5xdmG6QE
OO4pbHTVL7g9/woWf3oByS/Kot8ks+GBTeYMDeX6Qd+KPHnOKby+ShAlSVspNhU0LfO5RF4jxqT2
JWOqXbA+zHVG2yl1BI9dNN+Vllq/m2qtczCs6/Xp1+H1XuefLcz8eIrs3ECgeW1pEdR+ppHUf78J
idPxds5XxyZJS10GOP/IBDL72QUmBrSmZLhNtMoasXAU8Ab6I44KP6JM6KSfgwL2NmESZ15p5mB0
N1wu7xlH40/TWXLbpRYTKX4X1UoR07T/PUhRdnSiwI+pN56iIPyLFkoA8LatBG4UU6t2lBetKUqc
OLzwpDbM074xVmlx3NilmSMv97ygTzjjX+IgU3JgQhyTuZbwV5jaKbXgD5nrX7DqjUe6K1NkZDWn
pjJIDnqkj2qCX/8NjCvpnScE6TTDTIkf5L50xPkVXGRYnSPejeu4Wprc3a5wqq89EVDrHku7+C6z
9UPOWLebZcrGGu38o0CV08dEsjWCDQ+C1JN1vVAs4DZYHE/h5Rh18ppU2yXxHqIKRM0ylZUhs1tH
QYya7g5cbWwQdoiW/9VOZrE6HS5a1WZ2zzXmdsVwAvyspXW1F2SsDTEjLYfCuSqQWGYpLWgxKecV
3vPvpzoVhACT5kqUZ8qP7eUzmhB4jqExGhrb64+/P096w8GSpM3c981322+M/HJv9qxpplx5tkul
oVIzP5yt5iyJ+k2lMOntlv8varune8esUVzCS52y/bAjrjcgwJh5/CfnUJfMvcSSn1mik13DRld6
T/T3EwNCBvgdtAmrK+x1W76FTl/LpddGkjE4+0LBJ7ea9isLD6UFUX2K5SpwvFcIkB8yhtPA3wme
TvwfOvC8T4SeXlYJZbEeM6NJvfma+7a++Kie46ju+BVN8vPvg/pEWL/QUZ4WjWKuz5MJcYPwMv81
jURMincXlkqZY/c6t8xfeDraioYYjJSgpgFE5uDoSDVHYipCpCZU93CYFfX0A0zdIzJeOk+DsVNO
DZVhlAf8Cy3qYw2uQUKoCMDF/nMazm42YjDeFShr6WQLyoF6gPGRwdThjyHOlfJVRjCbYmN8zGnb
mJ1UmS+h8RakOQhNpqftr0Kv/0ATD/7qPwhmUm/PQdMk2uHQaEHWL5yI8vi3djB0elhvF7UQ37VL
/Xg/q3rOG47R59FIvWtEcJpxxzkguN6WuSkuewxcf3IY+4aW1TBiAMY5s5gLZfLDGqI2escuLiJo
O/FhpijYjdM18uDngkojLyb5veQSNGj1xBToL34GnB1CXt8MQFZDF4dWvXNztIyRpDusyAk5cVRe
1hVbfRfUcH5CpHnnqMZ84sB8dtabT/iNZUxN7XVnSfwwsAZMlIYHNU+zKmo+pMfNt1NNPBy5pmqH
PY15wzA+uPqoEcAIjdaTnNuWfKgcvyKddwqLPy6Ss+OreAlTbwsAAM2K3tZDoiEyKZDX3mIW9ZUL
mtjib5O0Et7LrefpqVLFyPpgpQg6ynoFQA6c+O1rmiXCfuCcIHNhE+knE8Ls0GqW2Pl7Uj79KIey
/swIoWnlsmYgsUJe70HiPaFtKQlGkDjy7qXK2RVGHz/zcWuxmy+nboLirH/XpEREFXMuViCu9n8C
QC5gOaeHIiCjex35HqvR2cX17F3i75LKKm8rVHkSXw3KBLOKf6Oe6l2XYTEHcA0KVVV1oadsW8+4
jRxuFal5HizWMvIskBp7nCWXsGwf2qSbSIUjBRuEzOcSD7PbfVZTPQJx6G1DfsADOGhJihfSodz9
NC4hOOevxzwIk2fQwgM2ho+p3ojGKc6/66RVG5eAkKzTHCx5qI50Ji+zkKV74RX4dFza2c0d+7kp
lw3DQYHQ9v0BDsJUKwR2IsVu+zLyBQ7lH0b6CQe9F8P72f5X2l828ueqk5A3agj4Bbn1VA2jO6cU
u/kXV/e4ZJztdQF2CHHJDRh3E24Gw2oVjxk6knA7pNQF2g6PXlmnnKqBMW3WTfffpUJ95tmYuNZ/
v4jNbq6w1ALQcNENP7JGP8Fa0j8O95PHXe0+08mRzs0wYv2C1q6DFMftvLbLjSKQKwxsTpt3YbXy
U14tMA6cSbaWGj7dn9VsnJPmTFSNTZ3c7Lk/uXNQHC1JPV26/rKye2CYSw7lVxGVbl1PBvdgzdfP
06h9uQ5sZU7Fiibf71gh2SOUFeSjGs5fnPoJV447E6tJkY8LsnQQ0BvWLH10FMGGLvbbyyTFYBbG
mRd5CmlBeH3WiQQdRUtRQwZlTsOclx43Flymrj0QU3WmGTXIWtGWSwHnRzJbdypRdjQ2tLhjYBZ0
6+D2K7fHt4hUrMOVbLD/Dzbzmm5DAKRpWDc0BfZOylt6cDcaxEBnK+V3ZHfit6upwB8Lvd+2QJVG
/rRbXQuBkmxZao5Dn7mSEC/obFX4xEm6B1MDwAhIJJNJJBXCb+gJkaONprlnNsiDsH5VTk2Kk1rP
vLMXK4qAyd7arlhpH5ZNpVCWYF6AN7R1jWKdh2z4u1qiSL7UxbRK782n4AgpRwx36N+RcNW9C/1L
9wXUvhW/RjYNtoouOABzEzTJ7lBLODY4qH8N/SqpTBFbilxct1Bx8tAVWuy0fzkzFle9JVvafTrN
BMuTRLY4sABcfcXDMcLt2IEspz5J3Vt/Y8r3war3OfQmBoHtRXKVq9HeAwRSe1Cmum+Frxk96WSZ
hbi8JTjlDBQVVkCECxEEUipCUTwf9bVj76u6Zlwd1Gg4si9R4r8YuVu8FTjTDI1pn2WODVyZ3+m3
3kRz9zYGOwei04WQRatJBvW7OMMZJrL2AYqDWzhiy7mvpGXkKMLotF5pkEfVrivDsAiFJYsmqezU
DsoRBwWHBuILwveXway+DefrCKFvaRgmqMAPVJNW0roFJKPGms4aZOZ5jz4ZEMC6/6NzvXoqV+8M
Hc8cP2qZWUpBsEym3gC2tnSpCtJkwvO0jm/EmmfFB8KzDEiudlYXEyn/15PwheT/BEuV14MeVczd
D++nFxCittdXhHCELgYseGumQdkPd7w4QBDNo9BpV/44wjjxEgMzkVrB2gXpYh6Sp7v1uGGyY9X9
TdzWMGnYrs2rXUHAuxyW6z1GDRvtRhGjwROV+PyD1W/sFhSfCAkTRRnyqIA6yHLKcROOOmrjSZgs
OKyqeaxL7HGqtXEF0oZbiXztSYlF5VZoih1COcmaO0zAqbSZdWmdb2Hnp49ksrXvkr21ojzeHaF1
96Rd34qR6sp9X8ghedkAQyfKGSDvkWgMBxe9maPdaHp2WpiV3LpYlS858gj6vUGuB1xXEJcaODfQ
bHojfh+AFsqaFUdkWS1JRfge5Psf1knW/RCENFuHbK65j928L+ctGbaURi6k6e23fztAop9oV27+
BiVbgqRMjXThfdLDleICJSfzehv7WdVlQz5+FCtqmp1XizhdMY8S3zSs5FvEQe6r8tICsUu0rqSP
fuGnpmYL4dzlveowCum2m2mgFBtDfDGM6iDCpdQCrAWwdUv2vHQxK4wTJFQa7fmfTstlhHGLk4JH
VXV5r5TIcCejP3sjkp8Szp5Dbxj2sK0VJSmE+uA+HP+r/vFR6KjILJntZeo6/N/jPG5Nfn4QRHtu
f3Cm/wWQXggT9oO4EVn7X1nJvz/TXQu9+1aaW3uWNvppc162FvciCBUX1lTTKgXQVbyzwGgOXoVN
bx/U2aYlCZ/EtREReVGoYF4beZfmEpQchSReHVJ9/KJxz2Ydp11OAPBd4T/ooR+Tsp6o6wxASp4E
u8ccoId7ekJ2fIIHOSZvp8sTveWkEjxFNyIm8Ea2JN0FDRYd86B37Ki2yl/u5/+5uPRv6MeM8XmV
xJzW2wUBetUgDPXCuKEEUGx4/W+BuVeBd3v4tmE7lzQOaRy1Jsn/O9vEvPdD3HGh83Vnrgs3AD6+
UDpWl/XU22DwFbyk1CAwhjKeQ3Ft+z7T5cnuTlQMvTlXkuiXTnhd7fRW4d70+xMuuyfew39p6eu2
Rw7IVZ+yz8Fv/LG2hgfaWdjTWfRxdhXhs61QPZpQYE9B+02CdPN/a+lhSAZiE95AV97i1Z3oI/Hz
PVJ6B4txnpPw4zuxiRYOwvFdbUL8lfDd0RRs14uU0oV9jTZv5qNbLU63kWe++vsw0dX0dfddVfOm
K+f05bYTC8SxUxkXtBxD0woSy+0ximb09iQ9QuFwzjKLEC6P+G9YuMW/hAWHTbRwnvftM0bkD2Eq
dhtlFi34Gf/T6jqS22+kPG2l9gMmZHxhXSLbpCM4XOlXwibS454pDRv/4HovhYhVPsYiGQd4EEeP
MoJcWyB2u3y2MRwTuUoqK4KgcWyRcGotm6Ne5dXvvXPNmIMDHMU9DtCmaTmEvo2YVCxRE7myo0zQ
lPVIdYoQkiU/Q2dO8kQonFX6yX/ium6zF2vPgnuMt+B6yxuGhiEFf4H/n7WzEPjqAF6NGzh6NBNp
i8+YdRuEF9s+KguFIHvv1ZEFR8dO5U1iGwT1tO3UNHQ3x4f5CUNcMHhbV++ojux7mhtOsqS//gzl
RBHnQTnBv3dJ3Lmeet/6wKQY8IBih/0c7yT9DV76N3+wpQ/+m1C2I8y8CLBTBMmzupfWPkq1s9fE
5XnoWTnKrkwLi6cQyQ6tosy96bH4/lgHcdOAgGGrszEzbyZs5AswAR/YWnpo4FI9/jJ+7mZZ7qr8
98c7agX6iUZqu9h9/wvVDTw7xGMNNILee03Y+OeGBCtFoqh5mx7tius3BTi9K0WZyqIKK6SGY02r
H8kl/Gbm3v5dn4oO3PIAAh8A8cEICp8aM/+bJ7DNoMcYZM4d1/+4aGfPi7N1CYExLwNdvPZ74oMz
XDVHpjbBkwsvyYMPsPhPmxPP1tRPm+ijxj0NEWdt6ZCWMzIj2SXrdqxeKRNpZVJEHge+6Fy4zsAR
+AKCJuIxK9Xud+ajwSkaE2xt2mYqR7TwJ+OjhUiuAEzvuOnH5O7OVZC3b3qEZKw1QAltazMUVHYu
spsragTpA83qliBd1l9npo+Z78pJDy6jin2t0r2EkRx9amFbTLp+5QIg3J7PmpIJyAdmBs8fJnPH
IWfaUmurmCONgYLeZbmHUHUVXW8pLOhqz7bI/thj3r0sI3ukeDFvdnWNdV7T4d2y8VqbO97WUW+U
jSTI9lWzE+KiPyl+G2rG53J38tlCpMMC7wa3lFI+yD9/ZMGSpNssEnVlN4fUXQT7bjvJUz4Bydpp
84G+oEvwtWiLMgIDDFUfu8UqgHC0Hz1aattZnWPCKW0IiiojyXrLVoqXaOMgUwES47SOoLJZfi55
wOF8mRxRdpXqYI6dm9lXZZ2nrCyuzm97XhXb3AeIC8TUQsUtkmELJAzMg5ayad50GO7XCgNZFYvl
euKHaaYLORnVAZvCIV1e0XBgh/v2gWnNDd39N/UTgrMYh2yX3KPwNBwrhSzT7yQT2QMcwcuGJTjF
Do7ndXQzq0lOJSrol1Hz/M1Ltf04k4S1UGg5Kw406kqFBKy+HUuV/OGTVUwktscCdTOJTEXU9iL1
H7UTYREbD810RJAiXXOY4FRyHNUGVO7kMgS1ux2I4LMkM8J9m2TK7ZcLahxV5t4ENrb4z5nOCFrV
IWWq+OyXmLl93TPQWR53wzz1qCa+ZgWSZF5c0gBB3p5qUql+qtGmyfXuJyAWs6KB+Sy4EWlvvdtN
BQ8GjfyrCWqdhRi3hSiU36tkekyY089PLszFkwmQ8bMPjFRjB5bD0ZfP75K2wt41IMROpT5ChCkC
0iRqeoedElhy7ThFJ1v3EAWGh0UEkK5ScLsBxphmrDCMWks+PdOVhSeCo0T7N5jR9FC2Y72tqWSd
n0lXRe4Eme/qIEfI+yJvxU45/gG4niWAT0VMo0uGKV4QKo159tPqZFRTxFM9R8L4W/Wxr6QPBSDq
+TAyJknciyWwd7M9+GnsW7KDucIr/llfun+YYrF5a5CAuX0ffwn7hc5COu75n1xBC3imKuHow067
+KdnnV9UcPnSqKI7P+Ydw2k+NwgRsWXEdvvlwpm8QdU/icB8RwBB5Bt+i40iILSHvG8v7+cdXaIv
A9ryG1yZ04clqv3vLTuOBrOmNso6bPXGuISBuj4Lsv479lyW3oSE/vWfbu7BztmbjRsciDcC32IK
Z+aDE49DUmtxhTSZgp1VvbSBkd4NZJ2tKVSyIt67TdSYHmQpJ6wFH3VPlxEM6vQmWgo8uyLe2Xst
A9b8kqRllo3HmTbeDmF1gE+eIzOs4ZqzmhJpMVFEdQtX3x2V45p5o2B9P4l9vHjD0LVwTh9DYahy
pu4Kjgy9G+pUyhOJpAD8pHQOr5xFIBGsgX635S10kadmeoH0eGVyxBaI65519W1s0YXzjMsRAqtb
c2BZlEILoqwC93VKy/YOYiH3faYaqehMV9Ire6ETN8l0ydmxgckqxk4S/i9xTHiiZy8IG8+FdIPu
CR4S9kO9EFTkWIwE/koIXdnQQfn5P962JmDm6sCVEF3HFpCbyHQM5S59COfzNSrABpUGPFVaTsz+
O9S0B5MBP2x1l1QBKKGoRhsBSsDRdpEftzNPZA2oXqdY4XN2f9NZEOjeoJYDBZoyO9oNbDgUw0qO
JLVJzbOV2TCpviiP1h2VlTIhEvRwOz3k4uZG4A5UeAoCnX7UQhttotG4nkcwYV8rDoA6NtqGEwvY
+nzTLtXCmZ5zkCeIIxKtpLhjUNQKzHB982owabRnMcp3Gz7FaDYuv9oMHf2UNSui//yXapehSjrO
7wPScyY7KqJpTSaM7iBizHDRiSsHiL7iWxOCDPk5Ptc5UbDHvLfEFoZ+lub5gKHMiN9O92xb1tLL
KL8k7MYakpntPeiWwHB4bd/Y9vW7TlSIMyqqHzf2hh++Y1szjT5lIukDYOc0fNQE6Tk9aAIGcmDT
0bDhRn+Z1kQss4Glza87nNq5gKsmnIoWUtk31lCooyzAFrmYue0qYNQA+qX/hVbXQxxj38XCbhpX
H4HSWDOuAdM4CgDEggSzDB4whUbyok6ZvrmmtGpqDAFrWB0suQmbUpMch+wK31mgHgtbP/NMDjVa
8iIvAipuW/hCN4J2DlMRU+sFqyDOVZwb6eV8JFp9coWG6AJemK1I63xDgdEQBgmW4jVcU5gqgMoS
aY3WaUVutN+I25saBxyXI19QNiYMkJPUtqEL7Y4SVJkpJYlV5McHOYsEKHGDl+PtJZA9e1JiVCud
rUmy2pB30gBd/gA54qKtBQxS+SyoEV/9zyMLHqXXRzst/AWTRyR22RcVojbXGeKr9G6AZYdojNVD
VJJ2dsoOba4zqFFcMg8KjjJITZFd0/BGSdMt3qT1H/CEg++0+HajBzE3S2x11rjzTLozkPbiL6z2
uDtnbCKYJXA+FzSq/dtg6lscL2GCDVrMW9qKzh/Huh2AVTkUqrWj3NfwXyi/le7aY1H04fclemnR
EIHO2B0MaIUFlNtQUar0d5sX9QKjuj1Inkmg/B8UFLpqdUyv+OunPwTyChHvvGulpMvSgpqPoZ+X
iFj0upXTk8vcWyZwC7qRB6Up3CIyqhhFphyxmudiXsyCQejFKdYPoOjUYYw9NkEXpqmlug4YLiZw
FKr5zUtv7NYpEw3MFralFRlFGHSQm5iC+0EvJn+XC9T8rsNhys8z1UdcmVm0MWgUnYbnqRtkyQCP
2nTVEC3waENrHoQmKNOHWiBmeZtohq+wtvzYy/0WxaGNJHs1JgGwGux++Q8wB5NZdG+TOcM4XPHA
NrUXhdZeAiTYgsPYq2SfXJ3FPAkgdx7vA6zc7kqazmmQXXu/ljNmKCNOASPAyuPbeIfXyBHEtLgj
tioIW/svVf609Td8DccsWZa0GfRncXoerCu8X/F1AfrTV9BL7wPRX5U3hdptTP+OS0ZnE0D1yEmH
4LVkMcqK/OL7XRqDtdMAdzGUo0m/WHuFCXhCwrVByei7uRJQO6t9QWQsDj5KDQIru+NXJkT5rpnX
Ip1lapzBcvVuQguNusITRkY5ovGz/tWDMhmU1dL6Bo0NSBjbAktal9EyPK0ntx67Orm7gpFnFpL2
AGuZ1tCsAjNh35q0JFchadxFwqOscDxaVRXuL9YxdV3VRM7i4JVCqY0Ac5Uyp59ddWLxOiVp532a
Prm0Nfw35pf7SK713uW6tx7ZPvvDUy80dNtI3AJ0uKkfSd/bqwSTQVnpuPKAa3ZjcGYN/soEsFcA
bKZxx5+x2NTwlryRZ5us+lHfEDzf3OmSAksgZ1TRqNrdA4er1rwztsKRXWPTHdUdCEhiQ/O+QZfk
2jMVL3V0mDHE6ez9k/TLZ6j+jBYouMBCf2DE+9GT4ZP7/CuugaCB6X0ConPTVviGPFMKBSiXuBKM
F86d9/aQCjNKEV3n+AF2UnRzWokGwS6+9LYKRIF6Gw+LsG3G+R9lkTAZd8BQRUFNC8dHYdDA1RCx
C4UEedXfOoOQVWs4xNa1j+YeNsxgELrhDuyZqMoq+VIGXKbSTvFii7sQ0hnEUFp1Qx+6GlRyLVWD
WtWBTyw+f8S8b7eDCjw9057dHx8/Gnonjy1MAZUO9H/tev7jWDjX43pYB39ywt4X4+V9SVC0gsTF
iCKM+ItaxYcl1HVRzbEIBiKPbtC+P0kg3Q/25pL++v0lGUpL6vqERe+LwZhvIRWHLWddqVM/g2J3
d8jMFAJ95aCIfYpMEoiEV01eRtwJwZY7gg8RpmeT6zbP1Zg4LHW5yYfVdVPHBY3EfMszL9B0I+/m
UaG5ezO+fo4XONe7hwkG23xJCsdA0O5rjcXAddAZr1joGswUSqhllHu+Sk9vugZXBfBRik9D6Z+k
wjbfXGPev0eGd+OOPJTy8iBupv3SXpUbsDsIrqaDokTpkoTqjtQyQP+pwoALvJ3ypT/TJoR8CwfD
t89eA6oUavqe92A82uMehIJl0sP4f8kSncSRgV3+0p59QgkqhvrL4jwjoExNmcztw24gQJseFuuT
8OkL1Ag0s5p1p7xZf/Jo6iS5Ozon0qXd6jCJUssnnJlLEfzAi4t/25K/DgCk3azw3Yhjrq0NWkos
vsSAF1I+bQjtBhqcezMz2v92UpTVTq9Wcp1kpr0jbzgUn7e9FsyTlSPDb5ansgitG6RJlfztuL+d
1zo+8kMI6JGUAO56g9VWJVESachP+xW7MlUwEacDrzDiKLwKRUErD5LGafSbCR8TGYwZfkLRVfKt
0oqtTLSbuSmsnnqzGQVFHcgZOz9GkmrtkcyuVvqgcjsgvmEwtzstw8CRB+NWhmeGYTF/SWpxEZtf
whsoHtNK8yUQS85c5GE0GeDvNiWOI3d72eG66TNFyeVC+iWCaPLNe245r+27mrcEr7z5+DFM0FO1
SyPCqxi1yThGj7/d2cR9XGrpVjsXfJnarV7orXg1Dkk0F95p61BcMUMvrFzsiiTrPmXtH7YyIvdf
wCGroXcBqluL/JfbLHHmG4Rl9Y3LJ9VwHJUL5peiqWFcuVohbO5XYFEzA2bh6GYlJLNr32HcNwA4
xzPj3bNvS5xXKl+LNC/q1PEfbjp+xIhJPzg1zsyTn4DdUJkUj4H/6cEbvlQbOk4obbNKAYieHbd4
4oOaLRfDozJ1tBdZVB8zwvtW5R7rPK4fcktOhyMJ+Lkyaa6XBQtMdhqti2EevJ0KGqMRuVDo961X
YrtRAy71+fXPeU9oeYMU0jMguembxBERMtA4mpdy9/hzlYNaZUVa4uuQHP0dLw7VfQkNEcTU2g1M
P/MK8fMp4ZUnOg/1B79ihZQg4LYSjUNGgkQPt8IYjTYEgrxg7ob2tiBC5Hj2nSwQT6SHD66zTBhP
1TfYqrK5E7aDztbemY9Zwr54762eXdSfFPadR5hfv5Abuk+0eMqF/1MI0Apa4OlXMZL+x3ferrA3
I83HRbYNMH1kyXGm+ibAUgRTHjQVlgEvJcxPVid4bCmhuFg6Ojoi1dk4h+RaET+0p6BJd5506lAY
mlsC8ep//dqjpKPeR5KeAGQvAWWo30GF9cOr+7HUlW4KnLziJKmfL3tyGRY5JGXLhZ8X8khr2DIo
/8l83Gwt3u+LFEVdJ5bM5N5QSO4Ur10HTuiGJEC1hc9YHSqhoHv+/jGzlMeVt7M95M/2NKZyTn0Y
9sARsp1NnWwSbSuxdiVlj96TGj9DxzbHqjHN8Abv2tCtS9VSMhZ+RvUqP4zGODpbrfFpoj13NYfX
4IMQKyg0HsC6W+Bbtlxtr5gwCSiqJ9KSWF+QFLc7P75qje8sBKUHqlNyU4ICi5vP0zQAHJmK6/8D
VIgHA0Es99kz1KaEoGhWOyWk6nWNVDwpUHFkmWoQZ16/0B3L38WAPoyB1YnepJ+LpnUdoPg+Vx5k
xtlJWP5NlOChPt4Zg3P38+WhTOXJjHZ2+RAc4skTsmsG3TPq0YWSldlIr/oisiYbZOyiNZsbpBLp
w+KHYUTXxF3Hsh6RUw6m1x5+rZ2T8OO4ZdP6g9oOPvZi3CCw2BGXVZ3VAvGvIg6nNfgcnwepiFhN
cXPzwJwfNwFxWFcGV0Wpn2Q1tFJfb2R2ByzUuMo5JCheX61Omv6UA9PBbrerWgSkA4wd7JeO0aS/
BfpEJ0NVumWaKzmT+VeexD/LvLhcjhfHRjDLxWaI5iwwuNHUEFbrPYFEDKw/8TbT+kjvEX4TfsS3
VkIerTqJvAwvoFMNkG/+jst3qMW5dwpdbZPjmo+4TZxkeAOexnLwYH2AtTFxMUl1bzPpl2MhZoRw
zGBUrNXe2CMTX3iqNWfOTvBMyIrr99eVIfNpVtu4RcSjt0zIkaGZ9w3KsQbtBw7gXf3xKrSXCMPW
twv4k8olOYi9wS418e5qKefGBr86VTRlZhjs4djJVLoCmrjU2Qz5d5UXNyjaq/GJZKiFsuDUsdzn
iV4zi1iPrpzne79opykqh6GucCQPmNAuha+Dk2uZ2Sir0GDS4Vn55aC4R15RzndC9DDhxKZo7KLW
VLnxutADnK3g5p3rjebai4CC86uS6ag4uUkEXuS8QptlpPH+fs9xfY5DsdmyLG65dmB9+8Ke9vsF
4OhEKfIphUxeoMUtFAKX6WdbYnkf/PzsvuV5xWrZsEC5J4JQm2T+xaeeA0Hfa4juNk9MZecrnfwF
2HE/l0uuRjK4rKe6tm8iIWw4c+Q9/+ZVrtpT1bcr2hgGRL+hR9kUlcnNmxqQoIhmQZXWZCx8E5uK
Cuf5Snxe17Id8Mbxo53Sn1u2i+B3IjkzElLI5oH3bh0osfW2rQFwaTjIRbAst/rS89Dhgv6j7cup
9mWCVK/E7Q1yvWv6AyP2jLeFgLxSXS4xU+UU0QD+Rp113xegxoDwl2Q/7ic2Rm4vAY28gzqPhCmc
zQiqhNSy9U/MVWMfaSjywpDMrtj5i4qZXorFL5kYO1LHFDQqMI9sF71lkAIhPl/h9ik2f6Dmtl+h
tAdtcnVYrjZUgsC3ooL6P5qu928yPKI5jlHmmnwk7fOsNcINJRiAh8txE130fURLhhEgvpb1E3aQ
C3WQ1J+e5NJTsxvo32rH1d0hFbWdf4V8uZSP1fUFoNjOPh0TGTqVMQg6RK041mNz7v7SPlD5hT+4
+DNGTzLmQrxYK8YF6xwau8TfnemH6F8En4ohue7amLXdzZ4qI1H/JFt3FYGknDJONr5tchHv3qI6
1MsW/r9so4zP6WPjiWA6A1LSCZ9IyVfIIxumI8h2NR1IPfwl0rrfrhDqzK7TsUbJz+tT+OIEL31A
tqrsn16qOov3Jh07wCCyzCf52EUupMAVU35UbX8YUxP+/HRhdXT/W4Qxq59RyvzH3xtwNrDPWde0
TE6U+NIW4E8wC0BSnmneU1Bo91x8YjIj+JByfnpOxtdS9xVoqBJGxrtG8Z01klKCah7dG4pdbt4A
cqt8Uru5nz8OFxDACPNMRziP7grM1vxzArwmwmvMFEdkzjP3N8GfnQ2B3Gg65GlCmtTu4u349Mwh
hviBxB/2q0uXR26XJbfJlU5Twd1NK9JYaBBa2/lT0fLsfS8VrGmlgUcTONSCY6fvyfQfd1h89iwL
Od7ILYuQk8mYh+eERlwQRXwmKEIyYgk4f1OvghMoJD7Dp9HApwghCVFiZFClJmU3eNZGIrwjXhWJ
zlbQlZ1qId15hX7XSctbYPx3irohXaJZ8g7PLqm3HYHgVBv9MgHZnRfVUxOfEHQI2CBkeyCl7PQn
5F6MustljFeE6iP0MPu4KTkmWSdHG83wpADLiVrvqPXsvvje+t9AkRTtMOlmEZbgl8Jzt5OBuGk7
PJSvjR8PhbFRxgvXjuoSHNXdLtdKFtMKN2KkILynhavCBkHrplY8rLatztTLJFB2qeuyduJevtqY
p+o3sMfjIoYujqDWV3R7D5t9UJhPrqYXTzgXrCSYCFvWR1PTHyvAWNZHC5lpRUmaiAC51fenv+Q+
9J5v4z/IHETqmL3XCv/EN9GM6Dfd9LVxpo9fHxutbNH2K2BaHA3QwpqQE5f8lKGFAKamDPfhXq4X
xzucqPNkYMSjVYvUM7Qko20Xm3b5JbLp2/UEnQqS/hoHBZM3Doo1HL5+psmh4n9vLjHlUAb7V62+
GhAZA5ov+lGjDQH8HIRGWde92R7L39hetN3P7kVjqWNPax+tU5gd1lkb3LZe5AFFA3IofNJ/11P+
1SpiokQo9gF7kxYUKBWu38ZiBzHO/eQf6PCyh2L5TPY250PO5poz5oUITpUYZwPR7ag94+/7LLQa
M+UHq+QhpjvZ7VBxnuRunXBd/k2B5bO23lGzUXwBPzlcrWjfjqA+7aSxl9w3ME/k0chO4/fAka9j
xJaV/ubm6SV7lSdM76YB579LZlHBKACmxpYKaELZN4M6gqLkzPQ8bQMhLaA9AfgqZraUVwjgaEBF
w7D7OXNU5gi5WmdxpCexgvCws858YJcXC/YkZn3kmiJRkaZQYkyedKRV5bKceRFhn5/6T2ai5y/x
ahMv7DQl6J5hwHpULlnD4kUWCJb9TM2OAwToAd4Wx79bDNC6zTpjqIf5U+BIwPAe8NsNm9ABDHlS
4AJw42rhm/vhD1LkTGdusukXE5wl0mHFhN7AyTSfh4IxMGgaNRfRcJuGpcxEsh4ttIG01mepcedd
65KpEV9b0eRA04CzlUFoGB2KgD7ISRngfkjldcx51YCeFAnludvqJXTu2I6qkkYcAegYDen+GDYc
vL1CuGemznL47mfcrTvOaVCac30B3kanbRWU+YFQ+WXf8URoGHlbJpspfq0LdOk8z28GuJXljPgf
ZXI1pnLP7REepQNacBcTMy7Sx6wcMvmhdk6s2OSPKvvCtin1+ievfOBSrasDB+ZfmRi7WyNPFYWo
0EoKYfOwFU81xUWZ9vOv0Ec+l30nrsKUl+N1KIfeZvapPnDaDxjUvL7k1Pp9eI8Zp/1BqvKwhD/g
9I3Asaw3OT+un3GfPg/m1AkSiLYAQHGuCKXpVOFcKkAgMjLHTCxbJ7Y3GfUppMvwBk3XkGCZ1Ro/
mvM0NSvhdtSXnwOvcDajqewF+Wp3fLPSqbYalaa0Q4cfx51ynMwX+2OTVOrpmOJ5kIAZTncbCS05
Lv6LPYoGfKcRbcmCbFqj0ZS9FGgpCAHk/ClZus+lsXoURE1HaZFaqPXiS936k2GjuMLLyJZE1tKH
eX1ezSRFK+gCtuzoz5dOG1rtouMfG4Q2StAVUYK94fZHNLETAzTXhaAWqd2lSEpi7PYyKY5EtNNF
mqt0EF+Odd8opm2QECv0mMGpva9xL8gQtbkdVCG0Onm26k5F67d/zKIm6/kzUHTplvncPlc3iyMt
RgCUT80TgUwyQP6isfVsCpm7Wl+QzadVYtPbFPMDXsgBr2GQqhoppggAdwHe85pZUuT3h9vO9xxS
XXt9aBbEh1jqokp3vMKYeqGgNJrXtwFKFWvDsy/rcp5X2fz1tzh2ndBDdClF+I6N3lYTqX5HjtfT
ScYbT7/4TfTkFj1a+CyJdxS337ZN/wiwUtzOACDkKNYmMnr5f+BmF+ggJoUm/3xlx66y4Ln/t6fZ
7CVewBaY7nvZka+GEcn+XGt6WUUu5n7fSrNgoFHuXAc91byOM2RS030lU5zps6OBbNAykg63w9Ov
zSc1nazCsntc1qh4V7WBE3HmX7Hxn03eWjC9b2TaBvEwfnfPlt44cX2E3+RH1ZoWnbnzfwNqNgj6
JuOqNVFNS94sOIq35GAcIif1K9BXRKG3IoQu3DWI1FNwp7LT59FCpfOASQoG6/Qi8m2FHaZx6lun
Mx6aHNraSEc6x1VMAK+7/qCFnMhiLFXzDy2eFzur9sY3V0XIsQHE73SpGPwPdFypH5OdfAaUealw
SZ9sdaRTwryN6GyQH7XGjl+Ptj5gatTuckE5QzNXeAcfKrqjQxtS3H9NXoDYU99xpTxTytAtbAY4
32U5KTpSJEqohcDkAiyLiiQU0PEL1fVwCn8+yC0ujxdzap1qGBIYI+qjpEHWfIJyXHOKkbUNDxeN
2XLKi5AKTShUq6BWr0syuDAAqSEirbI2TmnKcmi72N5jICOzo4kSIlapQY9nrvpwRT2y4aRGHPTT
Fsb9bx2WS5lgHM/bfzam2vHwTNftqdbLEfIixKT2sOUiFeaVp45Rw3/Dsr/FQ8SUFXYOSjbkeZGh
MvFLmsuLHgiA4GSkGdEwhEEe0SK4cAuj7HIaJ0Nzx/LYkDjuz6pwl0/u0SvEdfzXj/LhKVV46+5U
QEu4arRAvYuIPj8QpbhBFuKrB/wRH5QnCvQZ4PivK5P8tg3ZimCVrZkGxyvf6UgyutWRKQMqtMYj
3jP583ZqW0ma7JAnWNRB03Gbgq7UdV7b0RegzU21u7x+P+7JlGB6uxzjzVyAT/MmWoeMPF3XmUKy
A9JNmHCwdMa304AxYja6cifZIZmCYrqEe0u1I8UQVHVjgK+G6MTnpu3WlArlWJCv8UxjYgcOSmjF
6R1LfcU/x3Nz9Zx3z6rnFss50R7E4Fl/uGLigYPWXO6ud8yv6Uyty/VSwe8lTjIIIRXRewl20wSX
X+4UmG//ezfgCjoUt9noTbTU8NLZDT0IngQcGkxyiLJyrTIWI44qcjDa2vMYCoW+Bbw9ud03do+/
lipQmWQLai+k7wnqJ7ADXW/zey56gLfuVZAkX8UsjvBkias/30vrLXyIXd8bBA/r6O9jsbMACFmC
AaXtnXhSQ7uQgXCuVOxT3216ajtCFQBoFy6aYYnLl6rvCgwTEqCQrjbGDblOcCqjATPuene3oZj4
iAAE11GkMNo3/IdWQSIvDbDUSvMJiDNXHs0g7qEjMbiJQgux/HpBTwm/Tg7XPAs9idTJrEvMPXb6
7MxG2xr0aFAx+fuaJYbivLY/Fwsnj2P47/39Id6lPKhaREq5omp02spBOA1Cf+jeIwvCLXvIH7tH
63ijtt0PGBHDd0uY/6Lc053ZC3Z0AqVgXF6W7gUK72LoahQyAJF9AAmP5U9G/PMF2v2+x23Qj7em
Yq4p+uY3qXoQY34GBM1BQKjQOVglv4gd783QsZItv2j7LWUvOpCqA5iFyLML6we1+4ZlCo2wKnn2
kf2egtT1ambXH1ZtxgHm2ccVKfAIt7iwvWjHQwO9dgUberh0Ch8t98LJDOgwXr3zAhGAaRzwoPYR
fHBBPNHiA0+xiECVNECTW7I0poNSOO+/mAaXfLUo79dlzNN7oFPgbxV1djggp1hRP5WTC2kaitgE
nTfr0ghm9CtL9VjtDw0nPLP7HjClCnXRIuTpbtJA0h2z+tKrSvj6B+ZgNgf+vIabbR/Kmj7QDWMy
Bu9wfZUbeYKi1iX+yef47xpScNVDrobomRN1rzuX5+0gsDlHGkTsGOTmmBE245h0tLPI2sm5o+By
s+k6qe4idUcazVWxoF6t/0+oiiSZo/myAQvf0qygV8qqbFB+6UhgNT0Y80uWbpmC9PWH6mn3Dc0U
9kPTpYZjkfdR6s58xP71YdU9+cy7NlPrR9/qoZ7Tuv2J93Pytru2feCvyfHbTfnTxdl/MCSDsb6B
6YH3PDjqxUqMKO1U4EDFzq4fsOJylbjteUDw4UhHx/sXeCo1vVqEtPbH71+vH+3f0LRhhhXUIb1z
+xNi/asN+/ms1L0Ze8Z/Iq64ahDQ4GZ9nLpfMQFa8c+cj30EKMILRsAGX9HhuWCcZJrIhuE30f0I
LjVpCEmV3lrVXiGPvEBqdqphXygb4vLBRZrXZ5KEtOIkySHmmd9aWscU6ulgL9nJDK21icLbFs1M
vbb9gqfVU/1oIaMMlT8sAe5aiHwt6oWKmoKVO+akArZWvoeqBm0KRoSazuqGV4nmpjqq3QlQ7fDE
faNe/7D90jtf8wKWlAtkXDZz22m10kSGNCb2duQ+kPCZoi2jULnE+PWc/O5m9Eup8X2SHqUKQemu
JdoLqghlR+m/5kZgmwB9SoS+jWjk0ccRmqzyh/tu3sWOUsFxJg22ZOjexvqy5fvat/kDirgbF/Ut
rKGsj+J+xW5B6JC7BR6DWrutL0KZoiqkOcaeDbo3GwPlb1Atame/LMhujQzHGQWUjlj7RqhHX+Bn
uZ9RYBpCWGATw7eH3fwUoimDnjqyMn//x/NMtVHIPMKp+nZZdW4RP7ilWmfg1PpwNUcxOLznWwQr
/Dea/E2tckw/4xxI8YGU3eTnu4uuigLZDqpHPYMJfSZw8IbTb27I74tjykmdYmtCvP6AB5bBnVRV
TMoHJHR6F3+DkQb1WaXFIW0mIgMS0JUlQj3/pW3tw+GB30xaj7MLYiNVMT2J9F0T2uypBQ/zOWMu
EoaYX2bSNqESHHoA7bsACN3UO4IUFWrLTX8U/kCInSOeLk63NtAHiSvAfyo54QMOAT2t5tDDP8fO
oTkXXmqyo9d5kVLel1FDdoGFhL2lzB6afKyB31Xw3ksOR/kwlAd0q0gD9IDOg7Ge09c4vXYd+PJZ
KrET+zDqACb8dBLef+14hVoU2tjuvsamCihhMkKzjbM9jd+epU8lq7HEzSuMo999YVtBEFrYoLZq
+qxRB8PtEbRD3MSswG4sOSYpZAzfSmrM+Xhenej20lyrcVrDYeeWmj6cK4z/d2uCKp4Yny51Di3y
I0tFviznnPs3VCHUfgO+WdElMuJ5TAkwpaRo7qgchD9gVRKp0vPdgHO3lKEQNproh1PKnLnFH6H4
DpDkIJQqmdUHvvJkcbG6C0dIJv3LE06bh41uW5DyLzqFa3iZqP8EmyvOKm9nr2XYFnDeeGOZv1P2
6g4DpoAE8Kvxy64lL988H8ECki6svH4I7D8W8/i5bReDvZ73ODlxK74qewG6DEf9PRhaNMVRXRum
e3SvRgGz5JaOsaHT6VUzcrviMddt/DRprH9kkrKyM7tf0GwxfRwv29FaTHVmeXbG9La0wQko4Ogd
lb9IGO/ZBcXLpER9By2BCF7GFrMNSIo3tD3TZGsfguMIEAHgMQtxKHQ/wv0y09DUNoS2bwXfk2rv
FscM7u/p9/2CWX7u4jFDbGaVflOTv6P4j7KRHXM1Zo0lInqmavvLM61RbiHIzXQ6gU6qXAOPes1r
2qLNcG1LS3T7dIXZLvX6zLMZ6S/pwsnTAraojk3yk9+4c5kpXs46T5sg4RqVRVT+1Haq104AsD0Q
XbRoSCl7e1ffF7ALmFfGcx5cD7qveveB6zkcrbVrP1I3wst1D/X8AygJ90BGBLZuNzxWyiNjX7VF
wGCuY8WzMBy2JV11a2FLve38NA8WWlRCnwjT5CoopofkEyX89mxKKFVuyA/v8KLUh786JV6UlKfT
z1hoCzLmgrWUIgWw3pNXolHPxef5hpT1gOgA/Roixks5RO0kOTmOdf0CbNrtoEleFfMMVojG3kqD
mFVoYeX/kArbY2UvbDkIw9DbLQyHLcyhUecOkZqpqFrMcDkFUyJ5XoSh+yLKu/WxSyDiSJiy13tA
idZklbCrIkqjzWbKSfS447/ULeWVmAcbPuaaqWtJyYybxgtR4NMaFH7wRDlNkbbw7P0p0Uah2pXN
S+BAKbbepECSlqOX1O7OK/jcM1Y/WOSWVcdHEHHbBU0l07uj3xC6NmemcoZmLbA4mGHQFCLar6DG
HSCvShKlol5Wn7yAjqWlPaKiOU6lLpfNiIlU5YZtaxS7ol29C8GC0wuuDWbIX6f4RksFI+1YSigC
NhStZfiPSavdOTTyZv16AM8k6sgS/VyvGs/WKv20ponNgrKekfQXKFQle7HG8t8RQr8kU/Ds719X
d39iBTtQV94CLNfxVwn9FLyRWM/u4LINLnAUUOe2QQzzINAdz+rHWrTjDR/1VwTyQkxoIMg6/yVi
kD1kSx6sAqQoc2T/kkPRwZk3LZUf4M2qcwmqkw1EUF21YzzDUr24/BiM2hB0LJFDWyf0mgIB3CTr
qFxfiz8l5i4aD+3Et+IeV5URtZc0AS0n693fkMMaFVexAmE2PI/Ja3eislH9JeiNCMLQfbE4NlS/
2oUgp4KugwECC4iviflYISQNitGM1BimdHfvCsHq4uyjGd6J8kv1VtkUYC7FvjfTixSrP5ez+nlU
Bt9+TuM5iSkNWufSpCABYOdesQWct4wyeW9BL18xmzoGIPRm9elYgZuysNXRcYuHhJBXBNnO8piV
2UTmEVVudZILggDIOoncDlpFlEgEIEyMe253tX3Xqo+c+HUngPt1wvuMidk+aAtYs8zbe1gOd02Y
cVLnUtqYlBTI+iPJwFhkFiHJk4CxJjnxZgjpM2AuUaet+xuYJJHAg8L/TGY21v8NRHiLuYkUzf5h
Aw1Ogqnxt/uKLV1TjPc9SsjfQKvAA0qszd3+BNOoOQAX7HQwEiRI6ocunAKTYjWL8UGKfmPi2t8I
5KaJI1Iwtg5f/yAcyWNDwyMHKjp3o7jVm6yPHL1zf9ypPZ7/qgZz70gxPUbN6R8mAOlOTjm+pCG+
8DSXdcydeA6P/Zr47MORIqhwVBzxyU+TmjqBuz6F3GP551lGBXJOEw6T0mctZEixXp3Qvs52ptaP
jVhKbzhx1KySIEkhwA8HM0yZJ0Jf5BKnQi8vf32GobibePTyiBlputbdUWZJ5uVEeIg8GggWAXPP
zc97ABCs0qCC1Cg3DBZWMKi50C7o8tXBThBBISXA/VZCRyvxIaeiddUSbmg0YSp1Q9nzGnBs7FIB
lPsiGG/5//nTQo8xkLSP8c0u5840sMOg/sdB28VaLf9jQVbwGS0mX1FFPmK9ceQOISz6KvP7Jz7P
91DTMV1BmbQPBFnSXQrjtZonNFkJrM5uujA7ViumGrIXBXe3xqdzX7mTkbEe0fWSfh3bX+Mp2Nf4
hg2Lv4VBS+EP5mgOqcegZUaLAvvzVHAkx3SqW3hzskycI1QdMAqD/wbDj/eMq/1hJEi2XCwxpD0C
5cgzGSsC9iGqISOiN32pxfcr5krutUg4zmB6+IGWSo/Mh/80btGC6M84n1WlGcjQ599Eigde40Ak
88qKp8k0HERqMeaM/bJjbD6Kddf0b+D2CcMePI/5PkktNP/lEuhA++A6Ap+WpxdccwHF17zIvvY4
CmF0XCZxH6JiSmhUCH8Iz+9Lyc6gt1Gw1i8oc+asK5MDiKU3b+58CLmfk/WE+vHy7y6/3zevY93n
gY8quQb+o+KEQETzM150oK6JSB012wkTNXP0awEv+qWMGak+h2Aa8X1ZoLaAwru9L3kXcvHzz2I9
Of2bHFBdl95HeBZCBMzGkEY1MVGzCWoqkZz2NE6pSCbX6SXZ8063ZKJ8GpsguIxeROdhtxacnc/O
65bJz4sPuULsXf28b0Xfq8qTlCqwsNpbbj7ODI5giEd8PPf46CWLaTPvfC/W11/kEJeSuDFRDn5y
U1AUwAJ56oWyh2toSuZ9Zh9V8TMElzO+aFpkbA/nUEICJc2ob9xsyRnGCvFJicO6PTgKpZHhaQi+
b8vvd3cKqxHseY2cL0nyQZ919qECWRQIsHDqEFrbxn2ulAgaCl1nZzQT6L6xQeFNJ4CZ5AhKdXFY
cnZvigNN3oIICFXYJ5Ohe1YCkWSH1Kakt2dvZeCHRY+DGhQJiOZ70j0rW/lDUY2nfHh+qdX9+AzA
pbYQHOIRdtaU+07dG64lDtCnYIMHeyYzevuxoSPd383RTmt+vGaElKRNtGGFOMCj7+bKyHPTtkLK
Li5H7g0V0Rotdm6qdkgvdLfscRFWqT+oZhxe0iiSnIPVLanoww6bN9qUdejoA1ttybIGqJZI7Phi
+szxPae0nyvCwaD36xKJ7MhtYwHak2ENKpXMEyWU3MxKJHn4o8RmEdgoQiUHqobWOxsFvTfE0dLm
jaT+JAQRoUBKPvLshhTsbmQXAszp0BJ8b1PHJXnHdhzzKOm5flJf+68aCylsPxozqrA54bw5w4vU
IhneJeQSmw1dLVoEMrfzhNX3QoFdHpEYdBharrlVcA4F4KYwaUWKEw1y4k5G21HKXASZ8U1jY1FN
tbXl5XZhbLrgFdN4p8yDEykZrMDSBkNe2MOa9Rqa8zSzXDy8QIr5PNIAI5eYLVT1iEsUzcsT2cpA
9f62BkCCN0HeSljq6xbdZkOZfvPO+9Vuhlh3zI3XsLZ3cD3ioDF6cQpvwyPY3sxDTNfjFuxFG8og
+HntttLem5kS4GDYbfQWwAOvEDfPo/QXM/nQeo0L0DBxb0t/5Hf+JaAC1CBlLRBONfHS/x5Ececn
RUEGaoVsrxteX8HUhCCVWTlynYSfx9Wahvy0e8tuFJXpS5OUZMQWXuunjKpJ7Mlg5CYeZuxrVoY+
AnfaSNRqcMt/HYYdeT3s/h2auiDFpa2Z9/0vnT2humA9RvMmc0z80BpXT72VahrIO9/KuT1PuA1o
NAwxsdLgYmInjwYkIIkH/aY4cZkTTRpf5OUCIksHVZml257UjVqzopc5NXpcjA4w8sJYYqA4MLKa
IGzrwSg7s0QAOONeiTsnRSNyzIISxYpkj/BvrZRisLFP+P6NK8lt0doA80LvD5Ak7tdwV+o49mKL
jQ70v0Hgn39Q/TPtdSfQhkSWzcbpkq8SYwUMZPgYsWsEIwrTGk8Yjs630cEVU4wpRwUNhvTijQcQ
FmkNli2O5mb0Ig2qNHSGQNyZiAiRTZbUKclGFx7WSvRP65LN/EEiMpEbDjPGugVOXg//5oPYJf3V
cXUzUDJG5/iUeoi6nj1gSz29/uQjeFgdAPqDl871qLY8DH9T4zjo8wfyhTgVN5WmraRIBQ6rMLEv
OC1PgzsOlUS1x6HY2tMJTJAAwVY9re2uacYSpRz7ZaRLEk1iTzwxDUpUus7hUyg/XzPy7n4rBXRi
0wCM+Dr58SJEcqfZ5t8D8/IoOhDYaij5BqiydLPZqYZ5nNrwvgzFMdfHpXdsPPLZ0fVqTjxsn2ea
vPrCxsk7cSBfdJJH25SJHzpvNbLZi7C67hVTfJTbORxTKay4sOQWve2JdYT8dHFRwdTVw4QXgo+q
7hlNFTO5h3hHs3/RHM7n4BRkuI4xM7LOqPCnl18n8MgW0Me4ATiVY0aECywfivPRx6U5YwvtpqPg
kGLw8xOv4V1GUtgm6cRmP97WlSnKSSIkPDquizcItkHVgwE5oMigxPe4JGCoVkAk4ENDPqUKJukH
5qugqRhqORaAK+No4NZatgnqTQ9lV6eRjpLjhMQ3GcfaxBi8jh8sE95Gk2zUZ6AtpowCd2SWRsQ/
dS2BtBaQJbbPdyWiHrmZ+tmutA2tDyK0bCESFV+gC9cAwOMHRFw5uaBLbsZeh/i5alcHlYH4NpY/
9VS9e1A/V6Rf/jec3fbgOs+0+DL0yu/O6aGn1PFtJo7N0o05zTG2GCugPhESqGHSCGqjLVfCMai+
K7jwMxsY7iXnAi/noU/9WCRFubGG26E9YuxhkVtT/yH5KbhtvxKovha1OI5Y3dLA7F1CPI8s3S4V
ei+3B1+2KNIOrw/uyRa0O8h6Whzb7CEnfpz3cvLGEnwcbPqig5TEcb9tE0/ySo42Pda9YG1qekVF
JSLA0SR2DQRJcm+lflUblbYzGsm/+IXYC358/xoOs/nsnhGJti8tOU+rIBON6vh9DtN+hkJTwHPo
YIe3b1Rvbxf4gvxtYL5NbQJTueaCO1zCmsJSecIHNV6KYyQRscRinfhWkO8lVNZwqYtdQolLUZtR
u1No/iMu32DDPaxl8obQiaISbXGnI6364bwYZIV4xwExFqYkcxAt0jeY7DBA35tAE4qgw1wSwU7F
zQ2taKPkAM47tJvLN9HtB+bu7CgS5NfxKTYeiANw4boze+PWw9T4iD0HMZkWT6bAwmY+EAn/kHdA
5cgDBsxemWrB/4w5/XfAM7BcZgIG0mQ4Zag5SAkElRingcJ4lJjyIqRivBFQt19RQ8/Dy2lwBmSF
Fz4+9XBtNEse9N0sNg+Na3US2mqytv6DgFvuCMCjpgUwr7IXVAbNkr3k6ijjn3zaoAXMF2lRtE04
r91ncXr7Be/rsYk14FpgSCoYDUHswFnFPjXGUEVu2x/VrTVlClVNag64kNCbeGLPPoqIGEISThPy
eFb6hROteKzSamkMrsVyw07WpPc9C+N3Qcuc0oeTM2rd7rwlkQ7QJ1rJFT9/MaK3PB3XeUX8SwNO
VAuHZc3k6n/szNFYfFd5sOGzgYY4tOsYnWbY1w2d82T+cmZHr/35dNlsOzDNkTQ/rdQ087OU5Q7d
wRxmHl7RmwmVu3WcQEtL1peb33sNXTL7/vPS7T/StfmZlQuD7GfBbRPB+ig9jXJ70w99LlPC3DRl
L9KrRx61f7SNioqZEW0kckQR4BJWiJzBKTh97pGEvNoekFoP5SeEvTFDdaqSIccYg4rKv3N6QcCn
X9jLnRXgJdvUwqWXAPtXZuYuuKHcMTCrX3OksbmNL2/MbRvWiKbGu3WjAy/hywtDlP4i3FPNbGcE
jlh2IPW37ST9tFdids+RRnpbdr28Io88dcZu+/FOJ0dtRM0DfkoPpKXoebf3OZwXPBPkJUfQz4Q3
plpE4sp0t1mOmcZ9YYbgmB5Y34z0AYc4CRlDk7o4sclp+S5tDEVHQuVMQ5OjK9fT5yLof/h1k2K8
b66fhF2N/hC+yxPflroFNNhYwA6XnT8gqQ9+eYd51GnMe6jaci5ZfR7sp5KmUrD6QCJGIDDVK1lZ
47gxxjrwUxSU3+sImwHjXcd4Tn0SEmNFv+Qc6dVASP5k9cwxwxT2y2ZLrgj23loXSfnvToEHRpnT
HHMcd4ZuSumlLg+0BJ93HeFBLXAg6z8aHKFCYssbrJjJ3CMobQNWFWgT1BO8bEM7fCutL7L+Efp9
cv98gKICuBZaGV0FTFiNADJ/wDSWdnRC8MVpNK1ze9sxA1tpZJFZy5JbbP3dnzmO7kaHvVqKI8+0
kwoYsyyEnQjfCHMMGUMdLWbPYJMLAoJfqbpds3NVWaSGYeCE1jd7iGp+f+zalZe+EZeMlGjPpYsv
2Q+OzgMSrGqOeinlaroKDTTHU/DV2PrE2PqFg1I/N/2vuAubEuavpCSzeMkaWigOpAVUSvLKgFTI
cGJiLkPIU5BBHrPoydK8mCjrUeJKP0McDKuj9BmGCLr4/PfEFUkvOWIZUamhwrkHIvWz1DP425tm
6fXKLnYp++7npj5Zqd4GksQbmAonLV/O0bsdQgKscV/3Jhc3JG31RUI9pvyBISoQaj8x5qdfIbNG
aMBqFybTVCKYoRbs4MJ46L7agIWrlgH2HBSAmAMyaVc8be44ljgTUZaLDokoz9inwYPdF8HU917B
ECQQ4F7bO4DVSxptjf/6Duv1q70sPDfVfVvn7KGw1wuA7BBjoQMT4uj/pHmN1OzgjCcPlZCgYg3i
zZP2kklDZvV6L65jfUURYmPpr6xTl3J3qGVV9P/w/kms4Fl9CW6uTq7PBrLHFtc5NUoO9ClR38ib
NxdN2J3OB5RrmaYOv8VkhORz75CvuZXXANdZVP1B3UodjwAgR31S3zgl9KIcF2rBAcNhEINZmh50
OxGdeWE+AgnfmB6zCbgPZbDHvqvC3nk3V/21StaVGVg6EC8K1eJcxqdsiasWHr0a93evmfc1s9Aw
NPB/ngWR5Lr38hNa+IyfH5ptutFhpO6apgeHSGDwYW8CbbrzRSG9sMOlwtCQOYxVvIN/0GWgjwR4
cWjPwD2dTNfgOYafKLSw8eZmWeLnbZ3gkVTP9XZTGKQDgcYeJigk6rqVQE5N7Ug4OsNHhwBobTv/
7ChfjTTvVuseHhMf4eEDAqfRh0raAtKklsP+7VWvL+CnUwuO109aWouAwvQznFLEIPQPSFWERhl0
yj8YE4e3vgihC2PgmSHoH3mwvmcy4PVObztu4g+hDA+rSOki/VHLoCoYNyJuqWoPFOfl1ZZiQx/0
yZYrqvzagFJ6f+OG+8poGIBFR4/bf+2ijbqKHBZpYJ5mTT0Toqf3O1ZYQvHm2wyz5ZZgFPlIi6M2
B8IrQNLpKIeEIQArNpY4t2Do31UUYTNdh9B6r0VkdtqmBXIIvalL60zqpyDdVo8ufF9c7OAc7fOd
D8wTI4U9NoPnHqROHeUPNx+bZeTm5T59asHOp38+4vLzgI0rjDgpYrdAwzwlroyZ5iMp3b0iqC5U
7A/p65U5fDe7P9cnQU5aJb4RlCabVWRqeKZ8z2RBg2Sh1KzuNzIEVQr3Jq0iiouzzA2qDE/Ipaq2
Gz6av9eayb8KD0LqgnyTsUYV81wVZUOYa9VrtzB8/9MNWi7fcaKhVhqUg5AXLf/RMIUMYdmqM8HF
Z1GHAi27fS4KBvqeTJlIpi7i+nWxP2dS3j7BWzlI43GegR0msCBZhtUlK11sS88lW4vHIGqFZA7Y
GkPWel4OUTuGSs8+oXTBn96U9y3+CCKW273E+jgeiq2GdF+BvAmWPXETdkFTpBrCe7whjld9wX7J
HY62niDdcwRwBgsEAu8N7NHhp5rwkg+qg610nVwm5q1+7FWHN9lhB0k06IxSb0+RiFkegyYyN6Fk
6ztdaw3q8wbDpjBu7TpgXuSgJnS6+owthKyp2LMWfwLxAGtgQk9x0trL9uTHqdkXjmQCCbUduwHh
iATGKNugDFpzUsVSiRbJoM/YFHl/1anQPLS9YkdwkkL+vH3Wv/INbbIzGxwvwrQS3hWKHfKiGbGz
ToGjgDgOi0s6s/cbVjBRJwUt0eRRY+8MhJwJXKqAontk/0wTQ6PNh7EWA3+bJOo7HSW9fz+yFaOX
Rrx+6NvwUOL94z0G6uxi57g18CmL48Fz9fni7dVfpPbXfXXDfBEBaEdViJ48P9F/gZuj1EFk9uay
NhuF0W7ShH+j8YlWWwzUvo/JLhOBrFVvi+gancvloDFU7ztsMzetnFRZvJyfFZeQJdMQjXDTt8fB
41dgZX46F7bqY50FVZuuVhljpJ2ZFLgmQb3GuiwyDdT0JFDH0ApBoHYMmtv7i4CHl2BkQMguFkKN
cA1pQ6V0B22npNePJJQCxpPBUYpqimCyf3ppD7jq2KYSsi3UoApV1eI8ozawBEXgKIVQlLBY6vHP
5YfT0cYhwnUhN8FaFluHzxqJyI+NzI0nuaQA8myPQxSb2TcF659TbL8o07SgEZ0ORGH8Z3SAkxoy
kRLWx0JOv89rP7Wu37hVr1Z1fO9TF2uDhy67IVfQMv4vl+6M+qoAu3eymLM/eY9dqIRa0zHtrQa1
83i3obiZVkCshtCQ+nSMtpMhjLSKngwZ4D6LeLQHCF+MffUGOxhPkCQ1f5MH2rJt7PcXYiJL4v98
xmUhFBhxQns2FJ2rExdRypMNMOv8v2/go8y6L6SJeiFGavCX7uSaTIJvNgJSEE6fF5neczcHL456
bXMpndoONh05sfrZTISDECP02v1bkuFLr1+Ogw03y9HjgSVBgi+dIVrYpbEujMunAlD8+Hj5BtsC
z75Vj8YzdPJjmGp+NQEfhKIbey+WkEBq2kR5cPeDZKhlBNm+znjZ0wXEODA8tGxg1geXjvbwi8xI
X5Zkob2ycjzWHMMmTESPa/rTarxlS8cjHxoKEgiaY6kzJeiRuN1z+4zL7OZ7xAeaoPImVsWWC6yv
8l5K0FuUO4iGeiMbf/ToOcGwxu5kMlYUZpdGeOHDT58KHy6WeOqiiEnF21nEGu4URngFpGo78OVE
2usHgq1n9I21YKh5Ep+dCQXwAMJuN5S5sGbuDXAJvTNR6HsBZ96hKx/lWrwmtc0upA4nbvTDN/Pk
AvzRGON4tb01suQOhrIuNS+oeIKRmkJhk4yNxFiFSwLbEtqpjIIlHq9uafbVkNML+hqB4gtLJuqv
N1RycnIseqKgBs53SCokmwB5allsAMdnN6o0mw3mxuNiLI555J9qtRbo9rZnObsUSFAhuCEj3xLp
aU2wmc7TO285nmovTkbCUsBYWerc3B2c9voZFuxXGakjOuDB3TCVJAj+fL1wgFXs21wsmeqwbdkp
tUXgNPHTVZiBSSPWBHqCsJP1oUNUMibYtsp4ERwk+mYqGbf0S4hNXyJCPMl+l/M9DJEIMPlF4f1A
sWCztQdZLJ/ytV2UqfR0O428bmUNGSrgFWK675vS9+aC05zDKtDmRkcXxtVJUUYsXdAPnCUTFPtX
k2w9wBbudU3lTtZ2EHO8pNZYbMoKAVZT7O7I2xuH0LEL/Ee4dZIvr7V/holQa58hNcNFofadaanC
fzBYWUQipP5VAtxf22gmOrNyqshpjCYGFqhT9ZTa2tGLxj956UCBCLGq+rUZ9aD/5kcyRZqt0MKv
MyIowYwWlK0L7Yq1ythnRLz2DXvxBHANJiyDaqID1YZezn057cgdcVcu56/bSaJ18vSzvWWw8vzf
OotvHsdddkaIGSXP0Bzy992P4EdGy8nHCWwUkYM2+Vi64A+ZR+mZ/3w8OgODutTfRJAVhz1Ay4Fr
tjvb5XV1reRnkbpvSTCj2hExyyLusk7RWHzxlAhn5/kAmCmk4KDeyHwni7pjG9oMuyP3QVf9+Ik0
IN5rwcDqV0mVk1+QWqPTMy/BDmq7IOiFjKAxX4kA93boK9GOugjla5Dd+w5h5AxYvbh9gIAhR5ef
IeO7u/pTO0dq4q8pYPjg/yG/w/LbME3h02tnt0cWNPDOuThEk3s9thwew21Q0AjTYyPfIQoTQTrY
sOu+HCgKTdPBMdn5Hj+S09P4u5AnT01GIi5mYajFzhmDsRjtBn+3i+revb9rHOSvEgNQGgj7phrp
1XlUn6wqZNwgPBxZHlPQ59elFBwG2ipKSQ/F5NsM8K970t0K6iIO/zfiwD7ensrnR6YRqPXzj+LZ
jKtYFxj6SQRHExOM5hi8hFGAJ7v0+xmgYoZ1lxIN4ebYJeoVKVe5Yu+Q+o8ZsKFbjkdK5BgmZXEJ
jZ/PZrcXcsClFwM6+J3yzdMXUDNxs4Xa3BWaAjhtxT9xP/zrZKKkqdhQF/YbuEGSW5kCUwWrz81b
U9PSbVGyuzqwtyKEQTebq24n2ZAm1wJtAg28p4NGWU9biZXQ2fAYUx1HflvFHvZE01UfwOzblQcr
SN0KeXl7uX607OMplqTSKu/oO+iv8lQ4+b/HreB36rztQx5C0lA6k9QYtkJu/NAa3cUy8QPtlTBh
AOjTMc7xkz9C6OzSTwUOozSb7Cg3H7L1d4o6p77L7EbGjLEc3S1Ml2pr5kkSHlnpaoHyc7OkvjTc
FtU36LhzSwblH1FjN+K0vo0ZIOscwGF2KyuqrMKzWld6PdDfHyuDoZp+x0H5snFwj1QZPqDrkHhZ
gp6ilG8/IsrYpJQ6nEuKSVsDIMPuErop44mcJcrNu7+V0g+AZXETdjzIyNWM8Xt3Kb2LuFd+3FuK
VZ+HC717J9zh6t0KCSOngTQaYz8aFabO/XDW0owM7VQHgJV2waFO7bgQW1XytjDLNRzg6kZ6Go6E
8SzBFsuJgNd4zfQrhrBgBXhOkKSglYojQ1FhTIIlFIcTmMVwv38Blx/0AhfQ/4ZTLfEXfBUrgjDa
DTBvgvZL6j+P59ZaVVuEh/sjRQ+zRexvKoswyfYTGeFJTUWoN88du/ffW1cOJLPtTmXaVEa4hZ6t
CBb+SBt4f8dYNbTRnAJv6HQ9NAY5QN9Wjgp9MM2jIV0OUx2O2cuINod1CJuTOMgu1Zpk/yscGBE1
tOsrm8Uv078KIaOqhGWhbH7jq4Dk+ua0ySEpkEzhMqNhBsj1ypIIbukUtjyAIXg/eYnTBI/jkVBd
XYTDdoxsFUhpwPqqhWLy8KQtpVdMsbylF1Rw1kPPsh+QqkBWWLPYcVMYWfH19VCLk17+PWpnds3k
aZhd3cQfUSq3MK1cnCHOehoRw5WaSwgqByrwt2VEa06VI5RvLHs1t1b5rTyV3+WjbDTrbEzqfjpT
sGp6GzGzIPEnbtqG2yYsd1E+2lJfYWl5lG3+3o3ZFtmVo6YzhjDyBgeFsb5fgyE65q8RWf4rwVaY
yPmOYtUdTIoXTYxGHcVqnEaczswOvj462FdMpuqKbdSdw7qTpgNCBNL1X2P/qZrGSZ0BSbl7HyBa
ji3zNsevt5CfqalX6Ue7WqrKqT72coxVn3HbjCy37yAVrakNbDnbsZDR9NvoMpc7vHnZeZ/NZPwm
JonkbxZow10zyQJkGgvEqDeUcU3loAtG7sSlaxxIfCWCzpa+0NhW6DOyrNzIF7XcMxxOayTdniMh
wT7loIL4CIEYrLa20ClRjNqY74iV0clEnoSnssiJ+nnB+gJUaN33+cTuNMmAaxm8L3tByzThSaBl
TaOQJJqxrjAqXTevRombJ3ACKxwJ4QcpeIwDWZLSXixp9mG2kjZmkeNKxdDrrsf3WfoxkP5suFr/
eiTp8bEknt7pa4nz3HIjYgifTUaOeqasYki/43vsx+Qlb7f0DvSp2FcAtogJYjxV7nyOteZGxBur
hGCGyhvSoq24lbZpnDihOjCs0AYz0WjIJ82x//ZpTtVJUIV/WyT0weaj70pa32RZ1gEQVC/56SKA
gkpDKHAd4ZUyel6guwuSsd9m7Mp8amvgOgUl/A/xtPbIDN4h8Db+6+VXGJ6JtjyPzTR+rmf8hRnz
RDdOc7p/SZQaheC3soTMczhkNnijwvuBcrF0ttNpuh30RG72nu2fXahgh6hf7hlfFo9hEQc8bhNj
oQVAvulkVBI1wic0twKZZd9W7YvKsbsXSmuvigZyMv+Jg/nRf2xttMgAItmQqgruXSB+pT8jUpbM
gfs3sLZofeFvaXTZB6mzIBHk7oym22M0A6+VP2mqZgTZka6eFmLESm1KhD4BA/og2rd9OpsA0czw
dBWmTJMLDT7nmeUzDQ2zjoPB1/dcWbbakg/XKg/sAIRF43EYBclJ6W1aJtjNlLzhsaZ2BpDGRMtU
VOm0xepShDg58yhZQfp3hbKbFXNom0ml6adQ2qcicBOowmQYNs4e8pPJEHQrKOk90Z9+ULn3+sgG
WXB1jT6JFz+ocN3fSCq9jC7oBGR7NcEzMp0+NPagWjUgg7MUvFJVfYriC27OB8h+XkswJoSVyDnn
XcjLbb3hbzHtf1HL3dds2zekWK/GFOYKEzaEXVw2PbkxO/eS8zyY/Jbyxgg1DIjviYmyfdyeB5Yw
6H62QAFzdmQvIKe+gL67dwacPJcEiRo4/OWaNNXYVwswOVBNw0wNLLwYbeNF3LQBL0z6ECsTYB2z
MglPmizBMyhLqUVipUBCwbMrsjybfSFDLplIwKEMU2Gvy7YCYXU5cVSOAwC52TCWAHuikJavpzAA
jNGRPTIKViCVd4A7HCb21vQ+GUNqKZ07X8dC3HJO3nNL98YZLku2I95S088nP06TsNV8cxzbdCv/
JCx3z+Ps1OYd4X0wJJBgFDR5fucQGn6/MiR3IfjBdiuVdBC9KEoTHDaEVFAQgIjb+xluuPoPhJ00
GWDe8cJGCTHXZONqqXAqIZkF2WJ/7rp/VnHQwY5O4xvpL/2MPbhaPKgDHW22nGM6BCqHMv7+jffV
k2xWhU7j42juPA6i5Q30ae+G3wTF/HXHd78SNw4h/sjwExaQcQVFQw5bU2xvzxOBxgU2gIVEG1Fg
/e4Ub4upkcJen1jEyi+B6Oh8xcNFF6qt6JfxAdmMaa+/AJs1ruNdhEf4q4O1MpP5Pjlxv2cCmIw5
Mt7VGts9ZIlawlTZG6z+FyFoSFcl0l+x1uHbBa7ZXgSld4FO7l5A1Fbpbs+kM/qDBNvF++QlLBNZ
3UipsHitV/GRL7HJOr1CQyYBYDxRyoCzGnlc6cxl8SXB/qW3jWkipKNzEKjmJtYI3Jsv5t3f88RV
HzTLQlxS7H6my6k2wMYF/k+4K8P42FS3vGZx+9shN8ULck9QP2aFt4NEuUDYDsNnyg4Qdh6HBahK
5eSoiR1U90IKs90OqNAUO/tjlz6504v25gsx9lkU2RBI1VseMpH6nqqvirDg4lqwMlWg8FFDm7wq
gj3aCSYGJd26Mx7qp4/3wtD8FH/qyyszbdzCnom9as8yiYwaplgyT5JUGxVnzIq6e0iWklKA9zFT
lS5qa7SVPqEz0YGlXyLr9ga3F63loRtup+66JW9jjw3Egi4fWKRVqcXB3exbnXy3+I0LUXupgyPe
DTg7du8f+31N7LGTA5vxUYL4ZWjZVCAAb/dkVwcF+ZNkAgZm12s2cv2Ov49xSXgC1z+x9dVHTZsi
KxpLPAjOObmFYeZlFhtnh+UGYw7GO/KsLVa7UKdaQFwmhl0cNHEYhnS5fpfohfCctujmnLIvV7ii
VMKg+EV2GRdJrjHdjAA6VX7pSQ4zOarGj4GqERMstksL+ruludt6KrR1YVdY1cv3tZqwIBIr4jhO
1KZjoEILVtLoP1YcI3Vx1d8Irv7c2FwhbU8GMwOb7+JLjJjIFyVbEkXf+tvYKQXCdPAFtB91ZfPU
SiSdOS7OZeaLaUqESrvx/RYCSbLZ5dmi3OlEiww6CBvtFwV07+++M7TecMOukDRZ4qkcB/mqWj22
0OwtxdRos/i63h7E2lSZk4flU9WjHzs89/c1ZyLU/sSyj8o7WwLR4X/8wRknTTCzRdApTIJW0jT9
rxm/AuW2vqxJ7qrmt4lX1uw7pKmY6W1aRDqf6rG6V2DRZM3GzN6T01DvUl0yH8U9Bi/Y6xWOdH+W
L7wEGIs9E9qNFC8ZwtK5po5V+isiDyDNC+8vQXREM4v/uYFtqVlQMW92m7eeuYMDz8VRm5T7jzN2
0fHguISgSTykAtyG4V9B3ccdbRDr64WfKfNdAK5c8z3X1Y25kFTc3BdvBokt3gUrmvk5/wMcDe7k
k372ROwpGt2xJd6fPwEwksq9KU22KPgsjR2YfI5XGbNQNZM4Mud1S4TsX+emEVPJMpnHB/owrhPe
5Two4tk7HFoV47NLMxhdk00UZc6XiyEAsnD74ZUSEhqmnkDv057t8ofBDlOnvFDwZAU1fbcUvnhm
earXShGkeq+L/6irSc12EVfvtPy0a4y4Q3ZmTDTUQIL7uUUgOYNJ5L+bZlfddBzq0WfwQmzIAxaa
ym24d2NU31YDcuQgEtgx5jGNe08qv+XyeWnw7l5i0SWczubyd+QaP+oMpHX2GzUrsW5g6h+gaq0k
3YdO4nOP8ccrBDwwl/nrXr8xI4jIE7P+X/V16K0cCAtrvuWFLwvMzHcSN9smCKSLZCY0jfA7ACdQ
MvIb+N+a+1Olb/QRap2fikUzIIyidhlSPY6yLlyXkqIHA8M8IR5/FVkrbI9hjFvpETaXWdYI73bF
vVLgU98l+Ow/4msdfGYzhb4CKdxVFP0hqFY92CDkV/hSr7Wp37hmqOH3yNpf4ZzKesz7HyFgza8Q
IRmfOmZ9V8fTes1p5jdhqvOiW6nY9ddZiUhakGO2yLerCSqNLp09wGVJMiebQpgO9gD4iuK3Kkth
rrNFzdIFJqgy59FCiwSwE75HjNpzqGVSYCw6d1f2fNNDkBSN8mM4MkgoAN96uBwOKwiafphPsQXb
1UlvsreL0UksGMz3LVmaQnas8XQeCbEnC99ahnYs60iMkjwXSdb4ONNMvB0JdOWoYYC3zhzbM9sQ
C64ZrijJ3S1xJP8d0UyXxteiQ9mCvHrOExQ/FVigfj5pWgiVKXfN6oCX5M5ocT4jL4Mh7Ru82dZX
Zs71Y6jcTCpYjj/zuXEgO5HIFkdSPPOG9xzwTi5cZCNpqVMCUH7YTXVsdtVZuXBYM1GLpduWsAcq
ljz5bVtwx2dRufR6lWxbmL7xJ3y4asfPw4I3OtT0gMbNGZw2o2kQx4oo2BHNLhvse6bn7xjnBihc
w5ON9Ke17Ncc8ft1Eek3EIKRwK55kadqrkvRh5XpALU8JhrBSxMqJQX85O4OcCfxryJfrCBvJO+6
vCLBgs/Ew3Zm2lwBpsVitLc+7aj7us0Z3/bSUsk/H8JogjIc0ZhzOLgOkNntXGdVJ1hAKpIzcwqt
tz9Je710/jZhhSlxk6WSRU7s/eNKdbqn1VKfbqM2Gd4bQZtDVbmRTFoAX25TyRMOOpmS31A8tCkf
9pEs4LIbt6Ok0Qud3OeJKXXR42gQHV5kwKY3ScSYRg7wesgc72MR0kMtNIZy1Y+e7WTVI13Q+ZqH
zBd1cH2/e7em8VCvIracTnrYT/3s1gOMZH23OwN9/NTfLnYt900TsB3N0hqRhCqo3LIxtr4NXX5V
Y42xvTpAPdsPT+FjtbrmMsr9vn0BvEZEVrzAnUi4tTjUYgQ3AzKyJ6KOfhLCazZTm0HFdiL32u/i
GkaO3Yly37rPi0+sBfD5JHIkq7KtP7TzT6RbP2MQvsYH4JXL3uF26077b6BS7CVE7CQ2+WvYR2DM
BW0iNGds4LBXTOn3tP5zcpJNlsI5UcNqEpOcPgWUbbCaVAPQ1kdz1zQBVAOw9dYFxnz4q3twcTa3
/oAuShFx2VtEB7j0/dMs6m76XpoFcB2S0ANodq0iQZIOw+lwr8+wmZRDq8NHV/Mu0EN2bwU1Mgaa
OuFG/ovOYjFtxCVV0s4MdhzSsEAtti93bIdxobPZB3UK4nTgpE+EONErFfubtwtUIkBAa5tYeJKJ
PDPdUMj4KgoNTlvom3K86UAAj3TVaNVH35MiMFOOnahhBPmWI2IPB9lnpKVgTLXSbfHl6tp6ihbQ
eBRHIl+GbNfB1TOmI/k1T8h+quYmSRqNOlxIx9KCkhFJSMF3vWhS9tC+4NoqcjXpazXcFzW47sty
bcZ83ct7rUxThourf+9daq0Et+XW7kKX7uNf68OGlFljseszzu0uIPysFQGlJCcbnFKRoiB+rU54
YsxXNGEGJIipopqbmWJGw4oiOABcl7sv82T3ezMoha7fmZenDPSs4SM8jnLA6VOtOGokbeIi/VEY
P+vNQ/rX2We03l9BRdeSXc+xeBc0P5eumSqwOgj7Jh8FRsdEphcq++JxlMoVjemU0BfnPeBobPd6
Ybia93NOih0Ja9T3LXI992As+abE3rB9n2KTqRC8uQNiX9j9dSqNXEw1gYoLMm7tTyDUiTj+q14q
bkzWvgCuSTELg1R/peCXW8ZgZY1e8cZf05d7Kyoieh5ZkVPnk88u7rrJ5XfBTBDiFQyDdal8iFLr
8NfaEVyoeEAOn/UT1Q7qHFfp/C7GvleMdCz5MllpDZDmM5GRaorjPXM5DOgol+JVnr1FGgWfLzQp
G+6ckYypy5tHD4AQhh3HNduUV+REbDWchIq/K587dHg0oUkO7nMZEP5PZe5wwhSp8uV0nIwM3iEP
Jl9o5wp8TjlOPk9OXOjHswRZXdj+n70wHnnwDK5yGHZkLX9yC3vi/mPat37q11rXAmaqzzmk/MSS
IaPSr7nEdbFc4nwjLQRvy5JFgvExZsO+KxzO0J9eGtiVH20/StzIg0ZDxRMVXJCxt7YT6MFX1Z8t
2rSLBrEHto3R9g9E8vCbTKwGZDG/Aa0XI+5Rdy4QteFbbdPGHLC72I1lwDy2jXRRejivb7LmOJPA
YApQS1te3k30x7VwE5TD1Y0JATNXeFPlKZZqeFm8b7laxCOWlD/v+B0AsADqqVs3b1w6I6ZLvUAD
WbrRyS7/xpA9zK0zGmf8xjgq1nDKI851FcGHyjgy2cUpjXC+k17kJCixQqPcHusllVg98kSONC/M
mFHQY+BQLiclLlU35f7ZvrNCvPPfT3bO4ljg9hummEka/0aJDL6GefLgL+LnOvv35oQlrh96oYu+
CsYo8PbtiMVx0L/M7gk34kkkpz4N/kC/TxGzKze5QhELZFIv84zo8ahCkcbm+ctJpzMNXZ6BNu3J
m4JrPVNXaw8Wgt7pLSSjagAHrv7p4ttHI6V2s2YpjZ884YX7vRZMdMNfPhNP9JP9I/ExgEEC1Dhp
uxh4CMQZKMkLzfpsNQOSUTviW5xizpIklF35gVfmOUlZ5OVBIV9ERLadNCYcx2kMzjqNLZLVNv1X
1s+/J3fzTGMAOG8nfyKoepR8Kjep1qSfuWPFBDWZfQuig9i1HO2YN3ce4o9Y0KmFGLQHOeCT/3o4
e5H8cp9A+p+XXOGgSBXQctP/5jE/j4zTl2qeKfjN/DFovLQtNLTYuxXhlgxl+ruSGfcthTe95OX2
6Z5rr9ZSz9zlVXvh4qOBHZm2rHdfWPiuVlBnth7tl5YKSI2pq/eizy+3qfjGTjp0Wrh1BdLW7Pf2
fFEQIQ3N7auCOiv9CLJoaTFUzS/6H4q/GQ0pBB6NIMoAUezQ+2cvwwP/QvshcPYXUq2PLR6RIYe7
ioTcB5LMm+JSRzzqOMIeIgD7LT4DE4auTjngJQlNwVPDBwmvLpACkNHFKRdBlRyZriBWN0gyfF+J
aMJwA5G5o+bnf7Vfzb5S4J3ISZ0euboIySxowE+1GObQR98tGsuQyQeVPYeaaBzpk+6/rNWhuaba
YZQpdFkelIxYPDoXnNQt15N7TO4Ipj0m6HBT06upRlp4cU0AbZrCTpj2n+Kk6I1IQrkTXkomo7Yo
3wxDADJqznK1n0l9TCrmIGWGGgb6PFFFhhIdPcUL1dwaaQlescaq9S0i8wLBsTcOplG0OLC4j+lS
jvTZxOHoDK31k0MrntBNszhFBmLo55S85OgKBUv+9MvBVmzaTPhFt8Go8eIg529PFkVTU2RV18+Q
dQvUcQDtHPEWOz4Aoocba/jeW/xAJ0Gzwwnn1TIhtYynaEGC2MrvZTO+fW9xgWgJpKo6SkRNHOjl
AoQKLONUBSAWGOW+MxTImsmnzE7St/nvGdL9efXhVEP38H/t7a3s3JG6qJbxFDBC742wNMo0eFkL
9o9Vi+mZw6++Hipsb248DX1sCyLvo7jyO8gG9XiB/WmakBmp21hVNgGJiEgzqm7mnv+1GTQXvkf8
pWwyAONUcONo0/Zr6gg2RkC/Hmuig/ijpnmB1GwhwQ2xlSOB7GPNmtyTsJQ7UiJrfzMSWNYL2sma
XJfd1HGlrlnVaNM0vdlO0ebSgPXMD1kzXmlQs853/yV/wdFCdsC+KTVhaSTjJiemheu7B/djgIHb
lCzWRhTQv9rZXZZ0XklobOoiE4HWVEQfJ0niDXV5wDIHKWAd4ZTStshlJrD05YgJc9aJIBq5QyKN
bpP/0m9I70i4Xmzbu9ImUPGoVOxVvVWlScqBRS7XgDJYYH4vKtaRKp49oJpFghkO57H5VlFl0g8T
YiyCe6QJDBAE6WMFWH84FvRyOqpYRgYtF0GPI9ZiaYYygQzOZp7EG+t6JDMiKKiaOy67E6ZuiNux
336XmxeZiDcnaCbLv54jf6YkfBvmEr+5ePEUv56hNrx5K/4VUlSYuVvdUI8knI8k5qPRVlXXFAm/
ncbSMAFug6VlFpXsYUtGUUVYwa7migiioNc14pPevcK12iEtY6BovQK1i2sKM7XKg9hWXDIZ5Ouk
zdX4FYQa/V0SlTcCNvrMfFS1kpifLzJcQ9CGsNYlkHKItR9okpBw2XAXFdn3/i9lB+e9aE5HbeEj
jR2Cp40lF8QR6EipnWre1fIMmwgYlu6VtET/XODvzkmrlCKVVCnIgNFmPULl2VTvyNq6x52m/M6G
G5cl/vB5/RDqMDW7GocQrWytNUZoK0x0vauaGafgzhkRR3SWdnaobJqK1xvYoLBTgfQGfZQmkxTX
rn4fDCZ9ii860ok3Pws/uPvi6CA1kFc1IhKCvUbln2D5aqHgaAfjjSZbbSrf9OT0D+OfFcL+TRK/
cOG7gc+xbU5Vrc6x6Qx7B0JHEsYr9h1MRliYirvnFPgIrQkwZ9gI5Ci7cL6VFNKSEumr3JhCQUqm
mMZpg2BMT0XIcgWPDVXwyDfXFk3kQgQ2Ojsg6ZCjHQH0QtEgmFqLEraRnENrBmZzsyamJ7i6xFTp
O4AyxIMCi+4AITC1ORdhW8shG1ek/IqGvqpdfRZgcuKv2VoL40ry+3Ai3o08gcDxIcVIbZWKl1uV
NuqXiYkdzAQeQqPrR1ybulEFM3Uyh1eJwALU8qSpo0/5Gfw209FuKBHxbajGGH/7yQZlnEJ+nKr7
MtkUgEr9/YVRCe+mSOYZhE7qwPdG2ib4J+8EPwPRfG3TvwTJoGKNzAcRIZyZslZ9gyzbz5bLWvDO
UYlI6SgFCRSXCFPnT4MKZmH6Govx1/2YsRH2iQrBSV8wpjDCD5ScFumqiAooUNQXTGcQ9kDqk9r2
+wVrnm4JsC2E5WL+IXxjNj/eFZd2Pn94ujLx99yLRDRWH/ykikud5xxX0H0Wafav6NIdJMctHGuF
ePGBcW6j+KaFibhDCEwlV9nr5iHkSwLeY2SWo7Orowl2PfpOQxwcH4b9dS6JyN4CxwJxYvZA7AuH
SBpEjhb+uw4V2TtZ/TYHw5KBGQkbaRu+DMDm9Z8jxrVsFjV4NfDMygvbaFYInRd/I9By6JFbIgmg
p2aJ9QtnIumX74Qv+/Du65V4kDNOYDTLvpFqa4fye+qzAt0ib5OCyuHaTl9QS6D4VBsFTcY9o3Zx
qmhyiIPusg4Y+IZE5sSAlik3oEp9dlkln8qD+zXeTvz6n2BGKZlknwcr1v4rDfCvQj8jDkrxR3Wz
zVu05oCatpi3sTXznIz0cIAlKT/oR/YRLLM9zVkwzZ2iBK5yloowzpKSLfsQD9z1wH6lE00DeOpz
SYSRhwHcUsnA8+sue3XPZTYbgZbH8G2JAtX5xDabTBIy7W1xv0GKS7xGDaTa4rB5Mhw1s2Vt8Qqi
TPvyhADswdC5nMh24RAeQzOOFfKp39CdiQN5ELLlX8KPR/Zp6Xkbx0+T+dCy54+TuNbleDKbGISV
5eMLU4W2KW36in8XL5yKGq7+xBPGmw01M3dQqQNZo75hcBgXpzuXFzjtcOHjmG9Nih2QGhbxlEw9
RAl3JucRE9qpK/5t8bihNLpxaGh6NzZCgR70MLN4D4+mSwThu1ncTLck+ncm9E4pOJgP7k6JotGh
lFbfsLFWuZOeXlCCQarUs3aZSF7rfY7ABlJIrPArj5YdBoEk8ISFnAUwR2Y0+yV4HVZEcMhsfkjC
u4G7SfwFaeeUsPcQfDBZ4RLOfAa+7e4bp2hHlv848ooAoK3/Y6hjUUPiK5sBYcCmkhP5zV1SOFQi
g47lpLWyPs7QocS8zKfImGda9prHKOrUhyfPwbBClLOME9A44brrEv41O579yDZJCpHHk87n8vKW
hIVAI7jrSXzNzgZ5gKoOPBzCTMpm0gM+28mFCSa9dMxbRkLOdxDKyY15pOJwD+IqvfPhYbhbWofz
mSYU/hgbaDPcXfCs8Rfhh0YfQkqyUc+C+DJzZfh81CPFyL977s9lt+J9iuipQ/Xb7Ipepjy9oyBs
0q2g4EIZkIZh+EFRDxMXG1gP5T8zQtKTykJt64bYaEpWjgaqc8/ziI2p2TWDIoeFpusbWoMIeKr3
/7WkJ80vhXrz4VSx2mir161pPxiC45KJu+UZOz6QktbTF02ECRai1CKBmeVP6t3kOvjekahMsfl2
RPXIiJn4j3iMDYCXP0bzovORXkRElgSf//G3sFCdKMhJ2oCUuRtopH2eAezm3lwkZHkVtlJ7DffP
vgqqg9p5YmPO9Npv+M/Jly+zGiXfnUADHQWgdDIR/LsrtNn3v37BpFx5WjvAo8X7vVNNClwBvZ4D
p1nFKF4QAPCMnf6kem5bHSIsE45dbUgoMjsVNmGRtS1BcsL96mP4jjsleXSi7pZu1+lMU+f+021B
07WxWxJPucvQxXMCEsS2LsfPLVP0jTAv5xvl0+jrpGLKAyVnbiDZ+qLxfBouGXBRMFdyp6OTt2yw
sILdLbbJiEv0my5buZ1QFOulFn1gITyecmv2f9m4dfDAjiqHeVk97oAA7dJiKYIIrr0ZSWVovZHJ
29v80HPYn3ys8pPweUZ+mDHEIyMfZXTMptisxuiBplBCTofJoEgUI+Bw+DI6AXoZ8rsR7Nlaqsev
XQX84DXESsLxGZBkbsYf02n6zXeh1A9x7JuX7/7+ucNNE/M19hmB9F+Jh56iH4ejXm7fiVxo0dQr
2Vba9iKi3p7mCGsM039tpcUk2tEvwM43gUCVZGje1H+iF7l1s7HLyqdJ8UdDG/gwDqMam/AhkJjG
Jp9LhsKf9wfahh5Ip+rggt4NcwpizYLgHBbRUcrBQRFkR6TvIYPTF5Ahv2lOfcLOTO5mU8ZneNk9
HcQIwipS9J0XHMWDdMwuAfMUk+UO6RCw+vPPry6uX3yvUcKd5IG6efTcxiC/GqW6xNFP/lqw0vQf
K3jcjssgtEQLVAhtBTdBynO7o7AwAp9hKXCNuosNMmUCzZpxNVBJVrdeM8Hk/yCMm7OD9Q+/0HRY
3V65acuIuv0uq2dLWmA4xUoM/eG+l3c9L8nW+H+0aH/ZO+mlmLTpIqrgQx2ZM9W5T7eWpjVozi2W
rf3GrAHScbbfDhbTTpTX+UT7V+jJay5ue1ukGKgH3tt2QnNO9RGGfAcNHBIV/QZPdD6dKgZuK5Q4
ko/Aqq/49rv8hMEP5jajfkuv12tDveE09HcPJdX5PhmZU1gI6yVIewq08+oATOH4V61lbvd2+dtZ
ORVjMtHscQ/dpul2lyKWjvZuxBgXOPKPBQWZ7dUltbiTnDvBb4VZfEEjVuomtUVLNj1/Jq7judvl
hhh0rHm6eNkBRP2mH6Gb2ZbnhSOo+01XF7pDJAEFc3bGOAAyvJP0R+7ygPL0AzuSTvLmoN3JwqP7
WCRjHOKU3drQLC7Ogi/YPQ+OXJkZvOnK7HriRhY3i/ZjH+vHQqWILOSrSHfmqX/No5ckhKsNKVfV
/B7n9apblrKcphukehECBi0SP2iCQan4WzXOPe6rH0efLe6Dm0xK0bVZrXelrNraHt9Ut+Gs9DhX
+WOfYJYijCaadsFYkYqvNqGdOC9YjqMFLeAVRxP2hsfi0reAIS9RTYJhE+l/ldSeOtm4fDTwHbuX
uTWJj3t/lapEBrhCXT6brEp4BaHY+Dagopcx5n7QBwzSW4QR2Ka/g485WHzVmoowRfSf+90NKNc0
7TgTt3jkHUuZHJFJK4Zq5Ylo1mU+mpNTolRJqm1E2W6TvXaVd+69ZlGeJEgL8AjExG9/8/3mSY10
cANIwRAK+g0TsfeuH7JgQMQlZQkzNKyxG6YEhr5JFOmmOtU0Q9xh33htaxV8FTHOmS6xQ3JJFUy8
asXRFhS+LRcWn11G6hTY3Rb4O61a09bZqeueZS+KD8/lwKHD9nEFHJcSb0Iw7YjZ9WKGziv88uge
PyunzuWnt5iBfs14F+S6QWk4sAktNX7hz0cb4bc6ci0P36U5tjqyOwv2zkBMtnb+RS76M9tCfUmT
7jzDCc4tFuasa9XNky5IwKs1oKZk6vzVYOamNXgxNdj22lll0IdwCwLZ7rHUkGSDwMXg/D2s5bXi
U+8o3pFcN+0Szor4sHVt2XO4mGkapm9yhC5IVDI6Jg9+r6yjagL1wgva2e0LZD8wSy4sq/CAs1aL
asWSDEPRT44zfM2LeXykfzG2Exmh2UnrowcKQ3rbg63S1AsefEu8XC+uu6EhylUN16qD7et+axD9
x7hINk9QOfk4hZguXLXWyIsTow8OsZdMUpbu9CTG7aoDxUU0vuLoxmgY05AHOlaVtwPCQavAgQpC
wBBznfrEXP+XJolEZ7u9lwDn8+7Ogloa6yREaEAUgTEriGn6c+wYkgrhxktAn+PgrhsUgAQMYWxw
MSUBWyV2m9sYPKLaUdWKAktIP3UuCrhherrYuRX+ctyB8uCL1uebF5fiRtjgilJWN+x+obXiuGHN
UXJ71LWPkViplwhngXTk6BmP45TH7Uzv7DFEMoI4NYrEAdAAQJgLWgknf8HqqaxMyjdW96EBvnco
eos+lMpd6fcrqzJZHI00Zom6HdL5l/3FA+h6TpoXMTkWHHa+l+M/K1kdzwElVngXZ0KZNW1xq4io
d0JclmrXSkSi+suhZ3CvAPIKsR90/BHR6vbHEY++reMOMg38ILCZcWlUMzunW3IhLAWJiLhsyxWJ
TTodqoLI1e/yBdZxwJlpEEufYe+G5MO3URBjIxtcAhMl49J2kkRjVRMzdTAO+2nkWymnmZsaPnM3
tVActiEyrEW9y78ZKGIZQzXeVNKhtTyt6PmcEtD3QDL0uXaoUExWBPyVI2vOL+JHB/vsSQKfFA4h
ADZpYx4GbQrm3gIB1mBWPR6/gy33DdW93Jiayi0A2PMfbQAEZYhsu76Ws+aiJO2Zotgt28tFXb+1
ObkdUb+MHX0MZPxxRewKNU4yY+c0YkubsiQ7n2eSmmvg36pL52eRemjsmL6JNWMN0VpLJUa4tsmd
i/hcJMdXOzjPg5CaTPLiSTCfGYHlWuxxOaWpctwDDUj0MhgZ6J6s5Uu0aPumAPG42eD5U7S9phfH
FXGMx1BIsC70hlC5xFgEcBknQeO+uJ7iNG1Y67XBsMvlUKt5zLqM4rbGoSdOrwoCf8M+5gjOEgy9
e8QtJlv6uXzKs55Kv6jQqJp3xGPiv3rwqlLThS/W7KRZAfgLVaQOLDptK7bZ1oO2Go7l26/t+IcE
vxYcNFkl41rpwuRS1EE3cFIhkPTVR9esTJmOIHlKiM7mDxP0DMnegRmr3+Pfru0H8hwRrL+RB+ia
SMfDXVG2V+Nvd5RbeMSCpBMDX57zqCv9U68M6ad9GKeHykWHa/XiMFgdIzYgGxsG7DkN/oMqQ5TQ
24kCpkxCmgW3t1t5DucMJz1kYkKmtwl0jaXMPJ536Rg1Lo7k8o9yOHv66RoyvJsiaGARWUFnR8ax
v+KB3boDzvFhTk91QtSpNV8xuT5QEGYeAR7U5g790Dtn8PvmKVH3PHvj+LuUzre7ZYqRfyymJStR
sPUlR1QFQU6HWAaRwZaTMXDj/WB2HFvhoITEozlA2b1ItZMGpqSGUAypBVmKW+fhnn+eomPjHOBb
hw2bXoUZ+oQXIusQqzcM/NhAbSkA8AC0cWj5V/F9IJJyuyCGyzkrRFsh0ZbgXo8NtEXQxjSwDn4w
OQ78lre0brLKb+kwbOngJ3qqUUCMCQZtTBwzabgwrhvmswT7Pt43yLw8UJ9alT/a3G79lEJSNuhF
ap1KFShnfOZsKP+1DVucsGXfCGBqvL/HVm5vlIGkhho4JJ1ecHdlhouylNqTd3zIWfJDZRUBn47s
IVsaE5XY7UHOUMGBeLhYmePIUaef53Cjo7+VC8tdV24FBkCQtKVXUAOwPO0qRhbxgIGqog620xRQ
/iJzIxmlktSNjwXntAsMqD3gR629In6ANe+q4A2XCuPeMqOROnlROsjyUoqvDKFFTtziJyCL7H9C
xkgfy4VGLGSF3YcJoUEqjEe0i+Kjdqaxfrtx+el7ffCFZiycOTSXaxQijAUlo7pg2XwHDKRtVc0e
Y+rGaHZ7d7sxE7atp6SKfip+TVB8+Rd+jBoYpxoXBxemOnOvr1fF8AJKdcD8SyyXz7K+bwhWDofH
OYcoxeqxEaF1IQniTpmeAR5WfIR3b6SkpZOnCImTw1J43rpmX2tDBnf3sglEB7TjhPWNxz3sSulm
mtI375cl71cjtmxtavTpHCJMlUjHkcyG+eycULy8txK9mSqvl2A1bB3OpOzSfTU8fd+Omgt/h13x
66jB7oto023at9xmknEee2DI6Yq6Ub/1q4o8CD3ueZFKTwUgqwB0wy1UKRAqjl2NjgEtAZRLlOo5
Dd/UfP5UJWA+6lm9IVsITdGqzyp8UuytKF07tt9NtksnXhaELHxLoTFY1DcwNfiMR50NmLyZD7GK
MS31AXBr8wFUEbSiRFAKO0WZ5yxp/EC9f6ZZhyk/tIEHQGgZzQ/brKA97kb2+9XxERgDUZezORqs
I74l3T022b0XrSR23MxDqPjPv8g1X1XY4D3fBud/BLDeeKX4wowMP4F5exDdGsl4Lv6PXsdRq7Xk
ckNabaGS3kn4AJ59jCwm0+faOWptCMb/pwukV8mzXPm9TsLxW6jXjAtrO74zwd5Z9putM1Sk+j8q
GJ4Nur5/yxz1HkqcXc8VgsV9eVoe/wB8Qt8npNIj5SmVPD8qJch0rvnFKxcoP6vCEILRkFNxwf75
TiMRedU/xovGXHgKhJScYRzY2cW8VR8Anz6lXfVwiViWZmNfgLTjzaFCIAMWsWomCQN5B6bCDi9I
o2ZM1FjEf/ZFf2PEFLIObp4vJyAyG/12l0pOR3Kq7sbdNfdXfSfIF3JYyCyujhfgO2UPKvB+fGhq
Emmt75r2ZM/jTh/cAxqNCOMgr/5ceCZ3XmGtNwaCoDGY3ZeExD0QrmtjTRKT4apOzgdjZ13f1OFm
Kq96bE5efzq34+dEXGGfNKOPz3sN1nZdWz/ceibn0G8lQBW3U6m6PMJB6TuJVUdzsvUSegXGfRu+
cTbdIjqSLORBtM+TVPnyNDdfumQ5OL6BgpTd5c+EzwYqMu+i0pzi2Oa0SKHfGnoqmtQuG2af0Cb7
wvo86h2fcAJLnOm4a7HHgyDSzzO4piT/TA27oaeQSpWwpGn1qfRiwAkvsfS+YYWOstYNKtZsd6/z
+OfIR9nlPkh5RbR4R5NMonmHy5JwmaXKKPQCRL5eKlEs7EwcQfZRCR0UxBPzvqvZNjIji71miinW
gy7lUIJOKdhS67f6BREvAHCPj/CJXEVPBvnRLejPbxHqhD7HDKOYa+qMfqRpdFLqOyeRyrxBNbCO
0zjXNUqi7HZpFgtjYM22pB2FtTuLGN5JVx0aHXrIE7EyPmbF7euUDYygGXxd2JrC9B0lF7mk5uFT
brCeTUTcviTtZtoLuLJ6oqPb8WtUVuPLwVmjnTyEe6d3fWOf+lxA2hdvJvjBgqOE+SuHF7+SH/D3
PZNLibUNLruo3ZkVpt94kb4M+2Qu8JCXKzLMEN8u6ZkIbjfeBvrPot8vV8QZtS6eQ8HgFGkPTWNq
7lis7xFzs8ov/L/nobjHjydZPIfQ9DeIshgZMjrNyBPpF3aj80r6xYGCCei4m868bHOQCfGbU2iH
ddkJH+Nak4jH4DZla6m7Z7RZ3Hr7Q3ApUmgwjeBH7dQW4lpXm6JakkG0dm0W1G9iHYJgXhR3iVzE
mwmaPwGXvxm7BGwxMY6WS/LnmGW52aiJtOaHOX2vt0otvJYNRR3JEvRyGmA3uICGZI/D0EKPA2L1
pZd5yplCGzZaSTSnXn+3QT++rdwncvLo3mibboFeX8ldPzJUzJG+CYF51xCBLx/2rKF59+ts/68g
COYcOBzWI/kqSta4qO3BhVgfjVt00oTQpQglbl84IoJHFVxh2EWeZ5LRFY6dlsB8kg6OyEHUJT36
F8whUvJ5RKnq1G0dWfSFDAEGkEkfT0iqaAzthYQPYmvfXT+1O6+eWgMtaJqZWbytwDSjaktY9lQu
/muSvQlIEGNU6GNlL6fJc/w9GGs783JVgWAFZTfR24AVTJp+vBkdGatwxBSTtDozzr9BODmSWy/6
UuA7tBt+JUQmNbGVK3m1Kx0OLJV1cPByTmS34mqliPpw+k7dJfsTLzv/QjgMa4N5zTkdVh9A1PGH
keYDp3Kdn2vjP06OZrkzhTps4Lr4Bs2ICH2Le9d9iIqr6ybAMbKgF0GxNYgk9fJUDArmkI8YQmcy
3qSZMBU9fDRYscKpLNmYnIvU1Fd4vBI2rxtJq96ekPTTZaPzeGBiSh7X9p6VR6B92OXYbHFGbC5M
q4UPsS5jg3i+V6fl7oV/kSuedTSlMYAXAE4hjBp3sttukbeq5dA/owI9+rwqbQ/esKUXIh12a8sr
kZTlxVO/24g5KfHEXi4COXVH3yo3F+T4rXoVLIe9iy1jlmj5SFlF3xrP/gS+g/QmWijIMyswTAwJ
fyzPxoNn7BQKs/Z6LNJpUZr9tKPMI0tJZQuerIGOq6Ugd92cRYv6kLdT8Udew6i8qseIPwQMnuWT
j7DDErwzjncGRPSiiMjt1snpjmHoqwx19smoAIAstuGcvYKHmOBS8htE5MDZaa3mTbIPUG/Drd4B
O2F4MOCUZ39mqmG1Aq6hB6LAEvL6S62Ej0QD0yWpQOcohhBW1S9tvT0V/4DJPkhgIWl4DwWSvc8D
jYZAbTMf3WHyD4WW8rheCxSAY6XIj6P5156a8sadgPzmVqPBV48gv+/OOFf/7LtQz4+5gXoesSml
aTE7J2Om6UUJZxsB+I/HFwejEkIeaIjzx/kA/wKVyEz90EQ9jVRFatpNabWRtIny3NDZRSVpOeQH
RIonh9UcgpFYJu9RZOsex9Toxa5O8cEUmJFc/59c5mpekVzaBxGD6f19ygHhqRPDvavhatiG2oMk
IEuB5kYAWxhvb08FpkZTnZjgkfq58aZ83zezz1FiEJiOZcb9jyC/PtPSpz0OyIpl6Aqp5qR0KpNw
PcXX4kPfaXwfxujvnsZtvwQ2vO0cHcjKtuLZJ+u0XE6p5bY3FOEG5JF9JTlc30b/SkrJTJRFyNOu
vk6b7TuZOZdckkax1LxVYRvZY2J2WxmDQthI2DI3BFXYNEoXDbvZt+1dBCHxT+Jy/7a/xk9vA7q2
cEZrh9S93IgO7WToBQz3vqpaeYErtcr6SHV6wePu+vhe1wo1MLf/rilRi7OxQw0RxSGo9HE/+tq0
HhyTJ0P5R7QgiVPPZ2RCQNSO0iNnV8FMthvdyOxt/o+rpmxnD9ZCWek1q9j1YPRD/W+yq0c7+0uu
pGBBpz9mOHNMwv8kRDNew1vq+uCuUg7nHGD6yTiofHsRZo71P0UpUYsWNbYDFxnaPW2Px5ITLvyt
iIEJ1tlh5XoD9pVRQhZTFajFAxa5XmvhITUJi0QXNpK2r8p8RMx2iWerKEdSr9H1gtUbZNEGn6gP
AWyKM2lMiB5FLNHD/ozuGXEOesgQo36hDmIJx34YIkRseY/Je9uqV7vPjqvj8QbmBC99u6x1nP+E
Ptb1R2oco4W/W6VJQH0dLJNTb8JbILqLRrcWEkgVhquJm306p9PdrH9d+i8DnvXrKoYOgMKA32xo
KRv3zrND0wX5fGhDA22igXwjEcUMvijRjYQXR9OZ7nWNMuMk0sUssWpwQavoFWrAW7+ZSXakSZ/3
Z+pmGfMJWW883APKG8hoo3DKx9N5wke6BFzOqi+B1+hohoOynUNNjw+4Th2yv5j47qpSw7Ule0uA
75TY+9E2W01z0PhvCZzKwbd57b7yjg8v/6iGPlYcA6d8APGxaiDD2uDpOZKi7zEugT0GgbVejVEB
SmBi7gb6uxnqrXXwDde6p1w/W94dmK5OV/wUswM338e+HNE8pGsrcp+2MioWza8vtSxVVfM3KyA7
CGHrIarmHJYL5TyEpwbXYOEh59sSbC5EyyKIXRXA5GXAU7HUP3ogver7z66/9HjcDOhJW2astOrX
FbMtuI+o6jadQ+/vqtNKfgv4WJeFncX5A/5WrbOgo2xxPHPeJREKBE7uqL0oG4ebg1OX3QfxzsdC
w88STxohBS2OWJeWRExt132TyFqfswk3NU5sE891A6WFYzAEoxeuk+3pcYZY21z/4Vqts7124AwQ
41lB+u+shdddm4sKvmQepQni0XO6Y0bAfPHqjh/oONFyiydG52IwEVyZYSvbFmcusLKPGjQlc6W5
9YqV62SXMal4cZQgbRw1WMsiGwBNAHZVoG5hPInhXOxvPCw0CFN6KnXrGayatWcwt0uF8Gd1USx9
YIBxzJB/x3Z8XxtACt/FLLd6DXfSJ3jKpq5xxTEc182kl9bt8NB9ttS2UY+TmbMqpv839j82Yrc2
9r2mMaMpo5YoBJ8mVS4qUdn9lOYQRfjcoC7YNBAsj3/pkJP+lYXpnL4FJPyft1mUiZKgoEE2U9gK
KSzVWMorXAI/Nr2k+X45pvAeLqj2+XdZjAo8E+0w5KlXZ2wgTreTJPybMwblJqvThlfSl1o7mXER
Jg+I1gSBf8WIO5YCxrGtUs8npemOmhdL/JIlKfdLtE2PmcxKS6P+7dXxxp+BtbstPAvJP7zGZisp
MNm2ut00wEYqBYpHvvx6jI+t1GqrWJJcVck29U+P0S1KQ1JRv9P5qG5T+IUnWlZGsV2rcCVdPZtL
YlV/M//BH32AIh/JOA/ODldKuFff1/lkiMp0GfhMqovfAjzcHTJlv57c3cIbXYXGyeovw8qHZn6y
yWI/3sImICTTURa2LZIm8rYamoQo3QPKGrZh1n1k/SKc4KXnWCRPOW+qA4SZke4QXZIf3IOh3/AV
VfHkHmnj22rpug50n84lp+PED6R9j1qSKcm3q/W1cyZudcZ31XFip1Y4ZcmqPUssvUrCwJ2Ji3jm
/TcOX89iKMwjkk1MXQsK81GwWBETcNkFwnD8QkEIKdYmU2yPQY8sHrQn28Yb9OwmzTA278ldxRnW
ejc/7ev+W7BU+zTI977iyLYWdy7euF8pvmu1CJzIQmTL71c7B7tczcqQeUBoUJ4JQ7cJawkFMmWd
yYvTa5igdO4IlMaTQUweqEJxyDh7upf70TNEghCBRX6bg6WqyjB3mIuihHJ45hq0oW1fsXnRpUyA
XyXHtv/vk75xGC8cIUfA0o8q8g8dJ3Wao4SdjmfMbvqon6VcrJKgRMw1k0UO5CtqFXMl8oOgRQyT
FDOzP44jLdQmHl0EmuESH9cGYs/jCIx/OMqaT71yz5fzliLrej5QXys8ImLsCLUUaGhqYEdCZ9p0
2nEqCNhMQDjjJACNQrnXh5l8YHppUcLzJ31bycY6XOqgCurYpDHa0WOdKhz76wqIbKtgcwqQ2XyB
inMxuozhiwrfO7u7yylnsQw5nrI4C06HUOC8pyL9+A52goeoGuLOAB/wBOeaj+lZ26JU6J1YRkYQ
G4EvBSYFulLU1tPVGoKPZuht7WFZYVlYVfRo9mRcRW8qPHcBhMmjmb/NFiXdXaq6y9m2zlcESqzq
AKwDNvaP3nJ6aG2EAFTAQEWGC4tKcXAgizXLIVmvP91WsXK8ThGvBJSTo1H0OwMgFfWFR9NhTzT5
vpy3PR8QnzaLs8FvJltvu4HHIU3gmi/KrP7uYuAD3aK0SFTm+HmVS4F+bmbO90p+t3VI97vQ9uhl
37MC1vRJDTY1Uhsa+5w0MmoUqEsiRW7tD8ofNwm0vqoU5oJ9CGFFa2WFHt1iuXZ5dpYGz5zH2se3
+91Im+mw15XqUlz4V4Lp1R6Lh4PeiDwv5EKwfEIYbZWEzr19aPsOi+1qcEz+ehcKvy9wkMMs1Q8s
UXesn4LjvEGTxay1MV2lUX/7mY8yt6+dToxMfv5IbEChkAvhhl8bKl3DW6EoDxu41U4pH3d8XHqK
XiFyQ1MXwDSMza1kxh/0tGlVHyBnW+V5nIOKNrJvQMf95MdORg25oI+H4LqT+/mbVOg1X0S7r//Y
vHXaW4KtBZCNmwZWGt1ooGeYAtw64p32H7nBIMSsqomOwYhAX3gjf1wM2QSS+D8ZJ3F2vf6WCYb8
EBY6lH/fhAKawXGDt3EIJrStJ3/Gq5Btba/1Z8msYwlWTy92dcCunKnzSAxLUBYJitbZWmGTfTE3
0FWBOBfS6058seqGZ7gx/5ikudq1V+OD1n+8uvcJEO11xrHmt71McDV6CRGZHwN2ElHD7LpQlGJw
3wvLuFET9RzEzAuRDzG4oLztQl1XkwzQZrGJMrmYMdchryUivmUlSbr7E5H795ro8GSDG+PvBKhn
hXVwxHbuJ6AUROL4ea5U0Ho0QQ0GYzmuZqnn2gKCIK9c4t+xQ3QKn1LyWCpr2gixhioWu3BHnv2p
IveB0krfThVGQ/h2ETBWSZTqF2bziw4LH6JGieg22GPlJgbsxpwFiJqGt/usJnyn+qi41HqU31nl
uRsYx1TJZ0CBd6eOp2rV2MTsiNzLE6Vt9X/JLHc1HY+0Z0nMoxhoNBs5TH2p9DsWDv8cLnIhFRUw
Zfr3HWrcTQ70lCSVil0KJ4k0PIU5b9tdkFLO0CJtdspmEYqOOfNTMxo1QO37+mwPkibumawIlupr
fFDx4Lf6afALUfmlpOkLHqAUTu1Sw1yGugmjzeSyMaS39iZ2VYHMhUJadqHgMMV857OZlzJUx7KF
tILu6d2vM+n/UFHbUC+nhdPN+SI5hDyEls2DoK3osNb2zPfzi6ZlgABp3zwajeKmFJd/zxiDmFjM
q65Oj3MjivaJhFJXg9NughgyRfXJUYv1YVMxbiGeji2PHsiH4kvR/gOzVo3asErzfj2ntZLoGtGo
s6kRBJFSpUT9bajzqDq5A3Dc1BCT3+ASCW4AppyrxsjBgVrIh7fyFM0Vw7sdNjq5Hb1SELQi+0CL
6LeOdHyrEivl3OhvJprx+qQs1ynx4xlS0hjMRWQjP5+phdgCO8WUO+rKawupXRzRHIfVr0HVCM0C
YvHNbm3rJNUcHW0s1tckJZ2JgvA1xOt5tLoj4zB/hUC9M5KT/Jz5jcdBeB6tXUZ8K1JD1u6vNGZ1
F750+L9rsCCHSXNx2o6YUPDMiAyMqX/GfRZTy6VfF6sBwBi3sQarah/+QLq4SBy9lE2gsQkwnF6P
8hGmMTCzTtu6C8CLdoNLHlFwTXzF4I3UN2mCcOPDwd5YF/bGM5D6RmoO9R9wdLfgMaD50xtsLwFT
tIEgaoCtwi/I6P0CMiJXiVdPDJ0c8jyFXB8LW4W1f7L0mqv5VHuLMcg4Eh7H6OB+0PklL23PXQON
QKbFAOe4b1cFhfwhLIPWGWUzeOiX8Aq20ltQ4hf6wLHhnO+QmzX19VPU8Kx8slxE+9YfAV7/e3oU
8mHgSyxZt4Gu1x9YrDutNYaT4Ea0kmxLhSD6sDQrDe0iOtuztdrcOjS/5gFTuhPPPe2UMCC/NL3O
u26QtwsuqXwlUA+cyl9zFiP3NIHK9+yZTiuOon9eROGpWWuBYCVVvD+n+4JayrlCSh62Ep8gPr7l
xOQAX4efXd0314w7sBju2yqMtB3GtBY4DJNVp9XUOVeDHUOqAlO2pHO0hxeGG+F9P9KgDk0pKdwb
bOdcYa1/XnvscF+fQRP3ILdqH3mfYf+KXT3eUYqL9ywofLENg1laVGSxcEhPZ3Xo8FWZnqhcdjwI
oGg4hIJrcdAvFdCf0WyvtsNq/0tjelMoT95o2rcAxFcWDdkUxF06FG0wPvrZTFzHCU2KOJjUbuNd
7nWBGgjc2E1/xgOZZCBz7QkzbvQMt+W70B2WZCCO/7JH8jcDrZ4QiFEHEbuLM+QnAX4DWaqd7XMa
UR9TDUFSIzIFP9tqhE5SYFdHJYeqld/nhNz+FndYultgvK/kmy0K5G0URYz0hHTjbG/swaUT1q7i
3Zfr2sDtEQgEg71PkTP0XExuAoMOwek1+9cHiX4KPLUfHjAHUXG4luPvVmxSmaxvIX1eEOygCTHX
t4rQ+U2TwWmBfgB9J4F24O8VfJy75cZnwR0xWDhQGCFuZ8Q9C5Q3ACLtNO0igBwe1X9wZ6RFRf++
0Sg+BF4EaWldrD9j/AL1Br8wWx85s6uFbl8cZfQ59zS/ALzytzIAvzboSK/TD29zNNtyDYZQAHB7
+H4uq2E3Uww/fUZDTRuceGxYN+cXm0NdieFSGoNzzmQpuPDScG4FQPwhIBO+Jp1Cl4DSga+fW41m
ydxa6h4N8aHso8HRCZl/WO7fayEQWyvaax2ah/Z7Aih8FQu91y+wdmHNq+qlV5X7reHT2ZdBZKfF
JLR38pBXxKhnJwVl6YDWatAq/wyffMFuFSSSb4ewjQ3thNtZ8XypaNrg82h4t58rrEgm8+ypCtty
i4yy04JC7jLBsDollXuUKKUnjMLUFvQT8F0vvLUvOeWH4xCuDP7bAgWrulpNqwu+HPx5DWpS26GJ
IhD61qJjrm6IE5KZZyqeCVNWiSRauFJZfe41AAbLJrj+vz75C6+JVVDnGGSwDUe4mZXgVbH5XKWa
t5DPeNW+9nWGJiOIihRigBftMBR+Z/zRv6BJKkvPQqZgvwrli2uUgf43h2LC5kRxpkEh8XL+APHy
P2Nr1F80WBnsX6MjLsR2f/2mbkHQl89Vt3OZKx+Ibn1xOfZtqXXLfdXaGD3VP9YYgKGe5mAs9d5d
J8Ng//6HFYAIMm8VMWsaa2bklFLymolFCZxj6tsJFC3G0M8qgWia5x9Z/5TLN2ZgVtUNI62FGS57
X3a/ROZrCZik8AM6IjHGIDwOHrNsApX4ftR7Tzee36VyzeJ1vsijE0KQzJolHHOZAa+Jc9mHK0kQ
qujn797BG/6t/2XNMhLQiyBm2wZje58AHxQF0ZmNAMEqDLSl4j6iv0V+GFkRt1jYeiVYYVYlQLCy
Qei45Wvm+E/NzFOQs/tSONCg1bdEmpLGieOmhae26UNe2NHBrsEdCpWGXxIEpZF6Bdty+lGV1e85
5zglHccVo0m47NWfl1djKGSUJKC9V9LYW4uG26TSbRsiETs0872TsvroUHbnQRLiChSB+JCCqwLo
f8GddXH4F5MVJucaKRe4OjdSEoYrxR8HUs3YzvygbSlXrBZqHfmk09YdExq2j1QnQ4PYDDp4shN6
WdOE6j2EyFB2YxLSzjCh1VUBIQz4meAxGgSOiRXuamIoEXXVqC3whSdksD9JivJK4B5BzCdodJfT
benMRd1mDEppvRXwquJhyjuk/f75bP18eu71Drvx5nmH4G4VYS+dThAg23ojD3eGDgf3u+cpcUpK
VdqB9NDMBM3t8ruiALtYab9MImP3h1lbN5w7jggFpVoQCty1ch9PfUovhuA3U+N40ssLtXe6+U1a
4ZCigAtr42c9DHAzYSnQXhWiyeLyfTMsJAux5sAJ3HAzuXqNrOEtbHklVnBDQgQd5jIeFP0Fc18L
lqunJVDzd7GE9qVeSoQabLRX7eL9D5SRIqgmIF6VhzPnkQXjsE/POgYj3GP37e+JB9jtFXfwSinY
skeC99HRxaAGFG3j+5z2cI7yKPxVbQwzy1I7tHkuRZ/urCyYYFUhIW9GdM+9zO9NdJhpCYrCqXdP
XRQrCyHqj4ygH+E5CNShU7avv3QadiaUt89KHp8APIRvunLZZ7JCPEubXgE3Tqvn/DPOcMrpfq1S
xYN/3ucKLdK3KycFp7xXAQLL43hQ3e+z64BpALXC2KiymFT4JvvFccD4FZ5aQ2ntW7iAviDn8c3W
rf+LvTd0lmnFsup8Ng9mNuzcV7uE3XxqLV+k1YcVAZ/bzAo6nRtyubKBxEV8OvC/pxwO3jjS9kCx
bsDmSjAmJkPnQ114jPrKzEI0VT1BTUZUP03lZuoi7eicVfM010vOZ0Zz3yVY9dJ0KlkWtKlGeZON
9ON8ZZ8vtoGPQ01Mw2ezHoughvMFJIibtrhQaAp5oNbD5t2G8wUuVK7rKM7LMFGPrt78mHFeZl01
JF9GZZ+Mgd1VEx1vtUPuG2hjsTiqHo3L3CBaXmCDMVVc5lIV4y3Z6OQLV9ij90qtyx2AewDtOb+5
YUd3KppyM4y4YAukaQsXD73SsNPdXcmGJcUJb7zuvoMBnAcmKV8dyaApz1/YlA4vNejKn6e8FcKi
hm+V+NLeeNCrQg6TXENYJTawpffBOFHQfcgWPKeRTIgCCUzD9d4eulyTUlyNB9DxGEgKfKXf2oPH
CRhul/RmNfaFj8n6JLh7TBZABqu/ri93HnHNiYTLaS4Iy0EUbdBE5644p91hUEwlJYZRzfCL2Igz
jofHcQKasV+slp2DASoWOo1RPCsfGZg5nnslSi45SvKHVWNFJyXFRVVJ9nE0P0ci2Ysri45AxQA6
nXjUXJpGjRltL0soZZjuxiqVzLPXnMD4f/rf+EBXWA9TU7TqMjQGJhoUytD+wdxReMgIwQ+cb3Ep
WLn2YQQiihqsHktEatDf+OXBwbIL5ox8994NiHifIFjROkVfJq4xrNePDNhp5gvdWUxc7yQhaCVN
lN8X5WiA+IsBeD4X0zHzxxf32jDuqaRlPMSjgWlUUeJRBMvV2/Ut/pkU+mQH09I4Ygw/O/C/PrFG
IekpFyfxeSGY3y1f/Be2v17XpXVAcr6QxYcRO3mEt1Rv4DNOS+spRqFxXswQTcxlx4ixWDgASVrO
1eKzzXkqcc9pP5iQAWbwwxPMKLh7ZUuVGL592KW5AInnDzaFf5paL7fTq95TrCj0zQunmGBUngNl
0fhUDeHHdI5fvoAXWNUiMElA28qAHaQoRsCrQw7ivsKU3KwulMWTzwmCaOWtF5LJHEr0xykg2oui
QMj+jv4Y/nILc06ovnB3jrR0wcZELogYRDzG0g3Ii2BCGcBgogtyCXqpipGbPyoFTWIZkyWxDCCA
X2YRgXNaFn3Kyz1FDMdRjO6eooUhq3hdehZBkSQiP5PRs3M/vH1kcTHvUyCWX6bo1Le5XzR0+M4M
978sS2P+L1fEnrdnNpLQRwQmqCCNpm8/mS0VXJalsLl3oDQqO4CjImwMZlJ6aburVHbXCXZd/cTl
PKcsWyjrhTmURS/o4B6RN09vfWMK/8t59in8hzbD7ichQO5Vexb88n1ja+5nRlh9/7qMXYJsA4xX
L0d1ISmeOAkGPz8mIaGiNYUr0AbAJ6JNkcijyRuVLds5Y2EToEXDOyPQ5ILLYhaZdntfU7P/rSnl
slTXEtu039OSKQoDMgs2rGpyAHXkHadr64KQI5rNnvc6Oix2a/9wWKY3rgBIEbRsK3sngZpS0cTZ
33ytLsW1Ne8yTwLYFvKb4+ujU8odeDlUqkCU6HD5wn9+cwlrYxGFpCzjosfChTlAFw0awUXSGnjc
Jr3qNxAlzgGZuJvI/iCto2Ur+OpH9bZtlKir8iuZNJL/na7hgDBrEwY4pMJFggKBqM5qFgFCmiXy
U6MjO2vXVeMOp+aOFk5FtG2m6AuL7ykkJtDFcts31K62dxdUQQrFqhOOcSM3k5B49fkjMVYejomT
L0jN+MwpF6wh3+UfU4CKsOkX6IEBrgtqa/l6yJfCkj26elLsqyxryzOIAtqaZu5W9VO7pUrmWu+o
JrnlttIFSz1cedHScpWb0Bn4tKyZbRhdb+3ntcu8JuMY9Sky3fLUbqSR0FfGH5Wh4VVvYP9B3NSe
D4uLVXtfh3MV30tXjeuOYRFnCKXUIWu2A3lnHJ9EHUUy/wstode/OJDjuufqKO5DP6SiXADs6KgI
Bgfd1HQJ8XDD/rNUkPtE3gYcq93Rq5BVCNSbBHP1FOp0iUuD8OUY0x4TkxV/wdNkf358MbuT+lcj
sKYUh91WJXdl1EUDnW6UWiLLO/BJE3rjEjzPVzV9WcrGwhBJ0vEqCMsRgicIllqJbDJUZsE5LKvY
WYqDrHcl+FfAtJTo/ADpcLm74oFK7E38u2QLVuyLRIDS2IqVaO9Y7lTHRbxdJeoZ8Ido3CPE1JiD
2IUYJw/ApQdJsauu6CC86KYVgIZpMoJIdxG/I+tsWA9g//E/ibzfWdLFq1p9/3J10qswY0jJMdHp
GtDaCUMH2UgeZ8HAysVbxz5lJ8Omi9wG73qAEIBuHtm3K8v2WsvuRzF7mtY6idqJ15sqTfM4Cn00
r6fb8Jf3UIjBG6+4tuNOOEVzJ4nZJ/sWxbTlSb3cXrrLLMqYN4qdwPMHVw1P99w0NZkf9qIpFDQa
+8XoTb4ZzxYYCXbtg+9OSTPBOiWBEp3JTt2vIpzqu4VaWOG0WGjzP9A59VKkx/lpspvZOywOv8Qn
dU2iTSTCYPkWzq1BG8x3AckbPHpSQceMx/hsvJjSVed/2R5fzIEDn7OcK/Du0xOKQJXbuZJou3yw
ld00lRntyuH8wbhepZWavSQ017lekwaem9W8QYlBFP355DZiRCJLlhcApUkNMaPK/eu+cC9MiEr5
EwOg8B9BwKRJ+eQkq52waUB7ASBGpJeVGuCwKSkTo9beDNBhadDMAWJ+hYZgnp8Qmzmh/ia0Pl0R
8/nHTJxBCGJbWkkcQJCf50MzY5A54v2LZuIaHrnPnBA/MxHrkSZfbaGpFZN52TkRiAPQmmPhwLV3
9x5FYzGIVdM+E2E1dmiEnonCYnuYfzv5r9+FmhNkVOGEpMiKL3aWuzpXdgqAfG6KBTUfIfbvNJWw
H6wZAgv/w1lTBoKeQe19VEt39zxqF8M2pM/uhIaNKw+sof6RSX0t0/MWm0fp8valUMdV+yDSvh6X
9O0Z0all3YIKgvIMw8aacHFIut5LLTxauy7B1PHBBTOmbH8Lc0J0aZtTFtt+uYBMEsR9yXiCZcvn
7MRtNXiRPNFeXCa7RTyuYriFAj0+dVfJuBdsPh7IJb5ksVYvxcRJsMLbEYZXXrkFNx0BDatRKJu6
in2BSLvVhCnyWmUKjB0d2MlwqVQCxki8pBk4zWY4bL7m5c4MqZfxaHa0KzmeFCDX7ymwFToJaQMy
GE7D1gBMXGgbtX0wtm4PBiPeYlUeFn8/5/UBiJzkai33S7Xdb8/93/WrVwcalRiXANMk2dtHCp5C
QHxxF+RVxccQEHJgUwZ0VgRdoAQKaAODBXnXf9M7eQ++F8CtdzJSI7QGxINTDonGEEDoqtJIqT/i
VV/vkd9hGx7074E4dsVc1QAs7JTdJsjrygZWgUfhx5qaxdFt697JEcfDg20A7g01jTJm2b3bAvOD
+yrq87SkZChNpBZwtaZxwH64rGs2Ha9W8dhFOPGIWL7qAUUlLHOPt4b+hzCIiNlnEhG0DKw+BVR4
L1zLFwIWhQb5D3LGGqnfQEemIbTXeM14DLyWPIXG2NmXgPB00l2tUBihJAv8o5If0Xxc2lXrR9Se
svlY4BfLyTMXINcCDYYyoDmbNCUXs0db9JUN0+/+ZsR77VzZLvrALJJohiyx4DTJ28rw4DbkXqZ9
F0yaN3Hcf/m1+D0roFWrXLM8htBRxjI/85xthYxaU1IbL+0bSSKJ71SxoAktXvz7QYDKMqbfxjif
ZsVXjtLQ7XYxextdqFj5Z/O4yjcB2bGAMGOOjhzDUSvEdzHSGmjArqAF9Uw4NHoWPG7Q470f3zbf
bomaKudoaFL9/b5dN9LgtNSb/GkR6KdmBkvdBerB5yY6zIJPaaVCnMFVwQfXpADhT/w9uTEsB5fx
GwJbkgd+N0Aic5xsv3PFZF1Mtx0P0ejwwkvg2fuI3TH38NGS1/TJcECs3WK+FLclKnVCrsL3VW8h
LP582O5zeJ9xNBh0RWpcQEyf0Ull9PMPzDlL4x27lGV8h4s/fxeOjyz6tOCWlCnNpSFKC3raDagA
WbBKQlHv9HwTeD/q9TP05R6OCqmBDItMP6xGtHRl0qMSJ6AnY7lEMfUPS0mo62w9yGJ7WMkrWs5d
uEKU8pKDNnlRLGVsJeM/UE2xIjA9fMtVOEmW07AYGZOGscqT+ta6G8Ppp39yFsg3Xn0hiEutOQp6
EIrz8D7/SuP3dVWoxC1sOyrZcKy5IGfvUeFiaW9zJMPZIdCf5irAHF2RGPlBdvnhG85zqBqrQvIb
WMNo8KfYU6E7yPLNMLKo33IyRBWWPIs/78NP+TCz6ZIldbTMmW0mIRDBpWIK+ll8NAYSIjYoTenR
WWU86W93u6dXgsRqiTAlQ4t0++YI+m6e9mvKdRBeX1WjxcDGpNqxrTwVxICT4BC5YXJ81QoxOIyS
TfJRVvu3vVHaWIZiiwOxoq/YkDuvP/0Krxxy+D9E1L6/Oh0zANy4YHW+hXAXqO7bWaPgxLslKN7f
YLfy2b1NryExHqdkI+LjEye7YpUrkESleyahisSC8lkqkGvHfqTNYn+nL3JNt65AXCzYdV9dz6rT
bjV99zmpwdV9+oA8mtBmHXkmnO8w6XpY1x7GshqAE07eznH5yfprBhxKFszM6juQqCaGMjzhF+lZ
fRtD1s1beqOySY9MFOSVlmEOibYf60HA5GA1gsrKUbiFv9k8lzQF6AuzTIbsdthSM29zq6WjQqJQ
TjQLEtTNXXA8MgbcRZj7UoaQvO4tRv7dNxiXGAjzesZuTZKJMJL8nujAzyp3XPUKI8DMDZnNc/vw
MQbQyvC3mROYrrpSDhwHKx1ffztLJZHrLlYUfhVySnHJlR0nCfpGwLRCknVE70lLP1xmkBSgg+Cr
FmVCYttVqMJECheow8zMA1o7An3Z0nws3Tbhi+H5JSejkYTnp+9RTtQN91f5B7GYuQRuIRWW5knv
1dDAn2XzlO1JP3n6pMLeJulyc0/NJneu05HuJ2doGOKHK3MpPfQCY6irUJ22coVVyonPIalHT1FK
1CfZADV30txs2eSiye1wi64oCmCoLthrbKecXZkEHjLLDVgK3N8OJa5jsQfhQy8VJN1HqpTAfqHL
yO6qd4t4U4EJFjy7LxL0dTThNM6CgzHB3p/4xv1dERbO66vzrjufIPYvnv9sXqtPU9kfCrMP5JO0
W2FtD3f5O6Z6Pvr8GBa/6bbIT+Rev19ObXKnx5COHy0lNI8tM8ACgvKjX41k7ZHfqABL7NgLTpAh
ZieG1flwBBZfgrJEAu/t/mbboR1NkhW9R3jJzvfQ8z0axkAAgQK7b1wn5dk6EM5fWVCVHxfa+NKF
mfIIRfArX2bgd2PRgkeBrPFvDwEO4NO/QVqTPd818Phqi/h6rT5F1I4548LcgedPOLQRDHN1CmzY
IaGrIEas55wAbQmR2uiotBvZKtkQM4Wq9bojsl7VbNhjWS04XoS2gXt5x4e75UwIin3rdgtSQapu
VdSKlW+vi+oK7TVgmJ++1O4GDjcGkyypv9WAxZSj1ADHTeZlE50BQnnTFWqn2uaPRRinzLO9GbR/
m2X0tuKelmrNXsu+ysRiJrNXhx99jlDFLGV1zIRl0aMZQMeHu3szNRvCOexyRErsN50ZYtHJAyrA
aFUG4rMF9ogeiqNaWIcvXC6e9OlVfns1Uaz24CBimgV0x8ABwofY8Fktm53S6nsUrk2tSy0LV54K
KzKocmwUydM5gjVOJbaVpYruaE0UKCR+AZZVrfmN5V/v9pcRCvSaLQ+DB8+T+ZVBF6Jsg+bNmNdg
NXuTtmoIRdvUcZ0/JE+hApsLwIb2wP2jnU2kaiygwf5XsjLj8D9ql9NJ7LYDMGZ1NX4GpCHwG1u3
i5DvCqhbePVVX32ZCEt6MEUvlg8Y3zWXSfruuyUJwJucBNpSka2Rr3Oq18p/Y7i1P/DIUygx4j8o
fkqrpqgahIqbmfcHWnJTmRAPQe53UvUR4//j7sC+7Iey804FHAXQcT1zEj7i1QVef8kapycO0zRy
5ObbHUa7HAqGlazjeu4duE6EepB/6JQtnAcbukGnsCirZDjIDxKer4jz51fswhf10s/D5xyazp6L
ZwSTtjxZ6RGwNIXYbpJftZsAIH8nbXVlgDrONXuL5265/P9L+v/2oP00c6iRqFqVeRpH96qUS8dl
+ANUZEJ2lyEEwMtN6tWuRuKoDShX0LwxrbHXZh7YHidBg+pVWE8QcgqAW5YV3evIyakoBMtRUreJ
8Lf8dBrJ10MW4/bAcKKv0lXhtm+vGxlxJ1Tv4wvCKlHuNbV45x0kO5Tp7bSZCLhh92m+uVrlp2mb
ffHIsTtYk6t5mJVn7Eey4W5yOwTYl8c/QEaSklqq3zmwm5OakfwG18r+r7yOf6ytcnVjx0suDgSS
pKLFAMPoecFUF9ApwTbzxU1e3rncgvOLEajU93uFZWPvpedKIGsga+j60Gspud2dNxMrmsr6T6Rs
+foq8ATWn+iZzvZqdh3ZxBxsInY/Xc/gn5CHRUABn3MwD3d1SVvhKHoq7Y1qJ6aJYFn4ksNhZ5TE
uY2d4K4Ek62Un4SZZ2cd0zbOx02Emt9zwc8fph+tn0Fr+m0jP1xW1MgNsALgmuRLki7moIX972x2
/0bL9uYpkK3x86Vxz3UourJoYQCwN9IEnSBLTlGtmtai4rO/afwRhxcYbWUM459l9Z+78T3uESoO
jGShotUUKoWTqVjrdwCCkoKgvWFd+nqStFBO4QZKaT32fr+0McPMNPZnG6ySd/y8X1xfTO91jUnc
kL6hxYvF9RVAzi1m6IphbxjroSwUQ1l9TGwxv23VDB7wM7XNxWM1mkKvN20q38DmdNbs6sCBVA0P
yeJ6M70wlrZaodr8+0GE2Fktwj5MEuP4YqNQNCj75DfI8S1GU6cA97MFNnZIaaaL2aMH6+PgBmez
+YJfMiyQF9iDYtGM0Qel/ZrJg8V7YYky/9XR9tvxdxO/raXVkefu1A0OJtpjWjslGNwfpDwYYd75
KXR0Za1YQbi3Dx/z7FBctl9egOAF2CuRpHHK/FzbyZRemPWCZ6vsF400B2jJDv2+jzc6x/nCr+ro
mRSMR1rDzoY1tMngZnASyg8C6p9I4aXKS0xaogAvvU1aiLq3wYSjwvl3Y67wnK/ZnUb8WmRwRiFM
BLgZnVlCOZPoH/iNf578dntXTORZUTyfqt55hULXUcGSEJwFDm7ia5lprtjxIgnXoCkpEU5fBGFg
vEmDjIu+fyXSvMo9Z+4GaxYgB+z8TQ8fuW5AAe3nyUVIDqGVbJNRt7/H6QZJxgPppUcGOxIbnevc
objFfDfJr8qcC2y0PdEdfHVVl8vTSNK76dNZQU4BLlMBSnovSqbCxc4hZJ71Cqq2trH+6CCHYcVD
vQARaiKbp5LJW4hAqA1V5PMB6O0SJUrE3HXNPYdL2YDFIEBEqEXZCZ/sxqTnoDV+dtfpBh88X6of
rtGfPJQ1uXDm0e8JT+vBBXYhhmpEgF6QL5AClHK8wVxj1T6C8MRtrjTnVzxuvcdBwJiHNX0d/+eH
IbKlfrGtvT58q4BZufMlBAQpylA2lpRa8aFaN92obAI2PmV/Fx91xGZcLJbJvZ/XitzzR7I9vj/3
yfcN3/6AIVFcv3khEW7QozoteKJgBy26XrHKPZ0o6dLfsUOW/ZvI0vWurSd1h156CkODU9ZLRXr3
W7LnkKYL7NBGzZVdL45f74sixkmzw+m7JDb1a/Q0vCMeHgKRMJnHVQYX/CihUCEraR7SkGQQhoPY
8icu0buKRiBQ0YBOQdSos8Fhs22kcGmPb1uGb6u0n3Cq2mY3bdaVxQSISg0T1EDOhJRjk7nhSygz
uvaETowC/VpNvedMlYBn2qccZ7oatywbe4Qhb/kIGEgzI8wWlrd0TfoMMpgEY5ZbSeG23nJXLlmj
4GV0r5HZb9LyztgW1xDzIS46FTAhLUoL4GisRmoaO9SyRgDqol56vKEqWq1HuDShxRslKHy0MdhZ
aB4Ke39p3Rd6wDpnGmZG8Nm04g4INZyS5KiFnUfO5ElbdDtN8b3bWf/xitxZ/keJ5VuU6M4cUnmt
qZvnVhjbGQmXD9lWhaVRyIbM6DVD32CvOc+im5i5oLEDckaBlFs4qvg6plcPsuxcWGzdzzXXqVPB
h/8tIrKWmH0SFwiSrA59kZU40zSi8b/2WkFUcauiey84GED1k9JQJycXTCg0GSAp/dfYJL4ONx1L
/wtNPn9jBbqW1j6IlE5a6F883T83rIj/B9c8h9WxI26QIhZYSi50JgMP3SRljlRObje5+afdKj5X
uz5Asdltmw8ok3L6nI7khKOAK34ZVSnbGewiLflvg0PeRvYu5fcSExQGtfXZWrW+p6tN54eynHMG
/ieiu6+ICe6xxrY8fKaL1SutkoZCq6AU6OAil9BnYViSgfZpC750ZCgjrM45m/qU54726Jtwd71L
YIjDksVjNtJ0iRXjoO5SddmbMaoMDgn8ZjqeTc9gxR0UsK1J9IRdWElrHonMJNR/SWyj/8iv2tV+
ZOD4HcWzhMtLmjucYcDeO1gbe6zxV0YF89Blx/fx3wOzdH3ohe5xARZyAgtvsILm5RCmMPP/kFos
ImQ7VGcaaotLI0vu3j9/ncsCmLzLvesNDPurZWLyf3zavV+GnYKBlMfDatHA5zEAiqU3MapJ5psW
1TUTBv1o6rftzazAIZrVtPNl2oBZEzf9UqqAnssGaGei/JODOq1+fWKYdbWomdLzZ2yq/mOD4iq3
tD7xtDsaOOtq6YnJlC5Po8F0qlgGD7D9UsREja9oUG/4j/ZKKI0M2UvR7VrDO2ckP8JHDazs5WcB
Tb3aBA+ds8JI0YZCEmyK9W6fdL0TSRH/1C7QsBDAPgc+yPzWth52a7DQnnL2IB8BOjvJwr3ajLW2
T2bNMnW24TEAE25SFUP2BbEVM9q/Oqfs/ZJ3gsNlwuRtZukigqcvU9w2VkgCR0f4mUAjeUbwYYHs
deqHMA0DdyhKkrPsM8iDhayQpoF2O/I2yWezvx2raF6FxjK0B16ySqCogDcH49deQmCjv1mf4Mng
evQqM2SYxI4Rc3+R25Ebfi3DlDScphApycvYbwn5eDsOkCHtPeeGORsLX5x7qXzPalqBcZaYm05Z
x5t/3q58H7ArD8ecpyO56zUqF4TosEE8WELDg7bb55hV8OO4yeBI+0hxP5F4cffVtqEMtrFNhT3B
PGBrH7ibBmnKztlcJmQOrfkVOtZ+9BMAFqCCt4D0Lp1NRAqjUQ9hGW7uZo5EhtnudXLA+fk1SghV
ekclw5GhHhwUfSJnqK/4e9eEYhWR/4k2dAUFq9N1w8fMnd2jaeswlY1nBT78WlDhiK92L4eDnIux
3hSIFOTpTQlt8+jP1IiQi/MTYkntK/QHrFIPwvheoOIThaEYPKRats2hA4YP6aj+0FA5ZZtgdF6g
Kk9TwUtivh4OfKIdeqqEu6CC4+3nWfuuhkeX7JHGq3seg1so4WtrcL+UALmPYE4lYTgkE61sJhWH
k7hjt1T2Fu5U1dAXzjQePIxR1mthU355YwZLkkp8gkibOVhkFYLYnWvZi0/wA9Sc/UgO62G+Z4ze
yqFa5lkONPluF684bKbt/ctj9vh3PEhh1NNW+gcB9rlXp8iNWLz7TLd85RnuKfV9sWZG8gmkXDgP
SeOAVPF0nfelVvR75a4vnSEjZsXITrArhxx4BA8ybR3YnMm5WzDt0+ZawIjMKq2ybKCrNEPASUgb
THYVxHvR2StSQm9bn1Qa30J0kSc6rf7DyELruJY2XlhTqj9R0VH/IE1bJDTQXlrT0VQutMB/hOc2
8Vy0RHIjHl+HvAQ4EkVFP/tR0s2TEGInzbAtP5gf24I8iKJq56ij8brDYvzaJQOtSkUukspcYmPN
piJzt02WV7bn0n/zaECl4Nmxmm/+YNLJ6R576z44+21HGgG1nrik8YAt2GgKe9+m07SOHjsQ7HKQ
vh6ZVCoBVwtQHXVJ54hAbGY2XOw7lWHJsk63WoCp2q97/ySD+alv+4Ca6hwm7Y+IStsT6NJ1/wf+
IMvLTbyXAKjcxEKVjMQZGW9EXwltrAZfN+w+Y9UZ2XrX93Rwql2OUSYdiWbMt3Z6JVTizdatn8Lf
fixXpgfDUWDzg2OLy7Q13ap/gI6D/kBxte2rzeMxAS+HzwHm4RST49dQXqDJjAtZRT0/HhpMTwpl
b3u9mJaW5+GCXe2g9zvWUQwgE1ti+ygnHGJv+emgIoG9LGvY6s4HXNP3FmvXpIAmby3KX7+HoulQ
VChXq+Eb2xQvd5wEW/ezx1bC2CMcZaqmGuCC6qybGeItPxPuHq/OggK/NR6BkWN8EPFN/pOGs+wY
nekwQfLhgZsmvz9bsDmtHBrYUkJt8YaFSiZXFqZQyyv77wot6T8iVHmRgdb5NaYkvUG7WjTfOpfl
KBbu848KfyIxgFZgtdHvONo5uzIElKrJeoSAAK1tL7oE/3a34h6/uyhrjx+dFq1bQJ0m3KQG1t7v
jEH4nF9YzLX2HHi9NxfFPcD+WRSUSytv3BKt7wl956s30F5i2JeEVAS/x0Ip3RIna+JRVChP1EMY
OyQzqgMO0t3BFkryzlwx3KTq4b20TwdF/NLRSWWx0Ujwvx54Q13/q7WHy2gF/m3Yhn6tUzRong3r
DnqYKwNxi6l49OoeRYd2oef/nERCxQy8eRKju8mgSxfWfx8o0hrV1EnihKU72PgpBzBKego4KIs+
QJ+xZY7K9XetVsRG3pexe6qF8qFOQvAHuyh82lV6Nu7Sd+SgUhvqfI4Vitt0OgymsuHpofNVOhhu
+fH5Okbo44qfzgci+ThkOB0fcePdIbJfEId62gmXsD7tI//XpHFdu5QsRsVxklY59ya4WJiJJjDX
2q4yssMiUMhPLLAcrQKPAJWwuvWxnly1qiEZk9R0sDrBFgHrePkYK/LaRj9bYw7mgRjChZlZGRAQ
+tFP8i/PaDe6ie77dTpEOEeRD43U4OY2oykyZwaDkKFbc7MdOo7MXPu4UTL4Sly7pvKMQwti94cx
keEx13CdyXmH2c/GModUS1DJvc/f9d0oDoLrjiWlE5oBf7ygvZ4scW2Ld0nqMAen7XKBOVD5FQOL
mcUrjxGvk90B5BnyQXpTsci8S6GHCqhqNzee87U5AazS/iPZ43P5Nt+T5hRNGzdwaKYhrGOYJFDY
I1qml1JLkaYojSRRL24xnrInkPM8i6eLOf4WB51rp8M6TPdrBCu7YNBtCaYcbzImMXkWlZp9YCfu
idXeJRjxjlL+pn+0aZ0iwXhiX9Q2fxJkaezbRx3lY01WF/6v76Y/KGtn2siteLliAchWq2ILccvc
7LGZS4iZvQ7i4kbpb1sH2ZM0Y/GbGZFLrv++TvVE0a7fr7tZW2coE9wSn9cnpNCh4la2nQFKpGar
qkUeVMpeoMIrfpM5ojojBvIMCl/eSiNkBkJDJySJE/AnhrLuf9rxkcUReiaduSVYoJhYRwmETfJk
kP6Cfr5uYQr0sStCMp1iHmBL067jngDjldYsylxuiTD2PSXSmneb39kNqRiHcdYawKsQcb7RPzU9
QLLpOV1/9b1EKI6frSpxiMWX+HhTNh6XZNW5I+8Rv5NZ79vRM90ZeScIiCJCvog7ZkPR74954/GK
YS6uX1o0z0ur3SgMuzSvNxqNSvKaJZpVJRdcqD56rj7diotodLSEOhYydUHzR9sGacskONwgiU8t
dYlYe4aSLOZ0a/9GRRdyVIG+FXOqPGw0qoxSsEvmJmmbjsxQVS7zTnkJUH7JfIJloG8lUld9XV4F
Zb8J8KJfwJoKPb2eh6XHKu3QC5XkbWIGWC9aykPIOtkCfaYT4e3n7gCuywmG+KPZnuLcs1kDfEWS
LhoN09gWirncoA3AtbRti5Qp4ArnGiK8UXmQGKyKAoUKrv7+InZ9X1yDunpJXRe68WC6jc/oJ8f1
5rgPHbNa87vk7xJ+5YnbZRaFC5CFQEHlgVE1QaCE9PcjBmzUs3Qs5moMu2/PXq6eMTy0/+4zwnom
PVtic3cjgv2uMB3XhpEoMI/qJcNSo+eTEFN2RQSWo2zxg9iQo4E+foBf0Hv5ssxJAYiEMuo6W0gk
pWvP1glfLhjfL666XSuDcwYSSUzUQXHOQFZpmmebVNSCAf7X4Y55Vmg2TcCsJZjqoDcs8CihcZ8l
fLqmmT4o4zxBHuAaN7+mljRructzsh+Dcv8velPMmFFkJ4VJ4owrmgLclLZUXH/4odsT/jPSFwWB
FFkSuWgEvJUiv0QQObXSIukeGJBT2lxzwFp1zhVp2JBmPhqoTvh287vmCB4RxAuZUQy40cuBJ2Wj
Dphe9nGpQYvsqyZR/p6NHGVROIuuDXcQEvHvy059q16TcNAvYteav9eUPy2mTsZVcwRoRfRI2+h7
Y5xdtN6RlTlEfeWsYneEXHhss5pGZE9NvdLUSQwiYXjbjIW2LO/gCKGgGvZPkQBqxbUuRfldzZX5
moFxsSIjDbE8EoO+SqjiuMGTMnaz/D06f7OU9z00jHUnfBljsBySxjIBH39n5Ca0XTDjx+ccbawW
l8+efOo5jOPs6rhWDwKwU7gFNSjf+4Q6KlNnxrieyVB9JK/1yaqG8MoaKIj0tOr8a05Y5GDxdU9R
VMxfq1ehSMQWwjk2JwDclAWHXtEQj9FobCBKac4VIVOmWnrk0XBpmppPvOtymfDZhuxJuitoGiYd
1G/kliK4275gT4Qe57sDuKodoUGN0PyzcxEY4YJ9F8WVgfTOjrmLPVEq8Li2R+ovLbc7UFlRojuk
NrmtPH+z1/Ly7pr+O0n3w+xEmPqSBh4KZH1k5dWVfeKgOuYcMqKQ4RspByY0ICkp1kXuTBtolyCY
C0YwpTPznj7b6nrxY6RVzqnl9SEJQySyZap/69DUFvYtl60Ppn6rDc05QavkHgrFZVUodUDaaSXo
RFfUup5qYjR2Ih3IEIymicxhDF9TuVLxWqmwpYQHwW0HoY6X2pZ87NdrbM5IYUpvqNY7ths+NDth
ergvn/THSpLGNSeNyDR5mlT+wb+U0fG1+PD8cByfX3CJ1TvJMYpK9OkyyhR5VEXSSJAIzjXPPtEo
mMRvcijbSo+QiM95ibu94jvLmUX19yg2f3wJBrvIoL1tCdTFI+Hf7WNwKvpn1+51X2TOmIL1+ttI
cuRNN9HrmwO0mb7WvdK21J9Zpy+tM65lP1MImpU+7NRgDXRQOysqFN96iQ17Zld1Ti4Xx1ycCmRi
svZnQDfv++rKKkAzlEnKqV85k7i6DDafr+36gPnttNX5kbZD+s6tTYLhLsteMc2isJYLkCTS+XiA
IxK+Zo8fDul2GavjAEN4/jaFHCUAasZWWv7An10uywpfi4qetwKMxrT3RwgKO+XZizCFsaB/q0DQ
KhAn//yK0qz57tNDP69SefuhRn44/TzqtLY77gy3WlQ9A8axS9ix2V5ubIOSDWXq5MHYa+VCOSEH
B3Wj+lowlvp8oZoI6au66XlQRZUI19l1x0Jrd7PC5T680PiPZQI7dIfWwQBQTFs3diVuNd8eooLi
6OgLw4gSaAzN/jyMiVkBlGJzG2+bh+j0jWPoOPI0kolAtg8nh9vDyW7dnnWhcdTbQM+exZ1wpab1
xm38y5wWgRRUDQl57Qx9V2cOYnHipLlxjLG4LA0MkaTMQ0E1ng93CG/MuezaCUNE8u868tY3lJ77
RWBQt1loOVjB4Y6VXUGp5M7vAh8hfONCBGbV+AFksJPBzex/9rs+InXBONlfcECuwMX1NCNKVdC4
3eGggJRkNslAsfXRxKdDFnxkOCi1tuBU8JAIezPK7FaX46Chfxa5ayJLmWyPm3e8cv/HTzkdUwHc
YldeUCDPhUhFmU6AM8Hr4IWnsTDdROmSfxocdJNACiCmVeTl5LFWp4M4yaTEi2VG75uuSMt4XtZ7
7wlP+UKDcto5QOuDMgh2Qyar7qeH30/v2qY34nSeDmoz1ynBzZ1IB23317jKH9957M66GQ8ViYi2
dC4zCY4Tlr2UDVtwU6MHFK0yTvHzgEThlIiy3QOnj+GxTPFy5jWvS92ez0NjPxObxzbB6ls+Bklw
nsKIjpJonZwEiWKI5Zs5FO4SGeis4nZEvbdQEgu6kkD9/c9MOxUteg4SiL0W5AXUAvuVoJlepfLm
Jk13SfyMnEu1MI9czINlXM8K0VhpyI91j/SdOjZpsuDK2wifoQsHQSwN/FyiDQwDvQDthgXn6aBn
Pw0hnxWKhmynVuD2IUe22IDhYIAUccX4jdFoXaMXR/nIv1zEgYtjL7HPTndkPruXMgCu2FVeL9K9
c/pmNqm8rtvg67zeDeguH9VdycOBhd841+IvcmDLeh+oK0QQ08ZUV8SoQKcqE4NZq/njNvVKGtqh
eSn7uBkCk0RnNWoO0NDTRH/D7x9+GKA0A0MUlJvn3aYawZg5ee6za3LQXPBtUz+c9TyE/PMhHCRf
8WY5WIES0EApDtr+TrCn8SyDDdBlezCbZwADQdBcpe3Ar+nXEwo9XgSSRWbBCOji+9EMGlVpmmdi
7gPbng5Kc3k803JjzTM6Ik6DnrBpvi8N46M0wNIXKL+GujHOumAlD/G79RGJFECIe3DX9Kbumn4S
PD9wnH8429tEKwxVSF0KUV4rdBbC7nC4WjEXdXA5TuLzybBj2G+6tqiL3BGH+9MmBYVRzPxNAnhJ
pLmTUstJfS9ZvMLpYwESPFbPs4z1j0cDA215pMUYyXnOe8lznUACdlv6+5MgleUCw1jy3XrMYOZL
rIYbjsLNEpZMZrIL20Z48j/t22MRfK6w+xMByPD4OTzkUiDm9YALAWx6X++OX1FO/MDcQSkboM7q
GkvgRcjcw5ppZPjVEG6vjuEuEtaTkrcRyXYDIVsRrpN4weacJCXTBaXsCz5rmdDnvjmLQ0z3kDRW
C8+mxvUq4KkweUTQZCoqB7zXviDolfp6Ow5EX5lCqC3+Q1KLDycA0Ht0ZZybiFuaboc4x3tffqOX
njWCPVp+KKRMBDtEvITbmdARgR4dGV5EdJY5lVV0DiQDS0kvmMdM+xjD7hwiNf5j3PHuhHxXQQSg
zUgf4LvcfIpCgYcPWNrsW0VuUJheyKeHNa0tWZ23sBHrbzPRTO6XTwXlRAib5MIybvCLSwOfBmCa
/C2xXDRp/45mlPY4pzpy5NqdbxoJTSPsyN3ecgRdn0a7aAiECaR1Yv1TmHDwxq3aHzkbkxRp8vLR
un1DvahQeSiIAjT7nuKbQQwJFmVaAOP75uvLjtzrfvtES62TzrWYey7it5utt7YrcJBuq/+UtBGa
Z026FlxlvZJeV/I40k9HCJ43+R2GOeINELOSBi8agW1Pj9sZXdRgkeeDIebghOHiy8df+ZTmWMzc
pqAuKq0xiRHjsq9dfdBC8M2AiLeZNjc5FegZAB2aeH1oNllE+PY+zy30SBpKV8iYwzYaETd/KYsg
UFl0ScjCw97PjCWvrbxE7CLbkRc90IjyQ+R2ixiFnJSpeAuFfzPbwxw9f26TnzEgnhu/M3PDoy+N
jfwqzNue4HDYK36fTZhb+iILSBMcrB9DnIsXZr/X4tEptihFLIDBzuARJgpCmeClp8Np+vQz4hO7
vMXQZG1/hreil1Gx9Ip4OaeSsbbPeBi26ecoehSUCoxjbYTzCF04Fr2Ux/ZaVFpVJbJAUlWdJMJu
PSULbqlqScxZ8b2iO9uex4fOCVWz8KePSuxjfmyhT/aLW00TqT5TtlRxMJVUk2+DHdjb65yb54cH
faQ0GNIUGboP99DOjW4oNxqfyfaR5QeXs4sB8vlLtrhWWoURjLzoiXIAUC4FheUMCy9fuEXNYnuj
eKjD2iHD/iUFWijBK60sWW8zqMlJIiMamrXYvQmVFDPIajy2SppRXtom2EApvQdbCXdPuoqRzrCn
gebwAdMofqThU30duam+sHOqk1qOAF/NI4b+WR8bg4oX/VdkIXaeKceFscrBFTQFylxJYJaplD4J
jZGGS6mMPDNpFr7MS3O1JonJVTrrhR6f7j2iMoF9FbStxlCUGY2YA5sI+kNJgCqTHa4mN5GGsWZh
pS5YSln+YBG0y9kUdZb6fNAVAAwQVvZZj+eCaoxcq+FWsQAXFOXe8o//saFbHyt4CU9i/LxM10uz
FtGntagb9QRPx0+XAPAdGKxm8BSkaVKI3OZyaqTEPOlhsX1fQnF2VT2nsF2HgbVRbtwIUcgV5wDf
RybBu+C18iMfQpigP55TMsotSC730Ftv0ATafIpRnSyTQq4kR+iHY/6sIy7pMUaxRVR3QCgR/g2g
8s23kppO2avJKPeLaxZTx/e9m/Qb5BPCCn42JLTS06BkOmxQDNkRv28WoKLfFbqCr4RBkS57stM4
hXttTSEeRTrDEW5ag+J7Tc1dEvAjzlNnm2099P5iaLythhOH5gOwmD4piOnHOkg4fm56ygNsNoMU
NqXkQCyO7t2imoGMxXcDfJDk0ZmRq4pFoulCtHtkIUp+SfnU3IzsNAZEzRq73Y9ngLX2SL7+qdUv
9lJYwbUIAHmiJ4ngELHuU5BBwbBwzQ3aOc1TJWzg+rmBusf20f3FbxjnVujkRURsrFlZLHnsz7Be
/QmRke5Qj1VfkxCNEu+zquRGTyg8xZfEgHYCWwlVYurk2VKEcs/4JJwZXzH0qIp005BGcWHh8xS/
w+YFYtVYq3K8i2TR6mHkpRpfZM6KP+qs+s6T5RVKFScWmCcyqHdALYt6ZfUgz3VTG3R1ylip8isu
R4pVzJiG8iAf8iJvwX0d7hHgetzKQJLfXGL6hro0hjmMfw1/qmO4OXKke9tzszmODBdSLVHVJ+yb
uu3RixWWrokp5m2fhyUMmuXs9VcK9q0wrhpwXfoWrVxQrOoW6EXmfP0/PJvJpONO13/CQPeDKaN+
TFlbFQLXL8yqRT05eLdN1FLk0cq4SEh9rEAnoTxKg3SbaCTPf5hdYVn9l2a8RgcXrcjvjf1YuUU4
HlgqRlcSfwlCfeYq1CCFzJ4w20nj5oly27Ywm1SOEPlE5Mw7AMBxgDEGWPgZwr8eKAeL+CK0/pZI
C40sdntRixF2HN8TYb6y372ggp2EDehlpD6jTySEQWGB0ZwBwSn4CVb2WnBESdT520XzVw3KepIX
F06oKdCgBMro2hBwYKbAWgxmYK+CdcTLkZuNbUvcJXdWxKMGgFgzVvuas1saqNM9OrrsRKGWsOVJ
ncL/dj4B8U0Li7beN8D0cq7HRh1pGKKAXV6djl5ujf/2U8A5nwwv9PSyo7x3iwaT285FfMhcOnii
HgtPK+Mrs3rnFR6j0kFo8daYgl9a1DTgvfuYyB0KhXVVHfqngnq/G5lqw8KKHwwfLxjIU57oHul1
ydk2/p1QLqPavSJFJ++FmC7XGjnOLSzzHoOBo9AQG1HZ+nAbaWTmAGLEb+DZCqOcTzkFwUUXYzIL
ihTpYGXGht8FiUpzTRv3WiSAZOvp2sVk58dKiMUpiwe7To7F7b7qmt5KvVHdF0aheiktJoWmrhPt
DmNjjc0CMVkv0WqKJKYgCb2fkSi9QbpiajNPRcCtSbC3iU3lzFPN0nAEn6eetgiYy76e7SPbBCc0
0UijIO987/fMiChgBwFhrxBqTp935PEctxvnnSHHpX+TIG8RbGzayPQsYV5AHehnn1r9Tui2w9x6
uWRYKbIhQ+N4TL9L9HHwlDTGgBesI/cqSomxGoStuTAz7WIx67KxtkQjlKoU9lyz9Cv1ub+/mhuq
cjnAiigpIR+HHHgM2b0YpPCaWjckT9MLBUvIeP6akcuKHR7kmUnIQmyvOGBngdBBoX6wz7XHyXg6
nuRbMMRHJd3lzXO3ebJrK1jX/XRbmRpSdFXkfIPoExfHGfg8s0m11qO+Zxszi8mCGIjtgGKphCDc
ZFjWWftHzkqhOknHr4srU8+Bg5xYdErMWRn3NKWo/BDLseKADKwmxY7a2JKQ7vFlgDSIsE6tclf8
Rtw2lnZtoeGqNKAPexSm4BnIvk/z+1Ktq5mn82dlgWBS+3K4mdwswg6Yy/a7iclbFb55tHEwp9l+
evbSwMFM4ufVbKXEOl29Xp7lwTfAogBRDiHRkJUMCNlee5uyiSO0k36C63ubj6XdT50C2LUSSr6U
E03bB0cXogSj9nEbEKvfS7MVt9EEP1/KLOPoYhBTwj219E6k7oDLBtHAsKCrmEz+FEZG3yQy5azc
/1yDxjnicTj6sji+ydoHwMzSeUcv/dk4vT4UoXtS2sYEe2ZDhnzTfJRn7jnQ9IQu0nHHcpYPDgwv
YQ4urhZvijPEqlxAzMTdNVUWUNheagGmiVJa+meH6xIk45UiWx4qM+fIQWyF+fAR5DwHtZxcHg4C
22Z2Ou/8A9J0YxW19nss3uwoOyPM+7SoK0CS7RLQZNiPV550YR/tMHXDvkF8Jv5fXpXgTkMBq7e1
Zciu2RCD+e5ju25SVeeD/zQMZKUl5RT2+lY4lRsdWgARaXe/xkRyH+0xBzFOaiz0aYsLhvH5ncGu
8fDOuox9usz8+12xgrYYE2Gi9kuWR75QQn0R33js8wnoFN0VTvx4u3hDYFRH8N2Z2VnTk+6Vql/0
XpagKGPE1kKcAjl5/MZuc8qs07xJt8RYn1p7go6sOPTD+PFjM9gXbJw/1K/t4mN7tn4g7ClzlKSo
6G7b1iMPLKD9MQa2KEfASOznhHZVJv0IYvsPyUyVBLXWf2zsQOYDnmd7ENWvOfESG8bnxiCUh/fV
KcIkw3rnhq2HKkeh1H9VziTrCY+N/7mRTNYFa3C7MwcHIeOA2huouM7DxpVBKWvphMbV1lZyYbs3
7I2RVhgDKVC7DvhbHTO2Hh70xHOyM99YQL7AGnG95oGbjncJanao8RvKRus5A6xZFOSI4vccUAYu
ANPCBuS1YGHCQh6goZBYmU27PlZ/r3S/xBT8vvkKwOORLNvjy35pbXrmdh8tSzXb6nKlfrFd5AFd
AiCj9bYuhbThXu/U4OnXVd5tbJRPTclPd9lzCcIaRklc8e43ttk/VAggenahn8/6aEQe9dRaDjXH
pB2Jqf6EE5LEb7Lv/f+q+l6ZJM+szsUWFm4ZwczdsgB+6R+TlmY3bez0O4Bu6J5Xc7jEluQiMsSJ
yob49ped5jsUDgZWGmzTeZZi2lzjnBztkLR36AzvE/UgsSBLkL9BT9I8fbi4PfuiR2Q2ngN+J/N3
aHZQ/5rDiBFceArPPhgfboZlUra11lkUtFi/r+plB0qrUYphic81I6WVrssYGwzZSF9Qukf27uOD
oNkK/9ljcf492CnBE6n8X2sJ/o1a6aZKRkoq4PlGqezGmLG0YQxnPxy+bDDXuxRkv2pNWXg/FO2D
bSZ62BMAvxzrHGF31eVyUN/1VEX/EIhO25blpojrTOkCH1pDXuYxqkOVingtgWJp6DMQQ5iaS7fU
7+kdTkkNlyi84sqj4EuLQYpbhhMwRohUKnQopSrEs+pCd7LJlG3HER9iVj4kJvmsLxoExPihaLXi
vh+kZ5nbD5hRk4Npb3A+bQwiQU7CAJKIKet5zr1496P+MjouF7kwvu4syZkO+aakX+Qw+BgvezAY
nmFAsE6ySkdCyPS1/LX6fd5eird1Mg74274MhgxQ1srAo7olOF8QPFcJwPcmsOT1d9d7IkTUNvLL
upQmt7z6TbVhB9f6FMbUbMXMPNQgrcYfbM4OBKN8vo993ZJQpXYtTMSun2NnlOo5Z4a1zSmn/H+l
1meZcc4HU5xzGEeEC+Zc3MkIsP5RTJASu36gyU04PMlAB8nvLS8LIpRzzg3SIJQh7pMZZSUnMLIB
dLgowuxChnGj+BsVTQiR5a+ouVHeibtOPHFGz32GUO/bPK9w44XUst30sQlFqFnTGlYoUiZvGmVK
6jxmjb/vedXGM1vHdp1IH0n5LFDG31Mif3eKK7lFrz3Ou8UMTaH3tflvGqLzYvmCt23uWGI1urV1
55SJ37iho5nnJRucDsJgY7N4F40v1dRyMfySrnx21GiMqbKtyLkWOY4P2SY3rb9AVTFNRv0WHQVh
M9blDHTbPwTApob1NPt14BHNohLQkImgKFoPV0gLCVfj6HJQUwpBnz4UtfR/jk57XVbR4R4cyrPU
TQXjdZa/v7SiqtAsGyYeONQCf+n+5zlARlnfDEMYYBeRClWbwkB2WAlMtzXZkNFKotnkKY7G8DUd
DO/ED5mIBAhxKfw1qMhFIjtrN3DBlcTLA12zdcKfZjk2Q/lDCv0gbwiX9L+gd6WKDrnAlNUgZzHF
cjkGs9wP+9o+IPw73dybznhU8DEF7Gr+hj8T56g5VmHe7I5Mi8IO2pZMbtomAv8AOi/s2CO/2VLI
XxlH9vbJYfJKn0EOjJmOHCEvGs7Cp03ljsc7xwP44XZZjpbL46si/rVRknecrsYd/v37zS0tiZSN
UhAqsKFaakc5SIqTUhe9f7C7ROhyjk/KrxdJG8n7ckpNrpWBxjA4V0nVNp1E3BiGrMzVMxZEoUm8
qm+obCt96P3WQVtRAzRBoGlIEDX9Y/nCwiWtE3/7YgF3DOpbaKt5UdlyIhHk3yU4wYoeNXXXc5B1
jBqXFjWwlqYkPDLOnRAKwXj32vsgBixmG9AbCKGYNO6h1AVCeO8OGL2YDen5PXN1ZekUGg0I7Zvp
+LCG/D4sRHSPLWay6XzPkjVqV2DvUH3kEbmgp3gIbfiby5dcN/HvLlo/H7qQiXtxe3Kwrr5VIzPg
A6vnnw8hSjEzVlBPoTf0gmGbIVbkMvRGTboVtG28LRTKZboJWM2LQ0AnuCMBTSAgqxpdP58CtBI0
EIq3u5QqO9hZMlX0I0UrPxbioqNYAMQ5GjJmMxOwRbIklQMdeQheWeAA0s9wmMiYPlESSnlZooi/
pSRAPRQGfEUtRr01JHLQJqErrW2x1nIaus9sFdoHu9kK00wTAv1w3f2RPfDj5s9KvP1eNR0kbJ0t
J+VnEupWIEHwSjrSrgLfciRK02+qtNDawBdCKIPrFAX/7z6Z+kSlkcNO6kDJDnkuvMqMTcAGvCp1
7D2G5Mp1o8tWDb9L1pquGXwS4bKhC68n+yWhS4qNCJ7tdiksj03I2LIPU2dwHa8TOSqtAsWb/Asn
KuAK8p+j8ZAFpRaoQZixisO0JAsEKvp/3iS34jFKizLoUN+zy4DukUTPs+C2YXNrGZy6jt+S7WDm
80tfi+HWK1BxC12i8ZbzFiQypbl6G5iEcHCxC6UxioYNvBLNUCaYM4Tqi0IYz9EevWnHb1llrnrM
dm37hQSb0qZNhpYyQ+Xvm7SOx/LGVEKhkI9LZYndnel0jSyRvSiQX0uivkEcmdKHWk/5MjmWL4Js
YvWxozRBQ9rmCX0ZXLhzN/ZHJ4h/wlasHHvD4J2ZqqULBMx8rJPcsWYTxN5ZTqZDMelOJVr4dVsX
BBuMDhDXOjR1JRvp1/A9/XI2gu4g7Gxj04bbfMAKPgb36+w23sN3KGLoZi+lh7ySod/02zVGlgXj
ersqw7gjRFmvE+kleDAaD8FMhpp/dKMpZBwxmQOpPkDA5I4Uv2eC0Hppl6uAYgIBuNwZVUkG1kdj
J7fwLprBFUJwzmEag7V7Ovrz0t4h8s8Y1sp2JkjKPK+JAs/90ksskKY1/dU1iiw+Z2j0wvAXD1Xk
w9OsuUvrd44fCskBepfbkZo9iFzhCaSO0+fJreSVnE8zAXecXs0U8b+WidHkB1RW03bI51eDhM/O
tHOPwf5GZzUvrXpQScWzutM14Rp+pv5slmJ9LKYghlYNpLKL0GRQY4ktdMacQ/NoNoMsgoi8vmgR
wtNdq9VSO+JSLZIit8CyVukv0amx3sGPLHllFh1Bji24WqSVaZ8hpNNP70MrB9mZPopnNrqAQrSs
izOrQ9W9PAHJ1sfmh9d+WjVB7+1AvO7+KaYT83FtR9hMW59iZvzwzxCQiWK4fsub5MNq6H86RwjM
be3+gVrtxp7nEpwf9sq+2ZuCU4BBGHVVEpqOavZRWRtn1CIQmXMVOp227sz7k/ZzJQhRqjngyKQ1
f/WGzicRtHBzbPMxaczvlQ2wbCBTTwis+WKcka3gsv/XPTi+NPDyaTq73IEn64qP2ZMYVCEAbi8W
diN4cYE3iomaXwnDzH17F04JLJisUA6fNwZTYEcXIwe8vhyiaCL8vpl6BGKcFEYRx9lbKMjMbctF
BdRjGv1JZE5dRxjv61xwQT6BQSCrTEp8kYGVHYqZkG8oUD2scs9tEyfzQSaK0DOdkWpNyHoa3SEs
ySG5PPloc9s3NT2xf/PBh+Bkpcpq1AmgA26BV7cynsq8riOkRg0d/ltUQsNPFdPw93Oo7Tom47Wg
6lXbXvFnfgI+AuB8MO1z4/6HVYG/J6ZjD+1FGExHf6x2gBDAwLUeiXKQfgbWJt558BF9bmub5xA4
5pA1AHjZj+f/5aCFp/klU8DWHkUt4nCFoBXO/lHNlaVm4WZAk7njMccUFk8SQcDeh4DTUeG1au64
WITEUQZPblB7uUwBtr/n4fL96JTc9WH0BUqggARWlOY7Qr2XC0mG54m37y8pAJym10hjvmPwoSDU
agpkzRDlVsBHTRku3w99+Hl5o3QYgLEw00bJ7kSV009oXBI2q4Y0pB2x5iEUtuteyfhFaFqdH08B
Yx9zRiepNDVEj1RPfAz8SIEHPxucBBTZX1Y4ev4nHkur+06y09je0KYGsI8oVhJTCGsppdkdFAhQ
bSCbeIKb3SIkGcuA/r4xt616Pib/RbmR/a6ke0vzv2XmNc/pj+5IV/T05OtXBX9pxpjxEqvMxwi1
vbLQ/ThTO15RbqGHHe+GcyfKxIN0bis6gitQhcxJ3soBCGosESj1PKG8Kf0M7zNQQBra5POYeMfS
yVLsRtxmmhkxnc+lrWo22XV317PxK+LaAWpClskUpmwWzPVM7V5sALj46WspKzNLXpIlMbC26Lgj
+zrehlqaYc6FussiT34MOuLuFO67d3LPHE4v07FIbvmQEgnz6ueWVzcN1OkCIL94qfcj5AWhEDzv
jx1cRhbyngYRkkrFPI2TsxW8XR8wNlRsMk0D0mHyP+opf3jxBSMYeNVRC//crSmzWqRwZSZDLakd
8MZrzygJNQ8vrYPaBYvc1zhSTHsgCsy8vZX1W38WhHjbeP7ti2UkCWhfN1PDViCfVblPA5y7tJl6
OeF9rJyQ2L5+NMhiER4/O4vYZOy+jMYjH09xd15qxDlPq2+BWd7Nz8wS9lX3fjY1iSEGfMqbw4Oq
Pw9hHLcWEpHo0E+iZ7uSQYUpNOTKFkUlfz9SPgpWOOR//xgzSReb4WFRXu53dZwHXLJwv5bSnyF6
NSBO70pXObXryx8RQyat10eGfI+04XJB6ONU2OMlGfvMSoRfTLRMjq2X+hA0x1yKHKLEQ9m7Qgkd
ikqe5p1qp2HhIMHrnY1vF4p6nZFaMo5rcv2eJRgdB2R3m7Zl4albEH+kdDk+l+sPSDcmg1lnUdcM
OIuemFkpd0Zl3BQ5wVVg502yoAOHbl/IdrlDGtyxE9vrFkvzggK2JYq5YEtnkfEmJqQcVcSW2dS7
f1dYZeamhnwQs+i1qE7m/6OvN3I8aaJYzJ8gU//uSQORmU5Mjg0rN6+MaSK1Cgaf21hSlTvBoRTt
FuLFmuiDZe9Qh8D1hu0XlH/ZO5DKxicCInZD1F3F2eyUgceeSI/2zt2zX29W0YBsK49XRdCZKw72
fbH3LdB7E+Dugd9BKREXORl1FarF4sxb4Yl4szaUENAAmAsDizPH7MSMopMj3vrYs6axroBlpRmD
vSyM4VzlkKF4puN5MNAf8DWgx3uIYFRRAw4eEkBMdbsD0ABhB3WENNH3LVwMa2vBWV4/PuUyMO3T
xPgHxzfFzMeKd5rdOwLjbAVaxhKqrpqj2aZ/XpytTDjRA8SJ6cCHG0Tmq8Mi44ENN9w9aaSsUmyJ
YWdNow8iDPuvpPAx0lnBEnodipjxyIb1wDoF8BlfB6GMM/Ys4eiDmS+5ZYRMNRX9ZZsqJ3CrhA4W
q5Y1nSvIs40NSNpS3UhNLZ4Z4z/cuZXpWYKzmj9AYnCb4mL5VXNu/qYJ8eaETPeie7eCI4Hs85mW
8KSeZriBJRlQpC7OS/nQrF+hX1JHc6gz4VMgnSRHjon7VufF0lA2DK3VICah4/52mhdtGNGtYVfx
zs+0CWgIRd2tcWn57erA2XWmLxZKSDwIjlFQPpC9kAmFJjCK6ojEOPj1dthOOX/DaTgvjmajwXj0
8auQOC4ax2/7PuayQVgSB3uAhzWOx5bJWjuyZ9sQqAUyk+ZuSymjneYHFZHKvcg3b653Cnioq6u+
dF9JYzWKN6rHC3om0Eg8TMMJZhUBQ1Dj1fEvO0oLXqwKpOgJBIWY0bpEgd6cnna4XIvAG3t2OV1S
djuGqMGbJ+eRyS6jAbTvkeA2j3WRkXuNXOTgCCMwyz8TIhgaizyNnDUxVd+fIgdKH1gys3rFAgXC
08KM4G/uCPSUtyCJvaVVVu/kLNgnPYno/8xNSaADE7kMQF+I/2jMszjlqjNryHukdtiOV2//v2/4
3H+9luldrP9w7k7bV+kFGJaL0dDT3lq9IP+iJ5Hwfy79M4tDOnZooh9oQm/jSxB41BQGDkn8dU03
KTBkqRt+2QB4mT7dT7YcrWrgzZnxNSKB7HV3VVapmXVJabE3nrRwpcEPE0KjWjk/WLtwtZxIS8Sv
vmDgMWC410d0ehl7043jXR639Ip5IAbhxROThQ4JG9BkO/q7jsMnCYa+tDJyZACMnAdso0GSeGNh
BPupsj9tfHxyBoUTqXxaeqXsz97tFOm1Ou5fhUjASrqNm5q3VRlZUlpYQqlHejXtajaaxqOHx8sX
EeZHq44pTcmexCB2mbxUtyn083qXg1kiDGcrcWPhSPSE4vMwMqcTZe1zpRxqM3k/5BJxmGYQ5vnc
ZXff6jBZBVrcFFW31mZgWL7jCoEV2tp5UHlyzJeElst91F7IxQWe/5K3LnEGz8luN0Z5Yp0iE8vr
KwVScaIsU4NGvO24iun6yT3LNKISpx4fHfo5+zlAZQLq/MvmYBTp0MBHOKrEYEmVFKwqUOIUImty
HgbkCuZIfkSdu8vtpva3sQ8KlURnSt0l/yN0j3+D163nAGLQRdoAy5vAARiKE7yjWWTdLD9Wssts
3ISRuMknByARS+Xq8qYf+D5RKmX+nveO3nOW/dt8b7BnW6vjAyz8Yu9LYX5CLBZmEH5njinXDuKS
kR3ovuIMKr3lGHi5ClKS8z23tvaCNt+WM+n5WUUIN/ifLZ1LzrasqcRxOGnhLYtGTzKJVDiDwkRY
GnZ4amD0kIUDsXXQUatsHQUcbSpM60xWu0L1dqxFoO5jWzE5zzVCpuMoGcsb+/oJ+gQNU5KT/XPu
AZpYLmilcWUf0GA03VrR3yo83960rgdldyItjBZKRe06vJ1u1rCV3a779PR6RlNocgNv8+e8bHE6
sRAzNTyjgDFDkTdkZ5q5p0wclywf55A5Jb1EkDrxXEQFUP13HZr01CbZNyYnzzAIrH4BoCjRaMsD
WctVNNqrxSQwtC4jJzthVpTOGbh9xeniR//W/0nK56sRwS6HnjVKxqHgvHpEfwjByJl9xxFHiJGB
zTYCPN/fcjsifQcFajt7s4Gu7QntV/EN8Fc52F5Qov+G8os//89yrLXPBqe7+aBjT1+Wb2cMI5fz
Wyv33hewTtOU1Jkke1DPiWQQCqR6FveuhcmvnZotMGpoWfILUmTkDVRqzER2rZtY+UqtJHdeIK7k
Aws5NHrobfCdv9htfKoB4//W8Tg2wd6H5gvt3HQcZPdecaod1tuAO67jkdxSmuJSZKZMxrVHYb5z
4xKVV7jm74QMC8jJU+c1BRaCRTMhWimO5ZlLieKYEvUTC/j/riHbh66Kf36D3191JNtIEz9uZBXD
tBHIZHPwVMytXg8C2hhKcJmU/l+6Q+YaWPtWhw8/I7X3TZbpBMXebReVlfpTRVmqUYS99YNcsTZB
K50cttHCMbWgYkizqTI+DT7HG8zl0LslZLmzAUIWFil7U5klLXzSfSuGrnnMMzQidezZ4fl5iDJ4
ZEt4m8opaNAzhHyc+3uZCaTrqNg2lpvN4TTCHXygtXHqxF3hTgSDNqly/D9Vw4ip0WN1xqXqmpnQ
TwXhwCBboSjyGg1ptojnzrN64bZoe/iu6ND6Rid9B96M1Y7KdRvSJoKl8F0gna7Dlgx/r4VMH/f1
qnRiCAOa4mgdnPYbMhXFZJ3mJUyQ5MA4C/kDRQY8quBJiOiOkueH7CexyZ8Dqng92z7dQ2Jp+lDe
VKBwCfJPleKZdMQ7BE7NhyfF2AIlRWbnMDj1a/BNWKnzTE5lPflfRoFAyEI0Ol8mpmjdALJsCMqR
s8fMEORus0Glh6d4450Xa9KBtyKKTIdT/4PFl4jqdzpri/uDhLep32SO6a0hMcuwgtNXJ8tWvUnk
zuSc/7OaYDhAZ6AtPw0ybw2JUYO97e3pXpkNdgdOiyiGBvHxbigO8kmFWyMP8BFj4TZQj3ThH2Yx
QGkkkpVKeEyF0i1wiu15s39ywey0ZVWRWF+pEiohyfyzlIBIdWjPIVtvfpUN0eEM1IuLPJyCpNYy
VZmjzdUOWcV5tSZgb+fBgWsZdHt7nCnNwZdgDTLFjFpCKttfkOQ4MW+6jCdeAzl2L88HSoybrvWA
CZKUNMdDH1ssPA6Asx8cqJwRFKitKajt5wnGw0k+hhuTQZuqnlXRbr67AC0eqhVck0Sw5CgP8AVE
1rdEvv8GSB9hTvBEBN6jZJyagPnEqKqOjLLbJPOBkg/kZ208PvYFPELqtnqSQXfxya9L8iTn5Mw1
7YJTLcbh1DT2C5JGoaHiK6iGSnux7SrlWfbbGQMX3OtniPKb7al/NcXcnJN2dz+1radRU8PEpZrn
dyPj+shM3ajKSVSvljgh5FIQiWFa1evfZbTm6M05HY707WDOx/7Qv1yiYGtM+hDQ5nkGKSSrk5vS
9Wl/2ujUF5y8ZpEP5T9ty5Zlh7oOlOWZgMEkKIXEnEzNaXncv9ZEVfTqFH6hhTrVTMgKSHzD3aQY
m3LrwwNwWHT1tZakGqIAveP5w+O8rtHzi34x3C6fxenzFES7lm6peRD+D4e48DRNmKTzqEhmVd4l
nDxV8iKwqRi2HFOhQguZI09ajw4lBEuAe/Z6GCH6CCEVVFxJkc3pQsQpvNwyy+S0ORctqMM45WF6
/4614ZGc56IDR3RGV+O31tUcOTkFq+QrCHcqiIDV9qOY16YgonjxC5kwMZh+0AoVwdF55uUC1iPR
vYxiF8JURT2Pfeq+QGX7OSbkhfunJuCUxclAAdxxgikcX9krHTu70YNgceHACW6CyVGbJFzcwyVs
Ponm2CpuGHla8BgkXOAMEg/soU5mZpVP84BsYA5WbZExXS5Bxf2kJ7XfoMGn/le+m3yK0ev0d5Pw
vOjTV+7RiKWmJynJPyBBMJ9dbAH/1S8IIgnRtt6HTGos+ekBN1uXLf96/owZnU5TS9OVuWZp3uuc
dJCdW0gRP3QE/URkFF8UDN2h4Ujy7PjrX8vIo2J7QqTERdfegDifB/SsW1bWV/Z+g6F2Cncjslaq
FSuBYiVeAPcFuqENdW8iQchU8VQXp0LRB3fazQL/llt4p/frVxdezGMDDRNpNhAtYy8gWAp7KhOT
667jZAE6eKINJSX3XvCYdIvSGCx6buxf3jCO4wU//yUQ8M7+Czm+j8rWTZt63ORROLowOla0suh9
vPAuq6Qek2UP2JrqTSsCbEHw8529A0ZoOu6als/04PV9HxHyYfgv3IQ/KdJfZAJ5gMBfdQgDmRbF
AV+C42TYbptMAUZwcejc5BUGnbT8uvdSuxmzU4dxOldHPv1/JBU1Rw88W6gjQNHXMC3PU79VmcWa
PvX4FZ2/8EnWs48MLsgwqdGuNARMNd+vtesYVJFSh4iTUJrc1cy1nVIyXbJCxAh/j6tQjNaFJxV+
Vd7RB6aJme9m7H/85KHeXp54vAmvwuMg74+kndn3vCgeArkVsH+jISi6mlf0ozAlghbZB0D8+AqJ
d7Hy1x8LkhGtFAegqQNdVTlg6yziT2rj0tY64e4HlqkxcSFsZdIyO24F8+Bw7wTxorwEl9ZEZjFk
glRHJSFcrrze8qm07c7HDZwRZqvRZHUKOpKz41NZWb1Binlt4TUOkzHyVxBxaurXrNg8TAGGT1Ud
PhxYxKb0ueNdm0oZz+dn9b3kho8YRr5bLBNbr/OYuK2xD3EviLUJKJREP9aWnjCHoLDO6h0b49Fk
rU1ZTXkko0IaAk91hzflvXvyiW9ac27y83coO0q90yTQqrzTGnexuJrD7L+b0aURvhOnRbU9wTUA
P1c8WO9Ov0CEf0DLUem3FKhcJj2OPHXswKQl3ZOEwwWAPKPr1mfAyRmZ56jFgJmv46w99qaF+iIi
DTToCuxJIIaFJG4VWzI7cy2AinCUjjeCdWRNrJA7lfNsnOzJuqJ2k8PJyrDYuQYGxL0lSxf1rxqZ
4mWRxP3qviiAHNmpIhF1poxaq77r6CNlk1VT2Iw9/KTiL1QzF9dO19xiL9o5Hvvp7X/Uq6kocAb+
gJRq2ubWFMVJP2Ra506jlP8lNS2d8Cdv0Y5T0L98D3EW5k0tbUSClQ6rQqLNWWBAu/nVFRvNwRCz
u4jN4+4LIIgaLnfnBYsIgzbg8hITx2iptGl4xd9+pRqRxBgW1s+oFpN1wKrsmEpUdyKSp3M8hoQr
/+T7CSth/RQ3sOm37BgdcOO8cAcbqdxZ7J1tE7mayMi7AMdex0RCjJ+FBplm0tYcOlnOxOkCfpdy
IeVnHohO6e1XXuMJXWNjdSJPFob80f6f9Mfd9IGjPpWremt9jV9dL5FPfQcdm00vQHi6DtRbIbSU
hIFpgngLkYjoHM8/rqp4v48hkASyu7PKFNjlmE6BNOqFtIk7UUmbwLU47tUtGsCWB75RQk7upIKr
00tQN4jN9BNjKOMyM+tZbLwJy5BVytR5MWR0q2lPjuCOMGVq3Kudkethk9GouHFUPJH+RB9glneF
dbTkS85wOetdIR8/DRblHrK5NXW3FGdBire0UKHIXeXIkNslsfHWLMzCwrTbOWUYgcPtxULc5MnL
ElagDllJj+NeEHOTb0TOgdjKds6yvqNh0eBhYuwzWKJ4dd/gvUzV0HondeimS0d6Kb8gDmwIk6U6
2TVWpsqPJCWRxb1oECmOFPqmHysoFIZ8LIbgORwflNLxRuUk5tvFzMJIie4e6x6O+0RsqPtZVeLU
4/9i4OIOYzeNLhgnsEkenf/6iOkpq7tAXkU7XAPNCAyZyOqiwJgn6Ko44oubn1Kq7spxk8R5XPvf
N+bllzZHcJiCpp8vZBv53C++uZupRXRAH2tCz0jMG/RHrwXML2FdTiVkeMeu8IwYQqzDKpPmJBHt
FRs6vsizWTLi0ooPGw1cwP32+Jr7iVT+BlHubhdhFZdsVGBQGbT+UjyspO/opQWKNNvvId2pJw1u
s20ih45gWWBNJtLboaOXFIXN8M71RSq84J8gmwjtiNXZzCofCO2X5cWEJ9ThrVa3+jXRZJie/fw2
0XCnmxlmCXwjSY2jqta0dSZWi7MWAa5uu34zd1pTe1e6RMMn5l1Jr277EDhzwk5jWCGezZjPb0Y8
WBZ9ywhCn9OFIsBT9lDHEct3lUddLuYE3TA/nX5aGaTi8oADbs7brPisl0LD6Wml4dEWvt6cyrX3
d804zm6/3ekNixS6l4vj9eZvhiwkpVp1cDJOXOEIX2Hq9SQB3xKn/NWLOfK+OnTSZ9rT90WZJ6Nr
Y4Gp4zKSZd1/0afvYH9pK4FXbycFK/vnmmtm3zqrB1sqQxw6YAo/64mKlmadXWliVA2IkFyK8PYF
1d6a/YILxRKSEzgMD2TsHlk2dpRoeOpZRRYmYjapBHgXMjGgS6jN93W0hZqKLWmwwG40Yqh5eWlu
IbjJ8S/Y7KhGJArSwvOVKf/GALLsz0o8xoZSmwEz5eatvCQa10nNqkd6cs5uPkxHtjrEUk5oLHcE
M+W+Rn8BRC1ewW37RqFTZBqtTd60VlKjHGTqtFCbnwMQJUJzdw4QPrkGyKJt1ckm5rIW9pELu5d9
7jvPxHG2AdsZ+GxguJ/YU+eaEvjFWyiPuxPDQ5IFxdwgXUBQxb+ApcCQ0UHMnn+FeA/r5dro+8DI
qs5JyPTCgeaXh74aEJ9GGy8647o8VPdo+PxnxYFo0kg0WHy/Inp0/aXoH9WQbC9teMRccK/LStkB
SycC28MXyfjnXoeynKbaZbEshqRh4lUabQq3FofZRs1o5+lHJ1UdJ8tPQHdyrVWbnZMjMpehSLM8
eAg5IunIH2oRfvUmvMEkc++4YYZtDqMPPQe/xKhEtHEnlQid9cSXDMHPZi9TJOaLCNwlYvyXA4HV
Ohri2IxnM+U+7OcIUJ4lwo5nHGPQxxIJPJKoh79vlZ3KA0AxCVvr11Yi2IapD2dPfGJpg2Ik64FG
HdfE0OtI6YBzNJIydPAkL+XY1AODHWQWFtBlw51o1y5cjHPWGJ5Rv9xWxSoqwXiFYAa+Jw01Sfyo
BkvGo5/JdZZP4LMLX6MWftR+VErSORyks1l/tDSOlvoiZp0AImHLn+jwD1KtN+69oq2gfJ56IpPQ
XBfxhIgAJJReZPAvFci1g//NSmPmOjgx4xtAneHnzIfd6lUqp2yeAS0ChNJ6/RuVMLeRqfNrVi6B
8SzqYRSEE93qVooTTxS8YHthPJv8dXI2RG9b54o+QPFMjBmDdKtIcgFDFxVUBjIAYxOOZdN5SqqD
wne6A8gUh0FPeZNHIC9ls6NC/mL5WFavvsh+4WgerxdemLVwZVa2jFfCLYw1UmXEL8D22BXmju2R
iz/giZHLIm9px69QVybVwD4wh681tJvais4VOlD4RiwnSnMmQR2xxAvCl51egbr0Bhy/4TPx+Ylb
ee3VKfSarbx9R4CRzs5ZXnzR8qZ8d8BYgaaw4ihejNQvBAyCDK5IPzF+5+gILauTYX+Ktzd1k7UY
gAg4l8RNyaHU2gVnu3mfxdXBI6gamy2it36gvn1ugRlA9dXNBPNiyMc5i+WjJmJCrrjR5GL7zDHS
AAzebDBhnrXv8AlJdVW8MHZCjKmSG2yYa5xbmiDGPnvL8AdwUwA6Z0UZtFbuUxNdGOVRtRoOKhEL
n4uHIa2dJbzu1uhYk1QEWouKuBErMu6iQN9M3oNPxHKRWHLvV86YCrdoY6JC55y5CJoQJp/d9zPr
hZaeA8Is+a/Z+jQaYXxdfoehOe8CtM4OieIFzyxDeQlFJHWJjNT379Y5c74Zpfi3Ye0XwilIbotq
IOh++vX+sqwU4eJ+bs8fLFaHqbeuKR1cWtdJ9T7tpl5cCsv69G4dRKtvfVfBD9x2f6dnfnKgo6qD
W1kR+FzVbD1Cz1PVQTfKVaceXpHu/vS1T8g1gFU5BDoTdzy5sWUXJl3O2LsgeKUG4+nxP695mLVn
0nxqqwZ6R8phjniX2+H3AuOdmTQEZM5MTx3hoPhkmIVC71PgZLBEjJMhkpYXvghM4cu6WkxwQPwS
cPT4TTeb0ShGskgzEBy+KoV9Bdgr5n9VCIxvq+gu6gw2C1YjFKLEiawSMjW2IpFe/CYxBiM2V/jg
cy5rm46bGtq7ShSe/m8csmnSR/TRHQpYjYkTrzPODYmePtrdVG2UuDL/BOX1UO5J7LFII33C0h2a
EBbFsyS2NkzxNeAzpVa8wgJSxHJ+lCqAOXnmtowxigzD0PLz5zuYbN4QA8cC2VckdUkFszSd1iCN
pE+tiWs4WVtzMMYX0OhrdN62E9Ik8fLA/AM/2BFKi6mjZ3GlqckCgsmzXkprietOPL0Fzsl3Q6t+
vQnZ89iE4cgKLGZBGEnU8LKXOqRPvO6/B6uZvoJPS9mYAeafnQUYS2ZjyXa/KOrMDk+nt9SQd6Fl
rewR6+LOAw/lyj0gsRmTv5PqFCI7BcgcBKIGGGiYhlEk6cXmJAiE1IknsIdL9Ui7BJqpkNBg8cgy
F5nG3hDkr1cC6+0RVcgn0DutNQoe6qMJ6f0ZHbvalT/VkKur8mp6xASwzKw8u8JOQ+0+mu3xPT3w
xGnl9jn5NbVZe56PG2kyCWGjZxvZovbiiuuc+RwGuvtpJ1RoUfgJhU10r1CYw1XOreVuIif39qDE
NR2g31PmOBbHWsgL6yGRlmqbv2b14kwP27iRc7ZSZ8uSr06+5K1dI8TRbDvSMoUhkAKUpbar17HV
atfHBFnI8CohQHuuwr19Z09sbjsqaYjVPOEudYtARHwU1DGdjDYnqPPSGaY5f/WfDJLsV95GIo4z
YNjpzLOaYXjB5J8tV7ywrFGxvtPuQkeRDk70pyNNU1pJuIHF0nKxsBvSTijyQtzKdxB4xGVOmBxv
uif0C8n7a+3QJhK0Zrpnn2DSR9CQe2WXDm9J8F7LMu2Id/xxpTEQfbbGegPQJHSEZ8GmypWqQFTd
0aohcVDgy7I77enxw8/opOnhu/bbosKaYWSzcaOucEX0LcWKNW7GpSzrqJivWGop7O3KuQ9XyqCt
KYBocRgudyW3qcVB96UixXD5PKtG0ji9QcWr9RTl5/3hPXVay+zLgFMs4ckZquHessnk8LzYGcNV
88bdnGk7QI/N4glXPanePcmT+eD8XLiMCxg8uQkMxreaYH5NV0SHzkD0bO0iDi/C/yityZjROZp6
Sv5bG4r7BsTVGNTIcM5xzbLt6MOCR8wYFJw7WGP2HPnFaG87wV1BwFQ2m4xGa4LpMNdt7q9UFpHc
YuhXf0NrR/mlV0dmrpULFrahrmEbvPY9FyWJPIlZifoswO4hOcbCgK+DWmMWetJ9SyR7IWNgSXVg
31r5otStHo0aNZiMPwjmtsW8Hd2cRRzXsvBXj0zdaExl/A59J3Fbe/PbdKqqUGEdmNtAgbBxT66b
iHy18SRd/B8ME4BmGshiaNKWR7jkQq0eZeRr/Th/BMZRMEJhbsoTmSWsEhJfcgW4HMYZlSpLQwXO
RrS4XKaiYYfFavFVSu+w24jyzLlCD4kvZFI1xArbOtm6oyWaS0jUqHmy5eNJakSfod2nQ6pVDkT4
cWcIY372UADWi/ZdWyOulQqeTptZzh6pmWGB2fiG5h1xan2qC8iqo5nSP42X/b+ea0jGa9I8jPij
czSjF6RSG00LaqM8JsikLwxlfVx9e9TU+JHx8hCm4K/36dCacbcMlrzVwiZZObmxuAmP6p3e1AR5
hgVclW4MlS8v3Zv/ULNq9OHIaxbGVHcXNoYByRVbv37MCzDOOlU9bhA7lzpseevY3QQw6bdoe90h
e/V4UoXGWyhVyOZrEaz65nFRKbYZ8XyR9t4lh21wQI7pYSb0UgwM3MtwmMEoG4bRIAVgGRckISoM
R2RU/b8l2xe8ygxqSCWLXeF6UROJE4YoYbR8ZeE7yGbGfxzomtyLrRtCchP4moe3o/rzR5WjCzJB
Hhn8BH62oa9nVIQ7ILG+IPSM1PNvqxQN8EwrUKAAdZCvUFYywMESDEhl/ox84mul1YXGP6xdrXp1
so43RTsLcWCtTys/4YYUmbIB6regKI1I12+l7197es+XfF5buHXgflXmY9yGZigPhU9rSUCgqx89
lCQlDvQKuhODqeRd+kW7GVG1S6LhdWtreE3sM9nYFP2y4CiT2ZCKR0unt+uCTertao8xCl1G8yXK
cmX/zuPQNFz517IYtr7XK//iRcNIdYYCKiktue+pGEKCpLvqtvuLDl/nErcA6Q3Pn7mk9cmupWjg
wuiAwRQs+oi+0639rmK7rmrNlWjSx7No4aslmcqYJT5r1IyK+Nq/pT9KOVyaWm2EsXROAchmCSo0
H371cO28nVXknqn8ng+lBJQLL9o81tVR2f2WiuCVaRYGoxqhYccAuwbYssKhfch+8BpX4LzjAGpK
YcJHMdDM1v/BOdr7FmUU/Yz/6si+bI8mIT32GLTzuTUf+9uNQXl/5+u5sU2M19lAojvwUKXTqKMj
2QiTu6IANmq07dRDs+8o5arcwTeySaL99Q8d3Kz7kIeFjDvdeiK5PrbogO2xQaTMqfbkGloka5O4
sVLIXV6GA8W7AzL3OlwzY3jDPIJ3IEJ8YkbwLVq/Rp44gtr/aA2mPCIk/wK/sws4bqDfDVlP/QjT
zQKb+w+nd3egXMeJQrbbBp7YoKvU7xmAbAx7VtzTWvrjYN/jxdtbB5FxnJ/LFzTl8lLwdw7p+/T8
20A30VfAi9yYjPXk6Rk+VRtvHD4RIeyuBlXn7rOv6zuxiTR/LcvgZoIlmoUyyU85N0PMl6Mu+aIX
rsHpXhzzAdgk2DkkiALn/kpff4Hbwq4c6YKnPKTvbG6oJ/BUYmqYHyrJcjfOeUguwEDq/Zszr79H
nKnUqJE60lehasiDfL8q/Jc8Yrp/XkyVgCMi7TKNNgVamzpR+SkAchZedV4I7ASUE9G8TYdKSc3m
vF4kP/iRHcs7SUuM3J2Rcw0+Xs7u9RiQg+lZPzblK75RkTQ9IntJ2G4h32ijw2dJRWz2bpZdrU6s
YGvVR9xpMw2lMyNlVz5cULQIojdwqLKIF/+l9PcfGNSLT8wFG5NkgT6zAU3fu3xSQLjS046di907
kvl+nu7tYsba7Sl4TRCPIlWFrvlmsIjVOTFAacIw9qXK0pAtUH+r+oprZ7b9JuS9ZkhUpm23ksmh
ChUpuP7gvpHgn0rgzfk3PH6iyiuHlsyWskKHeX5ldwuDjaYbzIFkruWgKAtqTJQutUryP2JYnYet
v0rfF9V2lPZCaiT1k5SIS9rckSULtKQa7HTkzPV+2nk8i12EwfiKMkTNPn3xAA/fiWWW4t+Oy8Xp
i/M2xonALpt8AE5tVQeUTot/5oXDqrk8s6WorlmdLwmUMPWGxOUcF1+6yFIFgLbF2GA4uILYuryH
bGp1khalD0Cr4IqTN3rZXme11YJ0H+jQ/sgaD62VHWlV7ov7FrpQmBPllbkijTak6pcw4cxeCjw6
B5y0qTbLOpZ0jp7407igQ4YHj2rHElOG0Yhc/1+FrZ8uBZxfyZw0vPZWQfFUOWycPDDEp9pa+KDB
cUzbzE2N10PB4eA0iHp0IyCk7cZT++nmQkZF2qz2wVdwinCHsbqPT4jmW/DISQgxZM8Tz1Ke+TSk
skGIsd09GFJusHEjoVFcllUkxFR3Bw/fg9mL28EvPwRhmxGc7pL1JanOAD8giiaHUGfphOPjaN0W
v2EDyFsDgqyFHkWp6BFTNs77lCincRPvW9+SZnUUO103ju7w2Tmu95HgGYH0GDrdgybv5cNfjZas
6tJTW4NPrqVDeC6rue60H11koPBnTc3bLgOQ1AirRNLDy0SW07lc0LGH7Ub1FphZzhNo+Mow9tEt
QbmdnAAPX2oDJT91sguTA9v287Qdz3xP06/zj9Uqclbpf/P4WXBkZxtYzWizryEautQk8fPL6vvI
Up3ff1x/KLqGZOyJ+Ebm9Wj0cBcl2HSh0EAH1tSBGjM7AqALQueOh4N4zEX9Ocp+gbjcTSs2cLtT
9twV0LSZwcK6xB5Au/UXfq8BvFQ8GKdBFCfjoQJv1Bg6jBNDi2ux8TWuExigcNCHl34Bq8613Vu2
lvLlvuza43dmlS1CgMQ4ihvHTZIvkm9+xMJhd2exMM0rBsymw7ipsWU1dRLhoYDgd6DhvZiqY0FD
mUaAMZG/H5PiZc02fFWeyJvm+x5OO5eUA+jT2xKcA3gF1FO/e6LKOR1mBG5sgioZycTh/ASnzZes
l20VPEyIZDbigSewOcIR5680aXIfe2rENGpxOEefyOWxxGxOztgtjm8uSxOUQius4zVzTweBz4V7
GeMu6BDJUwutRDzWbep10W1WQ40gRCIQ4z36T8beUhNJN139a9sT+loVCrFSEeQ0K8IMMExYn8Al
M3tGv239N012eqDSedcF6qzCJ5DxnTsdYNJOlB8yN3Fvf1GM4v7c2bMTlebPRo/MZqyLPCFVasOw
hbpvRqPKojcAx8kk5+nPPVHCLEvG9NtyZPx+dSGbUxBwmoCymdNOuqgrZy0zg6qbWi2W9AGok086
zzT8t7uvzGLckRFNvVz/EvpB2fWy0bu88IsSVOdk6IfYky871+5QblSOz8+IQdkv2gB4zI+Z9sv7
h3bsbeaxpbd1HwPjqG+PO+FjECzK2+hq7ouM3mRjsvdrF37Vhbomg9QtUboVrhlBkFV2+RNbTOOw
Is7BmAxhVdEkhmlImoANuKRj1LxaTFY3wLRP7zovpxa95SCLq76GhBOK+ihJNIDDCZP9FyrWhWOS
8lSq1d22pYLIWLFh1yNTA59U9gs8+50BkxBbrr9rmp6bLnTzOLGOLZSC532x5/IzWj9ibsx/He+D
sxaXA6KTOyWAArxVSkv44DvFujuierdl/rWGiF7RP2+KdxYi7V9ShPved2uEtziT5j9PzYQwaP54
aVaBtTV4vTY4gPX8Q0atCqtlvffnk17iBxgusc4DFotFqRcKoTc3syExyMSDABePi+utwQW3prcr
r5URBF2EGYE6/lYtrnghXZJTQQEYa4RrueL/ocW2NfgWLdBIu3louzFigstyPqjDJB1HAHHEsnvT
RZGhmnErIcYLrdS8PNkpBt9EqZPNDyhj6tydje5BQWoIKANsKbVb/HT0tlmNjCO+ic3ljnG4Y1DH
5ZPGn2yaEaaN6SEAjrHRfNzBK8qFqnnJqDomiPQz9yVQHLnIKkpaWP4SS16sk9nlgDF3Sliap6IK
ivwDOmX4GNAfT9P1u7G7p4+H5mCqgfejeZywbwl+nIV/ZPkVOMiwMBCT2JG4eNsmIufUIQtfq4Du
81daWnqzA/4zwl15h5bQzKzy1zKR1hEBiaRVgH1bTJrSQk0m6Ws4IpwJZRj/VE9qfHnK/MH9xs0I
m/E3z8Qh7PCwRAEQkdr4HtF36uz6qeNCmqCubz5sukfEWf37YEctX8OjV8K7jVSzEkD6pIdDgSVH
WqI8dCZhToJCaop0yZ4dhphxSL1tATEtjHt32jeBKUrhf9OpQXCsEiLCxe/VKd2fHtxU8kYwv4zd
Kf9gcC5kKh5E9aoSxRG6JntgDbAPCfH8v+XRg9XanCRAQ49ZVdHg/LLsh8WKeUMwYg8Wcp1tFNKC
oy0JLiY2H3w+FkRkkdAhcihWWx4O8nPjzyw/oy49L5kXzcuDhkyxYVHdiuNOUoUGHCU47jU62BRx
Rkbfs87IvnLamsgU5tMv0OvjUJ5EnogwdhZHfJh71qLXA2WqQUvwNfJ/+AAHszO8CJ1P1uAPJZyK
BJnp9o5bY15dYAXpdbx2hml595Jtjzjeepwk6uZYfdPKn2oUpmg/NfmCMkdvFzZLOzrSTP+hlaZ5
HWN5s2A74BnKWtPwTg/ZPlVuxOO77mYwdapWFZ1+SDGTU7Z29heL0OTPjZZbnbT3YlrUqxa0pHop
1hAqfP+ejJGxJ2JUaLnG7vk3OTGv8HzP1YvPeKjHhAYxaKxssjH5wzyxChhj2p2CQFLHBHEWA4BP
10gbqSqkuIHKc4tn26EGqpbTxpoF6QK7DBFYsVahYRnRF0/VBv3lCW3PWtQgbMRpMxM/HuPPO0uA
3ihaNL5OCWq3XGnh7dNPgEwjI8QBHWmf8SSWi5PXoZuDQPIwgvuvPbKWo/hp1KPJMf7XIPNPmaPX
qybPdEERoLWJ+XWDLjwRS//lSA9QolUZIw2efTALj90pxlFO8Ji9jhZtGJtkDkDDmH7wd+9n3buG
MgqguoSyx7TQ5GwWSOuRKyqeelw5O55IXqe9nJmd8mkFKoG/XtHQO/TrfLhlWrjt+UfpvMiNYADl
5xmPcEmtrMMJkAC7vFtmSfqfXbh4sL3Bn7iiAbozYe3GED8fFZzbOWvh+4BC5xLDcpboXbftJTtK
0CyKttDZLjINHisb6sBceqLvN8kIkqLYQUR21UxQFMuicqInCofHJLOOAH709sF5bii556/mK+Gv
vFX0w4+bduJFHiLox8Ar3GXorZ7lnJoCpjDoD24VLcnU1oPYrptuDm7EV9dqSsWlNrJD8JatkVez
XoaitrULoYuLAoF44ECOvun1eYhiU1Apfx+HJ0dpNzfTVwFP+fe1XiF899CCi0ZbKJDJVvoYgNQc
G4kxOWLnB8OIWH+u4YEk2yD3JfV3/5jh3DozP8m2EzWa8XwaS3ax4qWZHBtxEEY+0hXakj+y2XUC
NRwFR8emsMcYuebuhLaDEerzRffbu5PeYUrOXap12V4mofsdEmB5XqWRSGEbVhXmhB70uM+29ewE
b7Wh8kW6mHPcLMFsvehi/Rw0gk7EliYjhrzZTQSOt1GLkWBsvHBYBSD5U6xFw3D4xRVjq8rE2ek7
5WjFcOubmA7AupBI1RMTG1XWusC/2/vxE2i6tsTKRu3UiK3wJm0W0Ag9/rlI78VnRCqpgPbpTYav
43obMYDQH3EkqVI9cdXY/xdBEnY1CbcI2CZ2SyPgLDIyx4FYc96RkKsopKkP9CGfU9a4EMisZv50
L1fY/b0CXDZlcI1OAbGd+RhcjooUfuHZCmmfib/6GvoaCqKDIBffV6HVwnt6KQsV1zHBMyECt6CU
Ul7a2G8NiC+8NTLNOY1ffWZOviNLcZuIRXnXe1UoEwpRNx+6rvF6gIWbjIUMtBfaTvghjPAZmZMT
WZlNDjBPGvASdr8nsx4jqF/+cAwZndmQutHo0UG4/tZcXsGAKzJaxQvR34QyP5Qr83UFektgVkDC
bLe6APpTb06EpOpaAxLBQAOrEoUOlZ8xh+Un9QstvLQ8LeOsK01v441JmgSlLnHLk4vBAloinY0z
aAn0uyGlUWXvQJjYS3xCo2N3nYxd+edOFyuA/ugDNC0fonJkwxmli9QOR11WFqkQ8epU7fQlvWgJ
zmTulYSnsidicWHg2M3yoNz1HDKv7m8FzWvGbmJTyzGGXJkveO+DRSrFnQS4JXsPGdSTwVyElEwl
zRhp5KVBPgylV9jZg8yN33TnPSDtrUwa1F4LuUfytPptwB3bhoAbV5XjYTWIvImPb+duypk6wXOe
n3dJ0yiQmkECwUMBrdhz2W7kpu8ENPg4fqTECr8KhpFCzjGgRLU1gaYISMNSeZdbrdcIM+n1P6/N
RZhqOrDxC50zTxIz+zMgq/15a6XETW7ZabeeoGMOFORofhnipYc9wFru/2jh9S/yKiRVoK28EUIy
VLfzzowg47AxGxVMCYqHGQGsOiAAdkgLHG5FwfvkvB2tH+UMAwZRnwHc1Lqem1G8Un4IgFT85g3P
jVwqeI27DmeOWxq9mrM4SLDyWjFFu8V9xNyII8jANrpLF5bME61X1mPmXJdmjdCcS2uZevCXGDTG
loWxjMEW7Twq3k5JrS7EzWbgwFSYTvNZgU98MIp2bjwYSet3HYN9sw827Fz/GAtvPeJJOMKvvvN8
39Qp/EOnuQThMAjjp3LZtPjsICuOg4Z8A/EY2a7lSK+xsAxK5L4hWW2K0dmFZ7PVBQEukYqOfhr7
d92yfleAw+KG87GhrIngVPGDaN/Amah2l32EayE6wYOLMOTc+DChFF9NILwv5IqfvGIh4IabErGl
90sbEe5hRNTNFIUbGqgxaCymoDZ/NjbLzTK+9uK2puIxyQWmsNfrf8t+ECODJ6r1BJBqDPL5R0eJ
p1k2x5p/TxE9le/H7mj0s23pQxzcwYzfTdD0iDimpE69hvXbEQzGmMT7ILbvQp6sUV4JyFdDdobd
Ulx9Z+C8g4E4G0ltY0PJv2w/lQqwIiY1rE5W46Awdw84FjKXd4QcBu9x5xJ6+/Sw0SSQ0RxeuLcq
sxfyeUI3Kzm2oHCZLfHpCFZ4lvbdSiBP7h1qsyC9S9w6908bwc/q7CLpqOyRC3W9uEAjMuA6ssVk
CqkYJsY0zhf+4/HXpgiOGKPFpkwYuPLzp/gzG1xyRJ7AINHWATwmsnbf9JKs5HN+ErBsqhqV8dZs
v3tkhzfW7xRZuYTFGba4T3WfP5hwwTIUg7/vGoWG+o5D/sJ+4TMWS0HyvhNFAMpMX2qUKqKzdccH
Zq8+Fd2Z8bGsAcSDT3en0ZZu+6In3/A85r7K33kilxoY9JzcQ6KE9vyuHwWS7I/3k9vys5GKegoT
YLJbh0PW9nWEIWTFGR45T4kpZseI9/9B1ginGMaol3/km1jZ/OBT20+hBh5VeJTcDVAvnSvQniOI
NScOuHbCCieuE/nKyX0XwXoyvy/bnY/Cgd5wtgMe2T9lhVwIBwG8QO91mYa/EnPKuLsu1dJozoLi
rAh8buqW5lFm/D6v6LOgSj4FXkZnH0jSe62eztdncI2LI5T+3rou0lfuEwtw2N/dB+N1SuJqrCVF
KGTqQmhJeha4CEuFJKUVCYZxiHHpFKGaHUrLtdgYyDSOAr/ASLOg1njg+YRizDapPXV+V5C3YFlz
wExSXxMpsOC52YzWy60JNLSYWFKS9w8uULG2kH/22ssrqa9xTBw7u27OudftSJoBFQHIaowpKvG3
yBU8h/Ltl0daryOKgKARgqmQVA8kRoVqJNm+CrVXCqybBGUfAe7WbjoZzHaXm0CMLlpp+ZMAbLB4
MWYrVuuG+35Jli/uwC0DWqPpMGxJ9xYB7Z/p3Sgp6lah2exAHYEZq2uZMiPJvx4lfV6TTzeqN81J
0V99kobB3XpsLMXslI4U0QXA1O7i1q92W8BU3QLmTk7SYH84qF+ckEVjcetdJpgXteslt8b0s4BI
HtMP8kNbvDCBXzNHeCG5A5QN68w6/iVlK/w2g/jY6LQH2Lg7db0VSgo2Nmkczaquqjk4vQK/e94O
Wv8pfssdIWYXti48HEuw55Tv9ozzKk6CJmyPeL+P3iEPsVzxmYJJE/5VYXylhcVOVv9WDlqLOoiM
J4Ssl0Z2LX3OlUvFJcr6yCqZSfxx+JzPrWweDocSMi2gdahOSFALpUzpxkh9lfjnpo4aj3itxNuE
u0ERKGaA+t0IowdLpdqstEp7+kHXpLMNdZBrK+DawGIHSMJUNwnAuB11HiLz/ukx6W+o8hX6yMsP
+h+a8K2u2uLK0LipWmZkdvPJjRqAkWsoYfBK01Vh4470GRqImTd1luMLmSXLxdaQqqMaQ79hXR28
aBIBd1i9Pn3qEVS6kUW8CjZGJYvbMezqq7tRZLOzkcajkJF0OG3Gx8siaXxw8vR20UIdzTl15hCO
GymMpiMFAhWkGTYa7vZ5TjtHZWPvEI2yeeXxv3Blf1+xpNyX+ZVtVnJ6LAJ6wVyRt3w/CRQ2yAbt
sO9ox42QLTQhAHUJMMm5ussiklAD6cAKK4LI4laSQmXLjKzWNeNMyUpkx+U3Eh677APATP0HGxGS
+bzKRUQftI4mn4TEbiVfdXJ4szvcB4rWpZZ4sijrqszebs/PnUlC5Igqbn2frDgezQ9UBG8LtNDV
X4y0z+/kopR+0ThVBLVaEi+J1ClK9jUkTcajTBD5u9XUvq/U6PbS21b9LkRfH6ntBhhmZAagyl57
J/ojrXHUHSiQPvfk+m8kNUaiTHjWbQWLtoAJAW63RwvnnIO3Gr1horJrrk0+dcwCQtvhAPonZuhC
gTaqc22Opk1uAGw/SiBsZ4RcsPKqevn0ATwpsUj2ZS8VduLClxeQDwL+iO6dD1lunh7ha3JiIBz/
XnALWQAwcdHuBf+n7tbqmA9zbZy3tlNT0h1fcRnXdeu6G94LAHY1wEpH+vuheUmd3zaf3A+lhToF
ZOSVk3N7niMvYQn2xYPWiM3T3RprWdu9xRwNs6JIPw3PDFdCI7TJFXE87NcYapFeau/PjCtLQTA7
5IlvcKe8ScT5qojzEXeZqL4oXbEQy4M+0oIj31iqBm4wFIk+be8PBmy8CqEmB4L834GPnT53bIZt
Kxh1Jb6hupXVpiWJZiZUAYVUrUe5Ct8yP4VifSimwXBs9DgyNoDVI5mICrpf/Dtsdj16HRypLfME
i0Nqt2uNNIQI5YyRwSLSCPSj5777mGMmbEdegNjMX+empSR7ZXfq/k7vstYACG76YVltW0RqhzJt
EAQb//bXcvz2Lqz8AxZVgzAxt6W2rYaz0s12144ui7Mp8lkjrPrXR5v3FT2qP/SV86J34pN0zBYD
uRGhGxwayqdGIdyyRgWDQULumb53CJowGCEQ3Re9L/WifMn/Zr3U+A7u10rq/95zD//ah5x8toEw
QcCBQZxpG/DHZ23+lBnJHKFxbQ0mX0RES4u0iaHpfc0cbjDRIrRYlKdqwjq+muf4qnvJjYWgw6bC
V06usEks52nKQdsU2rKNukzjxU++o2HBnV+K8ZJso0suOF8a+QHDCcnxJU4RgGpnyn8q2fxETV8L
LyPC0fJTkYJMvqoDRJ+TR5vqMPCtPs7TN/mJccrD3WA5k8PnY7yFn5in8qP5XXUa0YfADWPMEEMf
Xv2A3u4Cqb48H0ZfY2433R7xiT2Wnh+RrngnlJH6cjVDAhN3hNpZccbSbAhZdBq2JxB5V3CQi7Uk
s37KeTX9hVU2LtSJ55LZHcNDfSEuOKj8yI7TpYjzZjK08AaAKApUEGS7mYVi0O9n7sFu1ZlvX7+A
yF+i61wk4bX9PPG0Qrzwc/S/wlC0MncfBmyAaqlR2VSogiPVcCCEzbjr030HiXVF4b1xQ9kjumV7
K04+FzAqwVRc3naP+QqJPML6cbxlvcMcV+HXx/3my6YnQcf6rXXcCidxN+UYJdhBLX8K6QdRjCuz
gNY3VFQrDItlpWg2nsQ/zxg+S8c9g6uJOUJFdnydOiDL8CG4U2kjUrKGpwu2i9PDh+tw0SEU5/9E
+zB8rRKtHYTfpgTLIro9Zbh3Bfn8PSj0w32KvAlnUxf1h14WkSlNl/a61jmAAd+jVfm9It7x+UUZ
1OjCg3fNurQ9rm3HaD04nMdj8dfcoJEJFASBkPz6pmDurTiCFhdhSsuESwo/DQVRg9rpcwnftnKQ
rpTQKU582DYtQr0SKCngjNyei8EV8z4lNQgGd9feDS1Vic+6hZv/OwDnOWn/Wd/dyLGhTWIkqLcE
MpoR82RWqViq1g4Fr5qZFUliDjiSZDokzGGGG5auLuFkiM6tMHFrIhxwngWp1EhXVHOogrloiUhV
Lik4QsUmi67/nQJEo6ds/ZraMti8lt/mcHPF3m9fYzNzV80bbv9gNkSUz5rypALOfd3xsGGJVS0R
7bpANdi3Bc9ut/iX/Q9EZiBHuxktrpSgZc+qfen3Z0npKEQ+WLqmlpCkZvjAa+euiNlWvzJEcIkL
HX2bs6fQDcODkIDSxpIDuamyC71/VN8+0PmEg7Z5y01yEsnKWfssQpxkZmaglAGr2IVgVZHp1Q8h
fEubVmpzkJwwhNz0xhYqoY6sz3vvCjsaBQIKwobAIyE+JWurWfXABFJeAm/A0N8DOpGNrSOq7yEz
UX/XMVMS3YS1qiXTw/9CKtd9JMq7DruE/ze795VVj4DKJSt2sxFArw/DyHApzbCM1jK10/BmwhVY
izUb/sKgKrOJtqXfPYJJ0LyBC8aBEm8lQlY8AG09AJlTV0bjMwBWdGgdCwTbThDXZ1bjJ9flUxtv
9arOytLrrJeebKrPnJ+gHyFq6MeqsRGZ0uxXcxeKP+9tM0YPEQemOf85p6DMmA3FVBYkt8I6Pgdp
WTrbLcsHMGzClhZvU+BsAYeSD7xxh5D8R0pa97eKANAOawqpwWh7A/jSwUGZwT8wgebRTsWQdsq7
2fUFevzdJr+9oIUomzDiv8KnHCKc4wBrtbltQxd0B9lqz0xahqJ7ItedG9I3WosUlzh69hPXnac9
BHWOvggQBV4Q8h5ohsTf0pYDml08hM2Au7N5MYOfNEXzG4s0cd34ZDaLk2jvsX5Vcek0eAGfVdLR
qHolOY/5xpKDPwScAwh79MXV43i6pntGoN+GYh4jFrPkLkvB9NkHXvc5sMzkh4psf4tkC3aqZnWK
6tK7HTc7M2RZjEo0Fbplx/8iyXY59lC8IwG/HR7Q1zJPpJOkWr/7lGx9cpSpKMOSwqfGbWGi8EiN
hKF6485/AeipXL0wYnvt3JofG28zwvLXaRnkUBWSiPR4c3WvWbVvZMlp6Nv+EQteRrUJi4EVru59
p6JGgki9W32K5M4RfuUTHoq9mw54cQCdowbF/SBIH33AcBODxRjgKyl6xgXjSgx4p/+FqyiGTaCg
Krdhx9ekmqDlYCRqs9CrOjidkKJDaPDLx0mVuXyk9O7BaKzZ0qfvb/ZHvQhraIE/m+Ik9Zsomky3
vmneml9noYqPntwI81r3KeYNrSMlHeNC12zk6SnTypU2lpjBZoV5XnPbdbjj95Joql1xDo1e+LOF
h5/C5aPp+00qR72bQ+49xhSS+tsHS3J2BWQjja4dmraKl7Ih3EJv8lVSQmSiXqu+D7aiM5rkiHvb
iVCUDHxIdHoAbemycc1EIioiQu9L1jCbvj5rawcNPDUG3Lw9K4hEQMr7snMeqTHtmuOcFUM+dLfh
GyZVOJML/Y+fZqSjWKpLcPlrnceIRjG1KyCC117b+rmT0teYNP9JPvPMmKtZ+ammeMD8BJNPadSa
vH6RLk4xW43Eoq/Ru7v42WXLeWskN9PLo5saQBY9+Q72ewxVqPYQrmtAWwlihuJYWwTAzduizBit
CJO6MVMVIKOCpw501uClSZUGmIUt0neId+MOFYB3Mypy5D0WmpXszpFlEeyyNSBKlv21lXObEEDD
ihAyNi3IrLezLxmlEoCES8XLUc7Tgy6DMLOPus37zYAPk24X8QTW5qsfzIpWbQQpWdhlwMwwamdC
S7oqhK3VXMo7pOLi7hzC91qp/+x0ObbV37r9eF4VWyFAT66MqW2VAHmqISvuUZDb7pkoGq7A4OHs
v0F/viBghMJGHPWmq4k/j3Woq3rYo+Nqip1IWFO21+eE9BOe3s9yoVBbtEFpRJbxNztyrcy78jwR
qBFILEWuMzt/VRL4sTFDBnAKjyalROI9sRBjatKH+mgliDdWOksmfPpzLIYKF9V1ekreePg8IJJ9
Umr5NUkZSF7m4i2crlRsKEHejgk87090fq/GyXn72wI/wFYQZG0ok6/w2ITKGxtpFHMlNYWyzpQL
Ls5l1BDwYzuseXejPtvSaXGUmfp154PC9M+79iQiMhYS1zTHlcHeIIRDOtxjJzG8EA9CJA+EO5zD
LLAV80E2oI6qVv3LZKCIv/USLDOTtHRaG/3bSy7Za7IDQLA2Qqm6GfkoG1IFL0999oRsBe0j1DdC
6zS/0CmEgGbTOlw+c36004Z1eDvZTrepPFCi9jRBl7FJkYWlx/Ajota+0LM/WJfCeLjQUaYG1hK9
34UpNi0siqTEFOxnyASa229IBRNgELkKqeOohtkAFU0YLxc0cQfDcaLnqnqjSEesOFWhP2RPW1NJ
WsRAyswz4xdQimEvLZK0gtsgIAzpqnJ/ZG49MRXwgtvlhFkUW6NPa+2w9bg1O1tjg0SlgzhAjgTV
artu04itqmAVO22JbDNINjY246IUYir6DGhw4KDX8Z0s+8DIcQyznXuXg2/hRLdWl+c63y50SPKx
hMiT2897lJOoD5gsJQel4XexH8GkgVPXj20CDhRnlQxvCYOXxRULDDgFeZVdhnJsONX2vTdu0jVl
jrl/Zkh/MBGyP4QWvxY0s0nsUcFtcGAm+wnBPkjcNQvdaoiZJH9zHn2YbndzHlyQUSWIFPVoENr/
6A51Mn1C2XsOJGgVyMovzraMeW32ehYom1VG3xGoSsZllrJd4UUc1nKTBOgrHDiKML256YTSLwgw
84Utuk0QuMZVQ1bfWwO55/y7Dip4b7M+f/QsNBGTV2q8AfvYcnlhrj1/zZ3ZuEhUW2yuu33F2Utl
QZqOS5+Nx26gcO4HlCn5zWlH1CajCfCk1FnsEFNDxxBymGGSOFnB3ZXwRjIFS+8pkFRvbTLbo8gz
BQjVCl0hIbZsYhZp9edLTvaycPyzxMDJKFqAHMNLpEUmFAz+hyZUMw+Ib1r1H5J6jogRr8Z0lDzk
vJlVSK5Jn+fGRQaEPMWt3twbOaRdJ8Biue2XYGPwAojWBgY2iGFZaGwP14gR0FhoPXkKUU6J4Qxk
MFVyK0Ik4P1NHO3OU5UOL/HX5sHK5bgv3tTQk9lnZvHAzXBmBPkr/H2g3VB651cLzHIM4ZwCtXKc
qYUrR1qtQbzsOS46/B5sFNL0WTprvuEMYB4B0AkK4tFmoL81Fg4/F7pgeIvJbLbW7DnVWn0/4VBT
SU+MouPzPQPjlHMq4asFvN87lHgDtjAdYt1Qc+j+nDvGqgPqxmNMRMN6XSAWMmFfP720DmMTVWMb
I+SJqckILzKR6G/CQfa85aIgBCZxZV1YxF0HuVfSl7Ya3dMPs2qfqKXmauOORVcariqTWWMKKE4w
ITnkRIbIRWN62Wr0ThWc+VYYUlSuz19izDL4JygDTlCxmCtjvkpZVvndfW8jU+0rPbE5Lmu/5rUX
YOaTWLM5pihDOvKp8WkpImOlF/eSBIAI2ujXldSz+EpCUrADtULf0vOmWdp+RoLujSrp+5JZNe6h
IumOW4Z9xe/+OQpIgBdn7w3zaX/a6BnNOXiDioMDakUMq9L9XHXl1led8alrCIoI9Ga2VgkMIGxx
T72lfcddawDXl33mq3LQ0gtToErUCpntyC/ZyD1EwUs55sImGTOgunnlwKdN3msRYn5uG7zlewHy
E7Qouwn/OFjce56w9UXqag5UcPh5eDc/CZV4WGmQ+gVuaWTa+a64vvIQW7aGRgng9HpaQoyHhwg1
BoAKWDe3VXX8ZSKV2PfRmL4iTzK2fuvZ2r6RONi27W2GF53v3iKJlgitnlAUk8V18nVs9nDfRG9J
yA+S4NSEYpEdQmoPRNhj2lEkaREnfnJ0jyCvi53ZRFosoKKkXp77C2xoCOosEbm0PopXbA1y7bJD
R2oOcSb7DuSF+EJO2Dd0m9nR/h/MkoIokg9Uh3qcusOdtZlz3rzXQg89vKacbCBBw0EWwh3/43Qi
UwfRJHTVT+ZVwWPVd0+VTpBl43cQXNJffi0exLsFz1Zl2QlUGA64a4sPRWYMGe9VVPrnr3/AMQqS
ccD+BQ+WuEJwSxpSTrO1dBDuSKwVbBERJrfAUn76moGo/PDaDBzYU74AtnYZgzSSELAFwkf+Uki9
OUy+7hsl+j+apZ42wF/JlgPPet1uKhxzXHXpKRzIDng6FSCSTtDiufbmGy+ze6Ro20xl4prLtEkS
1HTwXWbOpi21Q9C/K/hX7LKOTs/T0chTeJo90A1VG+5B0SM/NOE716gUmFuX7o6wZOPqq1/nEyHn
Zfz8z8pO8UBy0HCMrVXJZS4RK/MerxWuvDcR7Xfu2RYfu6RRu5i+QzlgMiMwckYdc+/PeXqMdnkG
agLMVQUioumq2kBxdYlFQsgzoDAuqZgdtHXzlL6B8MoRfA7Ec9AJRlaa5SDAM5HBS4lTTD833zfx
nZlZ7KQu/k4RneuTZ9Q93kCkS7C/xwySrSjn9tvYD/H/DVTvWwXm3pwIGU+DwyOl+R7K8NYBbGij
DzpzEIXgrs55Vnuecaz5spsqr1AeapdRETK7c3EzJRRLFiLKoFvb6pIGEdlqU17Ec8eA9OPh1/TH
JzJah79bu/8GRWdTob94XDN1edHXqCuFe3RJbiopmjif9Oc6Yox71/cyG8ySG2expnsKKHlFuUC5
JrrZPBpYglQXE/kczjXZ3xCpAE5z160EbdFEkIv1Rnze1RSBfcx4k3gEggVgglGnyigIBMja+FXR
BOe5btUsh1m4+a3K6esLEU5JkGjiBVW/zRu0ckbJhRmOi55UI7to+xZzwFv960HsoFOC20DEVdif
/VUuOt3qAE56R+4XqJ0cbX1VM1IxOU6vncjT3ydVlcx2GZvooTB46167BfAytap194ZrgucX5C/4
KovxcnOvXesv+YGn97XMBrZ9Wgs9xrIrOEo09+7EJEuSuLRuBBViHgUuJkzw4epN4DAqXeUxf8ZF
RVHaOqDZRaMb77NHyNO3uCOICtHAcP3BB1yxm3mU89zxjM/lfs3uWvuyXo5haL3FyzmvJcTGpW4D
nzGUkb7c02coBOMnJM2c55V+yzGiTGdbsy+tBynazL1cT3gVoKPsOMe7dx4EQi6pFbOWRgDO7a1K
1JEz9AG5oPIsV0gl+DxN8IYfPTIWqCtaeq9q9wVj/SIO78CX9AKJnSyfkZzpr0OMPGdppQMBb2Jy
1uVmGIKBmM+yEQVU+1zI+UZnJO+SzBlJ5hRC2NPUbfVw8IBcgs5oxqoS7N94SrOYLxc92YPVi4jf
6G7F4+uti3oCL9mml2gh2pBemVow9gMATCmAoiyhEq0Qqsb16ShaohSriXbq8Bb3VRSorOkzYirx
NflTp5fblN5jRgCkJwSF8JvuWKQYNCwZ5wxpnaWJl/AXVy/RZvjpnigKwDwWLOauq89QUAOuafku
ICN7cbQbVSIC8k572j50clB+SIXeWak/Fd0Z7KpaXMlzqIRN8JDaGrjAdvEMQljOrUHUOQTZ23xL
l2GQqmqEQ9uSLYvU3vt2OlvzpV8mGz6ygTneWQ5PyRkc2LzQesBfHaEBfyJksxVkygoM7t2uf8d/
HWMZs3YXO8o9lZnLRTtvGXyeaSsA8NFIAb738VC7Gs+JJjTogcDJZ9eeH9Eslt3ARhyKbDCPfKqJ
AgQXIbpO9iVtiDB4CG08Gjd0dSit7gqnN9btcxoTB4NI6IXQheLslFV+Sbo/59p5y5DiKR+6Voil
9n1+LHJLik7HJt9aPutk1W9YN9xn3RnQmA0e7xh/PL6gfwQ3+cbp+6R2lY9DTloBnbgBGkSmn2/r
mRum+hg4ZUnEHF5OaSPB+4U5QF13fO08voPS3KuhX81mMA2DyZJSWn+A7tCKjB6Sg//IzNbAJyTR
Dl21ilCSSX5vncKtbqbkLYOzCTke+EJgiO3aSQuRG6+95gkA0J2S4IPul0iau7CsYdIuS/dLVidb
rzV7PKb+l0LRpFhjmRKBA6hIAIGyYrNbizxenkV8WnGAGnD0h7fISaTsux8pUpMvqsQtzUM6h4b3
mTq+yveKOkNNjs3GDdIjkUG1AnlfLiteO4RqYts0PNIvAuyXsQdsvEwi69fgU+o1BRll0ruX73UR
BlDVUE2UvwrQPW4rQe11O4mlTVrWBMMIP+ot36Vw+y31APhUe6z4FX+6hLFnfrPkj9XyumnURz12
z13wcv6geHvIXBcbvA1p5tyO4p96eWn4WjojyO5QuvCUsNaWHsB3X5YlaB0+zoGs4nyqCLqFcpOQ
RDKQttzcg/D56xFuAQ28xu7sKSf/RMRj3VYQC1frYoua9b0O1aBAk8wXKm4SjC3Te3uYh1iDsocK
IfLRRQYJDpId3I2a/8jO7xu+UWbrbOs9imMrvmIq+GYWM95jrBMTfIrb2o+5FZ1pF1JTYof0ngnO
yGAeYSCMGeCvwvNAQT7ORipetK+7tSIjIqJOM/pmPb6/oMnt7pihs7JWInMXp3yhXDy3lcODu6TN
GJcPauC9jTbNH21OY2vISmAtvRFi4Lsi3fo44A5CO8C1DkWgwEsQ9O/cuyy9ubsznairkJhL5XUt
w5s0Bb2RownFmwWWdus8Pie4kVqU3LWLfexql2g2MAiMgW9upB1bu2GM3WCuWkKg1IDcCPH3+Itx
b8mUV6AOSAY0IAiqbz/6+YSLW14lAS4lTFhbRGwpOm1tdDbaur3/z4r0BGBTbWj332HHAQzaM8j3
Gh2e9zKTkU00v+AvTjtTLlsptoBkZnTavr8dKRmj/MlmJuez/x8qM/cRG7c9ZrsJbf02NpM57bE1
XsD2C7nkv0e1xaeUkfYVfcfxINc0Vnj+Q3iHZi7ndoQQ6lP9PapViUEI1F9Pfx0CNjgbsXZO94oD
pI9V2FmKYJdK/otKhcjrLeudJWCBjzWkMiMJnQARxUcH7jKBIvKmgaLRkHTiEo279l2u8QDjgi+y
DoOcHnqxEkHjbPnAcKDWzktDrnM3lOrRdwudHf4sTyXR+tx6U7Z9xlYNkPS0bYSDAl4wWdqirsCI
d21AyZntvLGTkNHGMb2pe3T6pkZz9JEKLEt1ualRnVxQQxYR/kAwcYEMuM/risH5H4GEJaloKmGU
3RouRRlvni77GVAzUvyw4DS9Xq8gQQlqOZQ3Nvluy3gmXn7K+PECf8MVVaYVGreq8fS7EtCPKNvM
6MrDmV7HkLdKblGqnQvw33QjZ09H3Y2UnqbeF9VXzhKIUp27m7cNHfvIfgH3qkKvYo3SIiN1OrZG
eeVyOrl/xZre9HRxz68mAnZjm+PzxewzpplK8fWuV4GU5MB3n0QZrLYgiNDdxEtvVim0DTOovhqX
sYSzHRatw0ncmmZXtcC3c+0nrOgbenUCme6qNsTaP74a/ZgnNn7XSpg3WWNsbxjcOCV49CXFy2Lw
ZYC32xFxjmjzhLVdJIWd1Nu8ClcJlQwHqx2vbBWPKDQikfzzPaJ0YQGE7q8uvCBnSv3ymt9pccUL
dIurU3IEt1gpekzNcW0NOLbJ8fOYsx1RbyKp+CyJDmg6nLc1Yuwq83eFt7Ln6L70Gkim/zJwO8GK
1286vS+xuzv7zbaZcFNvfRH4AJC7cks4zKNn6SKRMsXr3nV6laFSZ8Xg8yPwImJ9y4ofDyjyJfOM
nY2kajhzIhPsZJaSsqemrMnVQ82tIUbCv8XfmhhiMqWj2Jpl4OgFoG7TU1+6B+NZAA74XAFMxXzE
CGZ2Y4oNO4eUu6bnCMcH43T4neDh5h+7oa7SYEw9/Lmc75Txy2pYaxeToSxwjatRbWYXcC7Aq6C7
Xg5KXm8HZDhNmydRIF2F1YvwW+dWNYBmZeO8gFB6D26AMNCQBdNLqLCHVeikKZb6AYlRTcsl8H2y
+fCu7Wd6c1A906VoljQHKEPSaJ0nEx4BiXeFZ7MtWn5jP2gPwzP0SiFWqYvzjKrsimoynw87SS+m
RA9VX5LrOX1VrABRs8QJuG44pTGD/2BCPhkzXVYZlqN5zO9sDBdIwE0YEjNV9c5LdjdtSFKCts7Z
s4ZNec2Ld6kUDW9aV2/JeEG/TkfP4HfK26lwf9PyweJrl1/yvsXJvk+MJWYfiTLh/vGP27PBJEFB
olsc/dgYvxnwtEXSXS/qJ2EKzESROFTk71wx3gbw6o6ArKH4kFxxZJjHYlrS8ENiKxXA+movN1So
x9bzgHfS1qElTyvjPpC/MT2+7/w6G5I+dlvaqDLoPTvab4WJs+JLGFh2QcAJeLbCpqPynJQBv60I
hQybBS61j14AGVwO9JxWP1tKQBPBpOJXRpvlbw1AyOsoD5ZpMZt5yeDg8hlPOsmPJUQUrWY+U2pq
2BNuTk3573K14f1htVKsd0tBW1/wS+WiQRYjzlfCrPQapsg8K7uQZnhE7UxQNnX+eVmriA3D+E9g
kVpO5M7qqluC2Nk0Sre9MwVQM9+HVd+7JsSDyGq8eC4qesoilcxmrQuwWrGlkZvyss3EC+qsXOoK
7f2k57giuF50vLbOV9jsxOHVXc3vgKYRL6k4dM6fN0DLTAVKDFxsnHF2ZCDrk53dJgjZfDv1Sufr
aBb48nl3K3TOecyf+s18inR7DzDDyxymX00T0YbfVZoJJJZLO9AF/HplN52zt9S466L2YPouj8aF
WvF4nqTRsaAOEKuQ27idZwy+5WDacaVHHt60HVtGq9f8H8xEK8CxoyIic0f2cE2iiG+bqY9KCdLb
Mhs6X988OIYZe4UmKmnInDL1u71EGv9gWU9pafckUpDae9vee6r2dUg6VEhIKVtl7hcm/zqqrmqn
PkKFYMVFSinhCUIIUw4GaljSMU1F4R2QwNZTWTxtxPgc5w2Cx9KxglwbhWE28Cyhw7QCwl6boUM5
2kQuP/43Ht4Kd+tINVhbd7jqYnYhgGdso8q33qdEPSvrUm0Pwj+gU9/zL/WwbbNBieVa7n/z8i2R
ZR6QSFFX/ey81Kls/ggD+c7lzuo8y+SEnUN58SmBO5Q3+VUMu9o+m9KJ1C7vA9mQl54GExV2kwNb
ni/+ptyqAudnbTRmXRXgrBtcWbF8uP/6z9McJW7FuPRft/2tbCNpTQ35m2w6rmSErHswuUb75ttz
qxgCzL2xUJUfugiY9aCoYEd3eQR0tdlohD2OE8SmQcxUShUpZFusLw0aS3oUBLCN71wlzvV5UO52
Mp2iSEKfk1u/8DY5+RPWJUfuP8LMAnevvntRNUbIFhRD70qWZmm+YhguPILjM1WVm3bj8NfRNCTm
S7XOPfDkMZYthlC+bJ3jEdPPnOh3tzpGqw7Wu2wJh1GjDwpY4Z0UEIO16ODe0D5Z1XAXIr4xizng
l5u5DkEXqyN5Q0tElbnibR/7SY3SqoV+mNOfN27mjoLNeFVwEi3dBvOmM4UWS4/T1sDlHpiNkCB3
18vhzfWXhzOullq33UzQJo+6K1qhWnEO1UbpMaUw8s06d3Oc6mRAGqjDgLlH23/+AwomBSZ/llme
MHN6IB+H1EtAt/tQUIFlBn/QA964tqXdr0zXxHCjdTqtQZht7op/RMd5jQts0gT1OWClVeL1Oax7
z8UYgYxeOzsyp6RcWlk2rrtAMdNYmtYn2m2JmfhrlADQ8v62Uk2r8UcuFIQ6LDP+1b7UAWgmOtmR
1G5lWxxOuBezErxrcP5MzwFkckNfaMnxAh2IGwyXcWBhBXWsUVm6Gi/3gOP350ERTxG8TyyZlCaC
FRL/ZNLmpkb4bhhNVCI6zguNaueN2QoglHhqP3AabqOw9HmVIsjlp+y5ECmFtREB0GrQDMwabtHg
PnJULDaFg84ZFzbpenbTi86lAnEUPV9h71ruKlyga0lzu9PRJZp+TFqcUPbJHHQUsWymVfjo0EvN
ZM5qxZhQZbuPLgPejKfqatU1oqCLZn29MP7+LP5R2jwVIm76A6UgV19iupsMCazW9m0mbPXhoAas
kj5J57Y7x2k2UwV1etV8ZcHnrXMErUJSGzlImvi8/ug8zNkwSKCL83X5uo791Dlreg18sgGnC0ig
samnGCZgIP1AHqrhEUH7MRnIrHKb24OJaSO6lGygenVFalc2EGTg0/o//EQsvpy3TBC2MUy4DbuS
iHs2SUWa+U6Mjf8pxQCap+5phzSF9TsVS/+UvY/cP/ZNOgccogvBTRk1XnMf0IGntdAbPwEED0CI
wuaTbT2Pc5tmdMkeBaHFKi1SAxoFENyZT4wMnBcdiI1VwctXiRBfW20MRE/qgVLY/HFTV1c7QdpM
goaYJxq0aMWLiPWpzzEh3J3NbN+k3A860usEDxVCyNgY4q7PHqT8KovwaAq+JO5EK5T4jEuZK8MS
+EpKv1a3ib/i5tQCGN5yQmLx3r+6+Bq71C/YplIxZwj5avzHbqCpYoXouT0QfGNuk4k8S7WLiYgv
Of+Q48nlz7QjCotVeEPGdFsg9HOaBZB0vHtqnDA8D0JDXDm+hkclHqlihTwFJB6pP7kx9Mf/aDf1
/fKrz5kvHGBSjqkQ6k0Pf9uFQHA0mtZh6tSUmZhJC+PlNxbKIwRbNErXpmM459OwuWLaTniUWStt
2FTLwsfKa8HGcNUWSI+T7AYymBu/xwcrN3aVDz0F5RpOZMIGSRMtszFvsoGfooVzcia/0aT4Dkb0
mtCuEkctMlU4RmUm461mqJCcfGkzbXMLv8qoj+8mpk36b5syWTej7za22I6fkpdKSbszOzGD5hGr
8bBtq4l4sMbfLL8JQUkeybdopeCJqC3u00wmKPWKk4/N1Vey7wYbw7AGF5PlOMkNYVxvbc6tNKS2
/+FiPvXemViyBf1dpEVqlJian2iVEwJqL0eoVfU5fsDeg1gtttCa2TSQ+L53qYukRhoVTTnmgkGb
d2W3rOYwxzcffgoPEWNGodaQ0LjcMYiVsvKpDmlettjuZJT+Nfr+Xg787KHTdVHxZHiYeesNZu0M
RgFWrtAr4wZwy6Tp7DXkUU7UVtZzkB+soDtBbxA9Fg9/b1bO4Mr15w3dMgoOB8WOLrjWFQJssHx3
AvgjjuDUx339KFI2Q3ChwGhmv2S84FknVglp3bi345heTrmAyVLStvzsUttgWb5jkN0zRlkiwSVH
omX49OT2xk74HHCi9I8faaK97FXN7fq/X7aNqN7SkGf5zQ9WJhN0vS5zyzhuWxc37A/3WemIW7dX
BQEMFR4DsOlTKQPjphExlBJhSAgmGo0D6vb7RPLJfgYWl18JVKvXisd2cxQErmLi5HKpsn4dTw45
j6SNKXshgRP0fOAUMADqnE59moBtMQhPWDSNqjwESi0AIKUbXS9XIzpYyWJsvIsxCYWW4OeuGPjr
/I2WAgi5Dt/xwlmblz1jOIKDD2iUl8haRDyiseQBHMqSD0d5DYdiLQEz7wN4HO2yDVGi41UgR4M0
2ex4QA+6fNkuIjvDgutMKnkjhu0oLyhtSebGX/7vHBrbaPhMI4T6w4we7oM0EIJGss6JLbrrndRN
+zYTltc/54Apo38+hkPK9J8akShR4zzAuwVXfY6JfxcO4lR5rO+vacqXmgWB8VHHURj4IkMJgyow
B3h6xneOtLo9RQ8bNewYlChXPv2KjAXpSjrQ5oarz0l6K1UQ5wcLRrwy8uIUx2hIIPVPLlC6N1d+
Q0l2z/bfUfWXWv0Rci8NVVYIR6LFSFab86wwXeLUVsrWnjyPJ1txng3wzt2RtYGrQlFjdMqW9eTg
pluRnP0A9jk0JFZrSLhIbi7LsbmeDcMViND2xeN5mCttQyrtowha1q+iZ/FeBFEcwQtx4Pqe8GNn
rc+Ej/VdKh7Um6T895Skhmr5+rCGjD9NC2G3H7WIDX6u2F5DN7ksltieUSZioXFjDQxzSwsNi8TB
UkuXpTJ4xiQGkWOjM+fHzY4JYImmBQZuOPn0lkxJrlSd9k11r5JYwrAcIOAaiukECCEJhQh+0UHK
wa4T9tBpjpCXWa4ztDIuezneQCLJEAzM32uHvfteDXG5EiIOzV8GcVJGcO3y47oZXlGmNgR3uqGB
4SxxTlbao+EV+moqNKARdiovp4Z3RpSBV2EmCrSs47T7vSutF2vqZN9A/fuv1YThoBChAzZH1PCq
bTMUTjCRubpJO+lPcWKDv3/oyQuLOnjijdV7P3lsPOrvQmccjuijxv9DGIRlUYJTD0Jwk6/XgSze
3wU89NDZj5cMw+P1cROr46BRuJ1lJyQd8mCzAW7yMGOU56Xd4vnglSwb/tz6u/OYcZnQDQsT949O
2ymHLsoNU81AGC/1fx+gEAPWCfWmxR9jEipWy0qZF4+I2wZsfVLmTMqYTPJ0gvzT005QLxomwHrY
Y8eOwZnHGB6dDQmCbscMEEUTieh1K8BH/OI9K8rUoVsMATgz3XazwhZ82LM4fSqjCJ5FwMk6AEtg
b8C4SLZZiJB9/WGv8uPvjaJqJw/mS7c2eglQ3788hAlBLPz8Iu3JZsAs7cLpzj2SwrLOMKM6e0FW
3zfCAv4mOAZsOuz2XjhIOhT0nvlk2zisVaENjHibhBkTTO08aGaWmPlWRjpTwpRhJdwYgbd2qefv
mLh4s0Mp6Xv46Ej+nq/Zw2cCxC+tNM6+HCsM6cL4+MewslVYctBnj5W7LGtGKp+o5TUiRAeixx0i
YL7NR2NwRm3VRxCaEXg77G55ys2yYBSIs7kDFjwkfvFRWJ+c79vQnplXyoMhf1n5aEZNF5YhRJ/W
3FnhvF9PSHpVY/z14Bkf5tQn1R7+j0KdQHtV9XwUypBmH7cH4hZlFQJm/PrQOIEHmJuo0eFhuLqq
joIuFTqlbFvOk2omBhvt/bKGqJJqxyFbtkkGKAZZ2aYM92uh/OjcasX2fx0i6V4/C5GpCE75/+rt
EFnnSCZAl6ieIsEpZv8NZAySlN2bwiabjfQmniVkF7BfiEHj3YFgQQpJkRWQgXv+7WKVpKMz7Ffv
hNraSuSd/HnGqNdGb717FT2/V6cP8O7qmnfOmA+WXRHVCNfXg0708cNjo8K7/ukI2CXlZiN5SByq
pwIdEwvQxyrdfdDWe6S6yTf5jnaKobjkqF3bFvuhCibK8SK0N8CUjE4aIprFV+MdA+mRKXG3ezK/
Hnym3Jxj1p0WNafE8FvgLUb9ItiapL7iEZjTv8CTVshHDQMXX3CClptmAKu33F7uz8hhyt1NKWbG
xU+aDfkQyGcyMNCIj0LyDcw8J4SwT2zy1VF/oyJViRyeReHDF88/T3fHmWM9l2nIUPjpMYRIpWZA
RjarJ9jSXSCZtVZ4VYziMEVsVRF6eV1cs8Sfe/KpK1CfL7jMTp6rfkk5BMoU98RirZq94WCRd2qY
5J4JPQhtjBiAvQCguJpGPod3qfcqxsvdwfu940b56lT3xuZy8YiOi6ZGPvdBAcFBIOwIPbqDIeqX
rl+Ckx3gFXS6R1RULBksFiblAdU9z3LnkjDyKxdPO2WsKpsbc5zjifCMQB2KxqQy2db5vkrd9pwh
o4j76mHyDamcSMJ4DgylGjrR1l6D//g/hTiWRmnc7dJlDfM96fQrMAk096Y3rh5a2wxD70m3tDrz
HPNirkOYNePPEIFFBGmpuUnLcu6kl9EtF3URJ6MvKLAWX1ErFWsKuQXL8PfNIOco83wrSTmzm5Li
KhBM3HSzah/vOLzDqcFXzu3DuhM2p+GzA+A+KzDuLBhFPBJrT+Q+DEYNz/kF2TMPE0o/kX2rGdKU
4UISIZke7o385F7UyAremEy875X6PHZuHXvxfSgGrprnYN0yai8iBEZdvfKasL5eGqIv5Jymbn6u
A76B30rwWz2I90aEWEGi5wkha6wqWdIEAgU7y2FqmdrYvfD+CIZCZmeQUlU0R3IpgexxXzNDN13W
fio/y00NOCa6b0AXkzsr70sMqZv6x4pYWKBQrOGrMZpjRlzwN1L82RmsByqyaeiZqyiSmOX4rX0c
G3KHeSFxw2pHElMFGcgXQXHh72s/JtrmHbTwt6HA3choZDSRVUn6YEOAeet8/R+4TZQj6F4B++xN
Qv5BDRkVAwvIKZXTTiMPVO4dMFkfB1rhDv5PzgrXGPGxvwDsJofVsu3uE6jTsjQZ5iESvwvSq6OC
kcV21CVWm2UMbiTRpmWNkINwPZYQQAknVXsgZ2HsIOsVgRf2vtCnL9ccs6qLgiE3lTrEPP7TDDve
DhRQ2X0qLqS2rYkpuDig9ocZjPiCbrjtdmDOVdeRcaCTmHvrRdYGj4O2Axazn81b058oJLewFsCy
26REsu7rOi975ZQ7EF37xghBQUgD124T6/TIWY9W98XhTQr+0eQ/axQqddK7Hn8Cx9eb6Rfl6M0z
f6EcdZCKiU/yls5kiap+bLdl16fLBfxjWKBTCWmGNBIYhqjG3wSyJBJ2PEnOuMlPDhpY69ivbxIf
LNmMlFtWgAVJT5Z+dnzn2MbbBXWV3442eEWMFhwU39GbmhjLFxJPTWOh3yFk2OygWpzPjJXnzibl
8wXbZDYbOKdwUw8f0hUm3Qz1hCb7vpTorcjVhW7AUR0kimUEO0Jv2RuNQ+JoxeU96lbUXDWkoOnM
/VDJgtQFkKmyKf0cje+D9LSi1MNfFSWnLrpFeEgVUktkKh4nCHKEqFbgJUkJBQNOe1ui2VFCKVzN
dJFwhr7E65oLLVBajGEaxWYm5zNoYG850cPywRWpk9s698ZQ2CTEvoOc2AqlYQDs+VMJ2KZSYAry
m4vNAp3vDFA14s3n84+6v2jCaodEvKY2Z0YxmUsRG05agkTIRPB6ieH5/f6+7G/C5RzBARP0wFVj
ZfkPm4L9J72OMsqluS9M2KahwrugDXCGCJM5kUOxFRAvn8hbRRNy/roVdu+61TCHmUgsXIDBwewA
f6ERU5/RnG5m6LL6zeuotH+22XwyxTeZSVUdSMDY/HdYEYPB7Vz8ga4/1bj/9k9yyebZT3VXYG9a
cYaNhF4d0CpFFOE4yTN0qcdxqjd4hISVe7s972ofZMbrdIxhQF5Tv6Kc9nUtHPd9iDXW6HK1l9sD
VyFHh1FWKdYD+JmXjoQPWJH0e9PfCjN7ys3CJ0vnT9DuEYzCLEFUXVjGIK1l2/IAtYMRIwRKMzZb
R0Eb2vUQ0C0r2VERwbNzpDFYH9bX5Yia/M8jYVoxxRfkYuhk20tQefxguEbs5k6pfiGhQXap6dfQ
04Zi+S2M/p2OTD5r23dT8Z1HV6wbvoGV4524OsJqzGuLIpJvOwroANebDj+TAwLwE1xlzvLtcCVI
2qZzgpWQQ0l1bD0pnJgI9ftpRB4sqqA83aY9Td0EzFZqB/JX5+FztOzlLPXAG6Q0qkwn6Ke07qlW
rxzIFWHTUb07cVYUbzx9o41xKyoB87lnN2or+DGrg3wPi2DS7BGrFRp6hjNKqEMKSqcIuiUqm5EQ
C/rV0rz4NqQXFC+C5o+3Q8jObDqk5mcWYz4A3LQovtNFWIsuMskFuLqywbMREwz5Czo2XNnaDsKO
6VOxIdJQMUtULG9xDRwvwDnfxBfJ7zILQqRkryiz26E1aG5l82YQqKumMbOOXm2MWzr7aHmtw4Zo
H4q0aIAyVHsFM/otDyReq0O9A8pRCUYZLzy2ShOntKZeTctCOO3g0hR1rqIOksXApM1R2RJ/MJmf
2Rb3bR2sG6GuqUS87c/qyYkiWvrkmoODVVnhIHl6YzDmEwvOUfQdPtjSKJnhMUfFEUwDtfBQRWx4
AUCOFqWCjxBTryXyvZPyvBX8nH4z8LnblfMc5+EjH964dxRfwwuqeGsyAtKOeCHDBa9rn/3YKyH8
UXU6VnZrbej1f/xWjH8SYRS8+86tl6yh7od5G7FgiWPTHCvsIeiC14KYrOcT5dCQ9DBs4evZqq5R
4TBgNvMcS8SUYn1hjxrAHtK4Qga8wmfAo9oQd3ZRdDlrUa+u3UZowcMMB5jXsCVKw4Twpwhkg5XO
nAll7hh0uFcj7uElVOt02LW46G3V5RJdHWkKZSynlFXbABQ4QzQy/MZFrhj6iNiyCk0RpkpsEG6R
Rxxb2pKYqunmySwa+1Rbo8zPIOtCkcvYuGHHCJCfYZ4lExhvTKAs7x+lUvT69p1BXDWVdFDz2UNX
JJzWZey9qeDFI+zTFIqClsyd4LjEOOayCl08ADTOUBe3bj0bnhK/oCZLCDKEcJBWF7IKgaI5Y7+y
rAZukGyP7ZF+WvktHI8Mx92m6gX43GcHlCHNawXzp7qCTd/97IMQ4S71gzPvJ/y+8TW4wJb05i+c
+xILgLemz/bB0KL1Pb5Jd14/4KNeYw44NYK7qyEDkcvSml8gOGiC83SDHAqplQuK8tWT/N/lMDUg
PR9xbCfEYwFSbFWHQXKkElgaEr3klWFz7b58oCmfCVoEFOqOuhRyX9BYZ4qmif2WBnxc+smEfrlv
s8iuTmCdSt1w3KDqNpueVQHTIsFVVtpDFg3RhDeIgDKfQvuLFZNcnE8zdRu8Gxc6XwfZ7fEyn9cZ
/Nof7Z7Kull/ifyk0iYYeNPHeW1Ovf4Msg0Q1fdu7yh1OuuTP0JmODZdagHjMeT9ARo6m6mhN/Jj
HE+c5Rc73kHW+p+lKJAdoV4ez6iazn5iLKEW9+IhOi8S6hFCgEImMZ3evLEzDpVIHzAHAYbNrs3y
psBMDqsANrJlZYBnxg/+tCkZygZlXBKIH9+p4mPZzrX/5WnA3wmzowsiPEGBXWaEM+XL/3+Ukudp
Dz6fojRwKNqzLSydL230IDuSDQJCH9yFlEDskZ46v+43dPIltzplQxB9qRAlsL79QH9XDdbUU08a
IJnxv/WbQLVG5Qqw2+kNih/h7S15S87bAPbRtPUuflZeqmbgBbachyb+c94tPTwX1KgxTJ2wt+QT
MBaJXK1cAGRDUErG46XYRcq/th7Me1PvQwvGGeHpUH9ngU9Sw9+ZW/GRjLRyWmVIT9+HLMviWbmu
Bnf02CJZ373bI8wHqA4j3eTqJnkhtrySIVhiGYm+DWdiXmuT0FwuG1urgkns/O34opSanaq8tq93
a9WyOpvNFrONCTiHBZ7p1WOexp+hcZt+6A/gkTwTmqBzSZLL6eMy9UqjOoPrwuHiserRAfX1ouhS
YKpbXo2oYvP6C+Gxnrcw7Voz5BC3bcWKFZGfMChwQLShFgUKEHqZ/WtvShrn1/rgV+GFSkSqyVdu
xxZhElc3X9b8rCgER/iaQZrafCXvUCFOvkA//h5ByoT8RZFdYc863TUVlqfhMPrDC1r/EdOjJy00
r5o+VLZNSTBXfRKDF0s1hx/GIj0YxVFaJlW3NzCc3wDvFsrx9+EDPFTZATNRs84xc0HQOHALaSp3
tIpcD9R6dWhEdXE2Ef1yxwr246che/ARz38ljhQ/9tgSGQmZ5zKCTvKQwUvZqCp0x+d2dWPhgvCU
yFt6ek3qEO49/M6tf+dD/IIEX++FcscuI9tMHws4KFi/BFdNWRNu7Wz93cgz4fvWJhDUTkTMz0Tk
twzTH+97Dl6Ssb5cmhTVyHF8uANVFQHOkt4YuYqUYypMsCey4eBZlii8clHxwxzAb6oRWPg9YiLW
DN67wBbyMvdmhOBOnjJnMCDtNLm0AFU8bgrXcoSXu1xISpJC/TcxmLqLVePU3fvj3kd+HM1tZ+Cu
7HzC+ALBEoZ+Y63/S6uBMm+ZSj+TMeG+zsU1ddgYZVgjWLyieZ4LwDsCdBLryOYM2hRA/dJvXVZu
O2PPjXc0SDYYBN2epkJhmsB9oE+x1pESNambeJK4RqwYtkEu+0jRKRYRPbJtLeH9KcIOtrnibl2V
8ekcNxq/OjZLmpM6UhfF/07tB/vg1kdtt3Wrf4yYnx9KcLh5XPPVfWc7WaKXBGrRKFF4Ik0c4SVO
S9XBX6YTsINCsATfial2k/pLCSSr35h5G9H87amMjEy5rhDILsyWEbd0KRv62Y1qin3f6YFANtRp
cXKCu+S7npHkbWpzBKycWjkmXy38eJ71QVR67TYvKyaMO8t6MPC4xA9K0hjivK+uUEGMeqK//Xyk
jF/ryIbZp9MtWyHYwVXJejinFbMY3prxzPFy2u+OQ/WOAGbbCv87HRNA1byHR2XHRni0SbmY7Dz/
vRrYpf78SESBjJju39/ZTh/P34/g8VqBv+pnVy0i4+/HLYY2aaqHPknd5dS1ps7bqDD3f0LbBo7p
A2PFpIdbswPcqmXAfKi3I4jk53PWZ/4G8IS+Hh/j4O2rxH6yesAyCvn5sCNxiOy/zhoyHK5oWrKJ
KYJJWGZmgFGokGyZem3s+/Go2E6A5ScqNla2HVeqqerN5UJlxwzw2KJQD/IToO0wiax2s3hN2wJ9
lxMycci3jIV0l/uZtF6Va1mnO6bOv1C1BEaVVz8DAoRwvyrjOMQZg2bKvxA0oMCRcM9YwLdo6tmS
w34hDssnf2WLETerHWYR5gSkAnDAHPEP/1v8VE2pJNLFVahjyxVRwAWCrzGf2RXKPvo72owFEJfR
xMGokI86ltKzW2JiSE54YXtc5YNp4cxaAEkUXZxYObQdjhLPEPuPZucHIsLYHWncPYetzCbNKSXP
ULw7iGJb6r48OzFNOyzQEGTZXy64Jp4NrOVl+owjVTD2keUHFDFr0g2CK+CnTwjJj8UAE5DLLgMf
cnL7TT+zZ8nzo+CBkMvNFkScxTEhUcnw+J/fKwI85YnhlOBRWBBTPokjqMQxXqWJh641c+LUVnaW
1xLDG76zLQKYbo/P6v51pSIKto7McUprFPxXfHpfeWJcPpw/OXydpVbyTwdXaGHe2BVvi9pBm2Ck
jgo0aHvqd/GSaF8FIWFjjMW5bO2tgBPrIv6sDOLbISvVASq03q/IvFEDw5um7+Gb1GovsOwcI14e
WI29A7l/2vHfWOjTUeLGxU1/cKxx+2pAlJfC2jtQj6s3xuo15T0cWn+Fn7ykDarC7S4igpUWy7jX
Bl/PpOxe1fmAM+vyx+qi3lAin5Y1ROKKRUa0YMDgtmtN96OPjB7EkFsk4jIP/3V1AMw67Sc5OP/K
c00mZFWO4vHwuPkZBnN7Ckv5T7Rl+UK4BOztJvERdudhgKBk464U2YeUh5LfZADMZ8zgEmBMtaQO
Xkn2Yy2/hpkdfxAZMonTVun2toroYIAm94kwy7LHAhFH+qQEpEqsjGASnDFflG8ddD67b6tu+cqQ
60D6Isv8h9yKE/YKBdAPRHNtlg8CQeHuS5fIINJVPnCeBT63U3jyNCWMiNLocEFXapQTo2bzQ8Cn
bMFURKfJcbQKGo7E3WfRfwq0fdiVPK1G5XNKdybtZBZcOnY1+RoVC+ZIBgsp70yij8ST5kf4swpZ
e7EiwDs+QBZKAJynj89J7FjiwKP3CMqX5TVD3jUvJwQNnSIXiMHilZaw3s5n9vHsO30cXuTmheFX
2JkEPP2eOVV9GenR+YL4T8lmis0OFmiw0to8pL9KMJqes42Sx5gH27Z/DyoyQANCnFY7+28khyhQ
CbEuvyAttv997zy8RxED1Yzl+KiuzE0nOb3dWMCSDOvD/amQs+kEhQByVunObTh8UnymVuphXPcR
aDYlQervWlCoX1FI2kXu1miAiYN97a5Rg5Y/I0CK0uF0/rLGz/XQ2ud9uSHwPgK8RlY/pqHCuBH7
2/aVBBXRF8aXlkluvHSLw9V8Jvn98wrg1J+q/BRmjelk2JkVz0rPEklEcPJ4DoYL2X/uAVtQMCJu
if54iolu1BP18dP3GZdR9PoKYV5kwvdKx2BOwbuSODF0csanC6JiifvH3W8TyFB1BbZsX9fdYGsQ
tJK1M4PT+DZ0loqJmcjiuq2Z7Ik8LtBfIZFqeIsmPnYqmimWdF7sG02lDu+PvSsDEslXoKm3LqNm
qhDME5qx1+nQHUUsDvtuDboZuswZ9ngSVL1+jM5pMkytSNFxlKq+fsiyV3eCXZzZx8XfHlu5/rsA
NFEGLC3b24FOPH987e5Wt789fgNDmOPTww/rZzoHY5wpVI5yO15OBGIi7c7VqwxYRpAE1RA2pg38
8hjuZY3bVSDQqaALBpGDJLqF+nu3zEGWzEGd4nZCO1GsnEg2qWyVyJ3dD6Dk4AtU/PtyXo/HPBUt
7JN7ICLJsu/XDYcDbamzsh09JAoglWYklmE03B1h4vBWoK7Qah07fItweHXBPuiZRHDWljOa/Lip
aU2OegaH7dhE1aHlp9rdMqodlolp713yQBwrLWlqLkCgvHK5Seqd3UUV17NO7FZY8VQtfxC3PBPk
f5R2oAI54bIY3VciTXseL+jp16jfPg0dFZa5/P+n1nNeE/hypJdJhhqHwkUEhFvh/FXxOksbyst8
5lScq2GL6IAQRNU94kyLu2nHiXJ6oDWx/xnhuHvA40vYia+wiYb+cm1a5zZOabDwr8CpK+p/nypw
cPOshkTtY8GKAXC7l55Jr4/l3W2u9XZMoFNzgb8HtNXhWoYWW0VOZtl0HTK/R64NigUF0aYUCTTz
yvp10cXKY0tekbQdq5lmHmtE7+bug+JOyDfYoF3CIrF8wcadUfiBZr6tuOvj1FZe4r5lJRoI8GyP
WnUHX2CSDsP/ivaTBVgm16FEHlb0CfrKAzTO7azgSP9rD/oom8COktpXDjo/ahHLq2IjGTfAGzUA
X/ps4fYSQlDzZWBxA2cRiofKhOsijRT4OEy4TEdeWnOob4o+PBZnIeE4lUTFjKr7fQA0adEcUtOT
K/ThgeqW3ybpsnyy6moEyHmCbS5t627yx4UQ2VFcxcJ+XNuCLre+wLsJoqvUFII4Jos6QKlB4SSi
mr0Ci4x3KcSC0DWPwmhqgcSzz8wxuswyC7okWpFgedma5NkWvdZxTAHN/zWEL3XvM4rtyblBLXei
FSVVRfzqC08/1k/kAR1RyR6sXu6b9ILRMLbmgILiFkeXmkOzVVDJ5xulcnFj2LhUJw9L+zDBJJje
mcmcb28IZyuk54pkugSFHT4Hg2ftnHo9EZTFE9N9oQ/Y312NQStrvJ5NSmKwwx0NIunEk/ifN30W
+PtPH9dCGmGdM6WQyQyb3py3SyKB1dSMx/wEB3NkdkIzmwE3icuG6v4BRaQUGa6pIiM9IOYYLTV8
E8RjLRwyMj0n68zXgzWoqoMyrjP2W1pee56sPTsY/MrjQ6yfl5XoA+gnb23xmKaP7W3Gnb0Ccnt8
0PC+scCmfiErn1PsOKnTsAhxbDIqd9nudC5hGjdebaJNwn7/0tj3L2+a8wzdJApGc5hm6ju66SIq
c/lB0TK2EUf9zuNLcVOG9qhw6sivPkh6MoKwoUldX8Ug9oBhSq7GlziQskl7Da+SyjwDuheYsJ9J
r9fgvkBmkWGPZ4J2ZDUKmCYzTJ5UI/aEoVBaoS+ivbY1MQlOikzbu+jJXryw9ESKA1NpjgeiGQRD
EanHBaN6vuZBW64O02/q0egTfQIXBjCF4Zf+rXrJOs/Je9CFgKPjZk6bw3LXG6SZr5Lge7J5IkiH
8kYQKXhtSZ97zdW2Kb4mWPbJ9eO4XTt7ck+Bx+XXSOmvnlh3Lb6h80vrOIwQkxvgO+zNgvDWLEkt
nM270YN9O9RRj09burnBxYHb9rlU6jtT5obE6fLdzADurhILFti5DKOTrmVJfMLSASmYf2aTJ2JI
HhLMVd9hMwg+921G24jTOCAq7zhTzEdeOaik0fIyx42OreC+TliQ8FHFGtmLGiI6nI95PPPiWKsX
8b1SNnV0zAk/HI4Xoo/VWSkzKp0zcjmZ33zWRxRqqfSFi2nc4byrAzeojlvZihBr5hD2R9FzyfVT
iOtQwm3PsxWMx7wn4MBp6dxPaPgFXK1V/oGfW4aeUqW8r/cFjgtcPOcubF4oclX5+z00FhL8E7bT
ZZmN7bwtYkgyCNCMCwZGdO7Oea3A/Az4yZULSSCXf4TOiZsFivcxG18OZaofnCZ2OOA7Fak5VJ+k
+bajqdzXN+NmIgSEi0jIIcIhMtOUJnDTLZS87xz+QDeUoI7aoomTWjJtuVYiYdG9U0ipcDlKq5Tc
uLbVjusw930PwrPhY4qpp9oCpbLJJeVFxaeAEqowvH5wDQlEtNy9Fndt3gpnwBZqnqw0+cTxwO2n
9D+8eg5dA1NYxLAxEI8JoLxNaqJZw9s1NruAatdizX87GYKVjyCa3qQwy6FYbTBxfF35bz4nvNP1
eueL/dzDkiGefg3IVtpCuGaS77N1VpTII8cSW9FG/sho0OnChZUTDGKF5POC6DXBzq7aI80Dw5Vh
5QJaHvd6GtL8v1/RSQ3udLOjbiUdOiDR99YC2bMR+ruML8oFVFzjY2RdS9j9gbWk4+x0ayvRJYMx
7r42QXN7BFX3ijofirmpEMnGMM4AbSkW3tPvIL+v8zh826rhQBeimvHatBA2iZWpWKim0aDblcX0
5R53bENtA7M4RwO1hwxJZ9CB5gAOZ+SuMJQe/62FWTEUVIeh3b8TNFnFzri/ayr7mJg+kwUmxtBR
3GP6SlA/YbOnEWHL9UyRB54MtewxNyWzHzmN151JhH5vtl5ku5XwynosDUTWyISHR1JKgXy2UxoJ
govVg6+JcBaPnlUpvSNVc2TWiuBcMeeSLuCRVHmjomvz+UkRO5dvJ7HCXqN4kUGOMXI0uEYh6FbF
ItRb+yXZSYZJ/y/Qd1fwdHLdBg+PluUHz6EQlzSmE9tKwTnhwmoek7JIZOw+dXveGUmGjXN2AEUQ
DUNpmuQ+WYyVgTzVeZHtHPjgG0/OyvUaSuHXb3wmZNfqWKPPd9Gq2PGw6hMw/s4mL2DzPbCYyDQ9
Pck2KLcew1bqZ4mz8xo61TtF98TsnQjpa8eKwRRSMVWIKCKWpX/Lo3ggplOqFZkZ8LTyrjLD96un
pnbSYMrFyv/Q8kmCUAft0oa8FPKsmSUlCRKuVmN7+dr96HaiAva5t/a7JcQqvwBGEsckNFkdq/TC
3Ekwl4dt8I0u61wrAo7Oglwo0Vs+krtwuiQSMWhT+UXEl54HIeEalcU1/IggGs1bK7HDWKZikxfL
O8syUmDqBKshAeEcJPUOK6vNT+quAaUEyUz69EzkNM+QsWWYO2+O3xhhtn1ksuw5pO1rQsNcWu1t
cglrdjp1f/qWAHnsB0/kQEs28xVCkphbhpVXRQJImlb3MiMLlXI5qdYlj3XgT5gmfllXkFuOQNjH
ezxoCyvtACmh7xXKNgNk+upPd7h0+AoZ1ejcRm8oGpoR8C1YvXTppkKJU4W2wUQBs4pREGpXDfr3
Vi3YPBL1W8DFIMjERO9db0z4xH8jiF3RK2qSEFoLLh7Ja/ZMJ462gWdSM/qMuIR/LwwUi4ul0+AW
jI/rOIv+V75WA3S73mX/r6QMATYcW8HMDjK+45Mkwyh3hjrNT+ccnv/E6M3340B3AtrYaZg9u1v+
7Wgglv85YXbY4yMAFm8Ypv9tpb/154sEvD8IjbTiKKNetsKI+1YGr2LfzcN0/dURr5qDBlI3IQvd
ajDqp7z7TVX5M9swNXs6DyfYTBQW2z/eZw8yqArt2C35fjV34tIP+/nGqFAQq7NsmATjXXGqaTtZ
1YyzprdtjAthLZ95hqdWYDyPeAy/cwM2bkXPHpill/Os3SXAD0NEW7kPUi/OZ0vn8ZTZFW2A1lPX
rFi4+kGTZAJPYj8MwfKsK6YGh4l4vWMOalI2RLpnaBWbpn+b7rqNMy3DaOH/qAasH3uGyMXy6jCK
uMwplE3EfNznfJODKLh4UhWX+4VzG8njw58oKzfvnLOZwIDNLzH34sSemFTdfpEV9EVp6fghgQUm
UoFXx27ohfnYUU6Pf9wo7E91JCu1hFPfkNNgY342h/w2zYp7MNhVl6KW49UqanVDLfw6mWLXwM5v
fxzWjkfYsDBlyLOh+Akpdqtq5YifH6aTljsUocngynHWT1JfNYIWtYi8oSXT3xqPRGxHRZuB0lpf
wvpQv1drFZHNVU55IwmtXQ88OE8IWw3e86EmlKJMpPG7Vs5WC47Gm5RyrNzBKj9ltpyjAVvgHa/5
jXZFZOPP2lWy6w5WtcamJxJF2d1PzUwUgqThNPNc9SU09LaXF+YaPFd43Qip0tJFL/gHxHwJ6AZn
K89IOTzCp5hHUr0R8/71qddfUF6BXoGEzgYLbRikT5m9dYSQ8rQYA5IfDSKZrTggJ/JJc1iXFAN7
9e6PwQrXjqni71vTQkcgyNUE95Q9RdLPcBYP6AyKIxd0OlaNv/NHuujEwVbMvgDxyp6xLG8Z613W
zVOI75OP+mVof8hEnvcueuUIrW+tzfNEf+lJ5eNi2rK5lGW9i7DQY5ef3GLjvHrxarv14xOIfzBR
m0CnNgVixcuYkJOijToTguF+iezns5OxPINjasjWsEqinkakC6hjErvxqi2nnUUCAi6jEOLFfEKd
qc9MHROaQn7VXB77ivDRns15Vg5jciWCJQE5QoBL1tmiAkhZ7ox3idHmfMrnGf+0FW5kDlFz3CiI
xiOxVlsunnjw/kKDWs/SP0nA3c7+LskUPkzXUxSEXD9jurGmmgKOMBqVGUzM40zX8dDzGBBwZnOH
JO6FeF33dxc2bBrbvzGH5VOwqVc76qkHEp/hU/A0fFtV/y3OL0/gkC0Ywc0QgYCz8D+dRELfUdSB
J8mgIC/hbyUP42JTU4t7LjbQ1pL9aHO2HXqKTtuRXzaR7wnqtqm4p7B7ct7mM35K4gI2nkVRV1QM
8J4RBcdCfGQd3UC9jsoTohmMo0T01lyln/PgAbbMneb4Abx8I98YgMkAiaJhDeJhGgi3QE4JLZBL
NEOVciocsS1HUbVfGJyAJNNG7JVQ2rhA/CqytyHeOYiVLFY+AC14DQf4/WC+XWF2RhqxqBzPWVM6
3NC31tW4+RUOOyPH4YZBeNUeAbblTLZNw5GGerQPijuKjPh31lJnUoB1IjfZUB5cyV5CWP5x34Ay
frF+ust1ra2DJuNwiRK8vn3BLNIydNA4j37SO/yFUADT5SV08ctibQTI4Rz4YJCMGqBH3A8QLFC/
dWoAHm3dxwh/+7UVnxldpvFU+OXRd1CAHLR6XGuh2l4992FHoHJgsIanHkVUAOFiDbXPbOrQW0/j
Ib4rM4IfszxljBDkK3AN3EgxXXNha2A3WW2Qz7Kxi2x+VBO8k1RXyioh2BdvgnvXYx5KC5m3mEZY
h7pr/ppPge5mdvEeUibuj/QU/tH7+pj4jy3ueaX6K4xYGoPBdg68KxKfDzQ1+nmg4yP322QaQRIL
RdK7IBvYUfDI9kWKONeWQWVWwBxXfYWvOT6maoKFXlzDhrdP5XGugHTVqWYEr11zotZ14b0Wlnl+
B4h0XQeKQ5pvn8bzbq+p1IY5tlWvYM/9csIF69or/jegKJ7068OR9cgar7Eue17cTEMJMHexAk4l
GSZD+1OK/vQoUjtQQ6e5g4tygBYLuFC4C/h4O3ztCZwe5gDeGK4WUzFLA8/y/LEq38RADdVzH5Am
DCaCluRHv31/yBgTr239pwG3cnNBl2rH9UpRiMf91RSWdmu0C/q0P9BscMvuF83kx3FerlaH8ZEe
7VonnNkLb6DuzpIkWP5ueIJaDjjEzV6G7W1oP336CGWUKGVxXcq7wYVILBxXQ13HPNq/HmVc82Qd
XxrEZ4Qeia3+LDW5QLJcVw5f5t0i9TEJphH6FeOGHBQQQbye2ObR9I/f7fjewhHdL0Q4LzhkQy3H
sgAk0Rf1rnUmXn2AfWGLDp9sIVkhZfvtYHitPxA5/wFltXSZyfNq0Ntu7mmrLZR1DYrFxx76Om3C
4ZRYb6UlFNVVA/HtUj32y85B9Q5WeoaOwAapcS8/WWTgYb9QZW9AltgD+3e2kva7d1J0edQN07eA
qXADDYJCVEWIcXCPXbmHIdyIMqF6fIJ3Rb4qiZNGYbuMF2/tw8+fUccNRCl6p/inoLh+3aZESWE2
Hce5aRzndbRAPlJkuCuT6H6f+CXicKEpJBYsC6lJzuSRT0RbqgWvJE9ZteQ2FxX4JDnEbVIbiwVr
rda27R8cgvdVQ/nZHG/KHcYf/43RKWmWHVSa5jV86Bh0NcNjACC8qRwpdFPRvN/2jMpyAAhK9Ze8
F4r3ZNqvcZ8YblwmFd0utPkvoiPTi5XAFsPrK3MSHKCYc2PHroWYaqkay0zgcr/PkKg6ghN35HKj
/KZJEUBHqCuEAtZoO6AnJPgmgeatT4z4yoPCP7mVQW/1sWamN7tvlkU+j4d33qOvUuBhMh0Tg1jT
1GdxzKaLmPwzV8/ug0O4cXQ9aGhN1ERsrG42Ol/hwX2yXLZj7gchpjlXQ/casXSiAUpY4JAzRFPx
uz/spVAncJ1+Fcm3WNNwabKmQt2bDsNAO7Gr2qe8Z8ocqM+C/RmNPvcOIiOV1h1g6PR3O4TgqkQx
mD4j+d8CPzDEolfgmo1yVXY56rVqc7vKzIl91HmJtbY/lQu6qhVqidt9cEfSxMNa1LvPY3G2NBpk
Cf/foVskzcW3k4I2T8PAqbsRuwVvTXL5PsLc7NWSlXqQ5MXY1QADBYbz9mMMhD05Sgc+AaaIjDoT
o5ECZqbVxompGCcBXzJ9o9H2GFowd7BSDbmEm7mpAPqnvSkvz7/eofBjyJlXXlKexLSbMrteD8V4
Ts/5SES4eeAiWgxXR4/d7fUVOSR8GBI3uLtUfTAI02VWgu7fd+GaPUiXnVefitCXEjXFyZjodSOv
54T6KZFOywO6CiMWlt+8tciakimJom0KmljGZ78d8bpgrAGeE6cAnURj0TroA+OHfFJmsJrPQadm
xiOR8wChgKaLzJM3NJNCbSKjiBMGTmeIC+6+wDhJQpN4pfqIG5LQ7QoX1vqjUsSCr1pJ5Um1soQn
/fWXA8KC9pNzYBqE1LwlfKx+j8XuyAKHBrkhcD993Vv/tARRCexvjzTVvh779RJhPCg29ETaatHR
k+yDNoeRlBKgUwLnV2WlCYBrcSI8AtcuI80/ZYkA40sxefGKQz1eILV5/EOv8NW8sy3NVJrGCU7u
Knp+ZAeFBFXISe1d2+R+jVpoDf705p8iIwds8JHBPZAP0D5Wnd+wBByauIT/dnbdiy1ZNQ0I7Rb2
Izn3IcTGeqCbJFp084CZ3cOopCgVtGAMMzNr3gUzzMF2/JFaZ8dfRsVw4kHjOFVz92qkJcHhiLtV
hq0OzC66OmhsN8nSDdaJbfkk8FFYgJ/IjdWdq1aHQNG3CwdB0hKFJFUvi8XYumfhknx4giPfkuIb
LN/rxZ53RVxPPy7wK65COr06ielWqsicoZIigOjdM3TlNVZWi8HthXDvpYTyoup+Z4eQ25bpeLY3
BYJlnNpZI9Gq3gc8rb2I5tA3bzdoWGqpK9yi09pF8LzxPbgGgOlCD6N2uAwyJSJ7C9P8akJBAMiL
PoR2Z4sTA3MFEk+WP0JuDH5QCwcA9WSM6M9t8cBHFehEVdYTGASgRp8QNDOjcndFgHP0OIHMoTn6
nI7b14f2JRdEFf6LSwkrQle8mPb98eSD6b41LCiONsc5fOL+ZoO77bvLh+YqgK21s10+Sp+6oHxA
NeLgFLITb959zaNHuulhNstAm2YGq5fCfxShjrYrH5Ak2EhaROCWbXQoX9CVOLfrGpUKUr2TzEFm
SbHC0ore5HLZ/lS8Ogi53uenh8+nBkKGKgu2JG9NjYAplmqR1WuWOI14qzr6J/Vx57S2GLXrnCog
89EW8YjP5XXDaADojMP+BT0rk+UtNGsLP1OR+Lv2F9ATb9uvx7agEDZjPf5I01osdeLUmb+cxJft
322AWUFQBmR4HPWmzuLo2rP6GCQl1H1zSb+IGNvTdY7wBDNLE1Ro8jFruh2TxR/xmVBNS2OaIv++
NhkgJXrms3dnpsg2WW/TtVHtOGRap/NgyIIZis/VKAvwNnpdlTNv9MP23s0ozD8Ik2GsZ49nq7fM
Pc8eEk3UYD4g56ybsZlF/oI9UWT5GSI/x8+PP/cIgne42EA7Ks6K8N5OA4ODF+R51ajNieFAkZ0j
2yn8PvQB4GNnzcaQ5FKpuYIMcjVCRFTvpgjMQRY97k8B1R24ABXrIE0O8nY4w+/1MOimhXg3LH8V
I7WPzLzWNzdVRnXW7FCinT5jxk7vl/yIpN/SrV+TCojvfAEALVceooM7oyvx8XOVvznEVyxSoJns
TZlre7wabF+956us9Ty58vNE9AOfp2cCtXHomlXUSvl6Lti8/H2kRd+Xpt1TLToT94ac1bMEg9xg
SB36W56zfOsQTY5b3lGmvfinY1ChPdPoje0sYEoBnM32OSHUm4sohw5S9PjJ2ONvZSVq3BOlSaH1
lIHzIybayFq7prenpo9M0cn8xmPgQKVb4jX11jcP3Ty2wASRls2A0k322lMNmtBFAg6/hu5qIYGe
tVHZ0wKshhgr1TvbUseX5RiIaKNCmovGrPBUgDfSneEiRG8ZedPXm12JLCfrO54rpl27gDwnDEsg
h+KrOJoOGuPqmiehYW/AMdD2TmwQLEwwodRSuU8WMeHxArFxrTppQfaQY5lwNQF6A2F4IsLkyMOR
yVHWuNRBG0mmZxTzvg20zV1YrTThR7O5iTGRxJioTy8o7jD4Lz3m8OIqu849p1/dBQAGq3bFLbKB
IKMLshM24dg1mEgmImkdVWeWHz8s+yUEPDCwo+Rt2Sr+IQs2WKMWG002nltnfoTyNRtwApkYAYu3
wvr/BdiQB5ysmJ7V96JcrwyjxSCAkOnicWMF1rXUrI6UzNVy6NgG1dH137mF3wVl/7xSIucD6kjp
hbHrZIexTDBEABn7yn73tdxGhQM/rIJPw3qiQAcvaeipMpjWLTMzVSUk3xjwn8B5l56S+TWBK+l5
QP1yt4q+3lpJtHnSwcKtfb1Sa1rDQvI1cT2hGnimrj7z6XcQSq9Dgj8HU7PmsDZ2Q/ZX3182xKoG
8h2QBjtOw+M3b/eJ+DfQ1w0pF9SqkKu6YGwxutMChfCGm3+Y7sfZJPUm4bwtaUA9mhH8VzyefHbx
hVO7VIWb//OVlyZYDIod5JYEpxYv5249pbVAYprUXeIMNsNwktF+DA7BI/symxTMAzqW/35hFhn/
OeiNE5MzLozXOagRX54PoZo5Lqq8iKm15tdQm+hw0GALWayofjBSrXPhY3Bys3KhCoHEdmQVzVmj
QQDi03fSRJz21Us3owsRnjZI81DWFMoaUuITmhd9K+Uvb+I3Ef/Xxfnvup7cF0kRQYS0aY3jrtaG
pSGChOCwoxzBXvHLZa9nVQGR16hY14gcdaYHf6QKu0r3sJMkWreE5XcN7IL2eQx+SXk1zIdaydpi
HCipntQ89NhE87P+zw/MDcU786Xxn/Ysy8AiKXr84bUCi24srS+TYLJEGuG+pToW1dsQV/nL9gfv
pRj4FqEUwX4ltU2r9ajgY+oQbeZ4TYXDTjWkb8KUyKZWfHg/mxAXWw5tj2kQoZ2EeY9tw7IgFrsx
z+AjNjYSQFe4NVt7fRw1f6Ss2tvI/9OTENbOXofgqcWHvs2Xf2K++W8Uz1Zuh4lnJiwq4wd1mMj2
d6d0SUybLbfEWnqpyi5r7Ux6gat5Iwel0qNNkB5pyl8RLiNJah//j0m3E+SmQZ02k1fkfC+3jUc7
CRBqvjt0ovp+C+rr8HK40xtIDuBgAqocKlvHLaBU2vnslV+9khr3phXJhMYuXUdu4PnsYn4zKh7O
ixQ/4RoT59zxhOCsPplo2sYoZm3KyKSRSd78NZjzDc+gxDjmPI23zPWlYv73TKGRujIGSQBvNbjH
rrh9An3iWGOkwCCzw00sSlCfGSQnEChJLDWkrOAVMUNXJJeU0VGpY4XLf7pjb5BZrDUDSFPMZrYA
/emqLMd5ww0HJK01mOQheHXJRIDGuyEoENiGlbH4YptM5bGfY+FwurXLAHG5Rl9qPW0nFMJnGe/b
IFijm4BokEAT7lB5PPRfx0pdU+7ere8lDVMQ2YxkCwfMWW84kj5e8i2mnXZL+e5DPCzHyE6cFy80
//3CXoPh9HEhRXWv455Q4s1+TLACapci1VWIiW+nAq5mHivp14/3ayXFEBujaIQIAuJM7Rw9FueG
NHJ/w4QE9+w8F2K7LrMZeXO5j9uT54MBkMhjB43qSWFp7SWZJ6pB+9Bfu+fXzZkpoqXZtQWhVSmF
mqfB/skXS2pPmzC5tdou2C+3/dtdNn3fNVpSMkY45w3naX6xEwKcbJ/hpNGTovPPE1/UVevO1rIP
8KuiUgwGyoGdayhVlAt8VeR4wwwneAJLhyCZWB03b28DMUL2Yz0F3zO3IcTHymtbh4tThlkZFdSe
wbWvoqm0Y08wY/zh/UeIiS+yq+Vuu/IX/mGKv22E+V6KzCcWtgUEIT13a3bqKjbKS/KLI2FVEeg0
7av7FPrRekloPEbUf+05w9Sp5WXsybrJ4SRZn0nkjMLu+aDAxApqdJAT2XiIK6WcxRpC54H0B9qL
vS3rPrjgFj0pUxr7Pl59uzKzgHpY55u3A9p44mXgdxZ095BDChX5JzEYdYgKpIqsdd//xp8CiUNP
AbVtQ0MEmtWoAlYjNS5MpTvVTb0lqRiPvOZKBZYRZmeMo2+B2eX1tNlVP4d24zrrSxzSxy0RcLY2
6qDWc0c2bqGGhOLoF6Pdbm0t28KhfYqrNAP+CCp6qCKxY94mpM/x65+h8XkHOs0x8My6KbArTc2M
e4heQW8xJHfjPdOwkfbC9BNDuOLyo+aRJD+dcgUFqDrG4XiEw6pbmyfpIJ7ifwWxv/YIp5P1Ejzl
8qHysekHjBkZ5fMa5PaYSLgAFd6stUoddGCKLL8gUNRus4WwucZTFwmoJLtr22CXV7J7G2nC/mKS
TlDpa5LFMsIp+kJbHLH+fAIdBR6iU9yusALhKDezRdMfz2AnVpzkcKzKwYXNtGMUZjCeqP5PAPqo
fP8VpuN0s2cQ991oOplvGm+ZBrPYzIkWq2rzbqim+FCDqzcgAetLJ+m6pthDsJXatfj6MngXSiwi
EBXLK2D4O7TDjkwyI1uZPg+SJALEEXXi22iCN0AoxxJ1X6b9aJ/+qRglUAD/5mw/9BY2WQ0cX6xm
zTlexLFaVkWaLFOSyUNuioOS9SN+LOqoRz7GZpzFdJc9lLRK7kjSl+yOLe7bA66lMKixhFQM3FzT
uemUY5OXSy/CyaZMCxiGfZYR8+UolHghvO4DNj/80RzlyhlTXpT8Thy9eP0rMvwe7e0BciLvyzmB
T4A3h7ElmCYCwFlOR/l8muinwS63tPe7dqVINF3IjqdHrjoRqcHg/g+Zqe8kJ3XeXq70SAZ68mSZ
EQXxH9gAtrjMWnn89oS4OUnXcEotRE9HnLJ8gD1SKG5bBweLz4mGuv5RbgfAR4LNwttXX/Whamzt
zYBJW/pT2fbOh8m+Wzl1STRcmKIg4ngr4kaF4KiRtlg7RGotBS6ENvsrirMf/+TOhGhPSwlWBSN1
jpykTqikNAywALcXhOk+E8kiGAMSUPj8gRWHG5ogW5uqqea51OTC5vAu42AEJU9M1Y7g5cB/PPl9
4kJDuWENfINpdPzdX3QWrukVPRPP9nJ7tiUDBDRDRSj6MADqXHpqbNdhzYIOCSUQPt/+GcAIKO1f
m30Fjt5R4rYLmesyNTnnbtMAZyghBq5JfG/33AmvpcR+XQvVtsfXolVCCDu75pwX4f0HCCqEj3eZ
Chr4B6k4V/sSRifYv73wViDi8zhbyorGRYpWOHwajfRNas8IaxYAbIp9DOkXQQRGB/nq7rnwTV/8
jL2NYe9T85slSaR2gaxon62HCx6zXZbeSVF1q+6eQ/5h38Ovpwkl+OYh91Pu4J7TGXKG115arfY/
6fCuDqpzdt9a85w/R8z8fcMEoideEWdL7srZuFf7ni+xR0XPZ43zLBHvRLTsHo4c62YGZ4uXmD04
dRRJSXfeFGI7G6ruEadb/AB5vmIQAGVgtdA1aS4gvWb95FJq3Lcc0K/W+gIuqa7t2gpcEnWnwIyC
VsJ2Smg7vKOSag9UT5Tx2tgphjRD+rHkbUtej/6byKLhmGE7mDgbD48DZGcP5ZAy3B9CA6DvFdEy
GNLEbCEbg+TxJ48ksliCJ2ZqKrrxtcGM+M1fWnyi/rZhuoTyVsmDVVfdVLVqtTR6Me/lLbBe0swV
/61QbKxqR2tVooHfJylf4F0LTwx3WyEnJPtArIfNCwESnTYmxxGUwycHpapv2XpszR90B2DP8kMh
fLeCpt6FU1m6t/e8ypaZ9Rdmfa77NNEztMFEmeUMG9fN5zFjdPtQvVpnFa5NHNs/7XskTXsLik/l
DRftb/l4oilNHOL1zdPVa2eGwvYHSCp5q/dAb0vs5OwS8FqN+EXOvw/Gu2L1pEscyf9heJ+DYQnK
S5cxHv7MSIBP2RTe0PHUsMvqlxQp5xd1+HjjmVP88iJTb3nxXf981Wb5bs3EzJoRSwkAcHhShONC
NohQczZMNkOHBui6WUFHaaUAyOj3NL4AKf2T3rsnqu9xiOi+/2AW/dJQ37UvV3YeWshOHD7NGOoF
GgNgnWgYVqB89jmgD0lKqtcCfoqi8Pa66t2McorrJ/kL1SBGknWq0lEbmqQbvY7EVnvfQN4TGvgW
v7dS3ELDVk8UtezUk8LiXD79SjsElIPyPWxJLUG1M7U1hTY9v5iOxIkhMO9zUDhqjTmMnnnY1WyG
Eai+krpa94e5sDi8IgD+MC8K0VtQrYVU04dUNfsfGVo+f68O1wIqCZf39CMiWe5EoVSAGSOVZ8Qr
wm5iRPBwRuGf7zsUTBLisrzqzX6IknQ58fwEALnr0qXEmFOpgdj7mjxQYLPhc+BWqGu5ZBgxFX9c
bPUCOdlgaBZIzP9AIaENWsphL0Psa0I7m8aXYwDrzwLBPQSoT3pz43tTUCfSF7Oh6bd8assPM+DZ
QaOety5UEmX4lMYInH7lpy8GkWNrzV0oyZxXqWbGKxB7HZl03YPYBk+1w+VcRguEL9JqSiNEJIFU
jhcTi1mJorX/xLy7D6GUv6yQ6aHWgGZd6LIdtbIkalQgjZxepi725kvDJ+VnbjadDa1un6ucyX/G
syO84KSpM27qOHXmF5HgO0E+k7Zphj9L2WmF19qPu31We3bRBieyZnvbMj8jDXmfeqUOTRN/MYFd
qTo7bQT5k1Dz6m1aWU0l3wbN6I2m7Sano2AfSjKYj1d2rJIEA7pEnBtHWBSCdnsMjO2SlO1vWrdr
DEi0GSGb5wjY6ldNU6nYvO8a77URW8mFXCn0HsX0wqpdEUvOWBmrJRWeXQSLPlN5KydoVJNaVr+U
K7DrBcqOz75f2BBvKeUWDH2h7x2J1wwqWqWju4yjiL2N9TrVWDsMmm04CtJE7svXJYtLSWvrXx/L
fLy5s+HDhCvVGNDd+XNLPb1QPMwn6umWxsLLP1e+0pxQMaTnnkB1xk4SW06C/YCB90cm3TOZwmeA
6GR9efdzR6HrRbRMg1WJGfs4dnpfbJy2SiHuHQJSQz9fFzFYnr2t0vQ7uC2ZKNeTAYJJof4Qeumw
Pn7Ky14N5vCcxCKoqovGDObVYlRxZbViBja0PDkJjIeElbJpM3xbHvLz4mgxIoHLuD4DRMIYM+44
zJ/kJAflHPOdOoVZaXU6cTwIjJa1hG4NTUK57VtXSRyOU8OS6PrRWpPntEWYop9Qzdm6IlKkjn+r
vVZ500FQUbt7wYDLcAOZCZUJ6bUHVWpPxwq8dKo2P4utmtFVXrkQ+w3K0ovkm/0xw1XZle3k0og2
0mWrzmoVZ7sWdLt6JRwQvNea0w1p2BoZI4yPcTG5YGoRAFvjfwYlZcRMHRm//e+SNi+3g8yub0+e
5cmIqYw0GDuP6++UEyt5xaoYVS1rqaZRb6rSUWZE5vwMEL/FH7L+RBvGycbCpQhsciPVBsBgRHJv
+3zfsUvT/bqanu0+fX5Fj3snT2Y3KOYib9DgCRRs6xXsAnAeVSvIhYuT3UeKqJ4BXgTJrbsKrxZV
A3M3/g8kh8E8QKlwufM1rX1aOvx+bR+DNonhJ0R1/n/3isTw0bJqy3pTzJrpXOhxct2w+Ta2a6KX
TguDmVU47hTlj/xLp4Cu/nGoQt63APHwZd2TfRv7l6vB/T8sqWUPhONIvwh99JYOvxYDb6zn31TA
IQNXGeIltbEs75yLkF2KWOblwizlk4oZK2DARgbnNDx7rONEhjOo1t6Hd82c8rM7imtmHKELt5BS
PjkwfOnUGCWVTBCAAbEs/HoKVsy1U+q7cV5XWMtt604aSG1cWAfkK37uijla4lvf8RFiSyAORNYS
CgOCaJFk8FTL78RsoG4jt5soFjPXc4Pc7zDu3RQufkPfjN9Joe/iiMsp5bFlFFWO8U/10U0mZrH9
olIN9UeayiImV69T41rBxKfk1GWodT/7zYYPcUO3En0JNe9CjiCC9J7DNGFDAu7fWAO8NNMbQuIU
/qFCGY1z+t63eM5imK52i6oBL8nEguC7fi2MFogbI4ByyiohYTH6v1TbyLiQnu4A9ugmuFWiym7c
OrzGLSJxi1e57DGWJKYlKV6dS5ymVetaQ6cuMBNdcI7kyv037csog89NDeDl7DtVaiITJf8sQ3PG
HlrN+yqPu1CuJQ9nLLM08R+c/7BTCsQJUzR1NpIxTL0z/6gfj6XlAbPMuCNrxVoyC75tciAr0wTs
vn9wJ8yMm1Jl/pYulbIHl2AbETFVhLD8awD78bFSSHVo5ZOVofoJJaI1hDqP4iiiYLreneQrpprj
nRjr0baSp0LI52drfYhUlJFXlRxNw3KMjyIkiE+Tn/fSaAxjRyQEH7oynXJR44g5xXh18411tl7X
hR9OTeeoNmla24e3ak8HI1uK2NfM1FpWeQ6YyIGhwR7vYJmH7i89WjMF11olqNlxLh1MqUluVy82
DMm/W9AtcVLeI7wzDkDLDmHuiEbrewlaDng+r+7ji2jwCb5pG/PoJ9OafiN5TQZd9lSAmKrksSwh
y+dT/yv4PuSFfaiayixIAAibgQaIgPNPDG9llewmqvWo60OUT8RLJGMJ3BUifh3QVt1E7muXrruk
q8bQUMM9BhgXPL27nQ3jeH1WHC3SHdIbk+lZEL8iyfA0Asdi8sFOpznYuqvEYgEgzUKXPL+cQs2i
zkLdz9xL8LyPiIwcnbT30jAPl+F3GgpAIb5eK2cSadiMGQc8u6V7IP1l5/LLBf4fNuiKyNUD2FkH
4KgEmDO6P9BMJvWtT7XWHveFS4Yr4rmEPmqG6N0MbQ42gYRRbxcllgafn+j6T4cMqNEv0Gd2VKAC
9qNMI/3fwURvGwcONKlb/R5iOHBf0wYkQNc3hHAaaSBopc2uUlK3pW76X95fHsjqb840Thqp6FL1
IRXgW82RbLWEBIpf1CNDkT3kpOeGvsg8/3SX+9sq1ry6BkDQbq725+IvRTu/8BR88U7ZH1gXFmbD
eSPyxut/nLv6Yre8PguXf/q4TCIq7hT2YPJpU2QRsHfdXzT0HbxvHYd5yQ/teBoMpko0o+P2Z93o
kvUlLF3bs3+x/FNVp95iZAhBZireqA4l8E6NuiUoqt8IApwlojDf5NsY9ysCKA0S2vZPrSzmfPRd
1umM1iKFiZf//3pxMzlARMJ+D7augHjM3IJrbffc6Subx/MH1BF1iuRPX7DIjxLbhzUmge3TJOi4
jigVHJtsEkesexEtFXO7z69A6HhZ7YZatlwE4jz7ZMa8f47IhYWE9R+JC/M6ULkwC0j7aSrF78w/
60fIwKLA0siOwHvScb6yI90nN5+GxGp1NKkeJfBQVUVI7KYnxtIZ88q6OZZPpO1EYGguyLdilzeo
GHD1gWTIT5QB6BdSPCN9MfCbF/SCrCWLeDaESv+R58eXdcSWhtDZBn3eFp+JLp4ZaqLmvas+lfFY
pZMxU1OSeggh6gyfeUYAOFlq1QF1NuJaqbRN0vEBUhU7XyrK7WzJfwTFQN0c5thRuoEqXBDogHLQ
q5xcEYrEEl09tSePAkDmmGdps3MdkeQ5ihskLLCHLmyFAGjjlfRQWYtgwtnhdwG4ga6AEwjBI/ov
JMr2RsnHDagLXA2tM3tNkTLrEfr0UESQJLDWsKt2AKdHbe8of7V7bNJl6tDqhYuiE0nTSNIfOD7o
BKe65kV/NAi7TAoLGQ8RZ0rfHQt+2e+ty/O9wY9a7PH8zvZYRJjwJ62g2upVfHISSFufZAyOEedO
Llb9LZYZOP+x6aFKZMC5Egbs1nkTp1WIMe81+BgpzTy3K1WUNfnjOeHY9JGU0Azo9/b357akgrTp
gMoQRI9Au3B5HAFQ6DTP8zD3U8I7IL/ppR2Hq5TyOVhof3d9fSamhINJfh3tk2NGM7iqsBjTqyET
0m/aA9UlH3RFUaZj0EX2r5MWOxh25MnCMCXrgHNVVEaHGoNUPzkA9znTGkdAmPiamxu6ZmctYBr+
g7YitaS6iAN89sCQz6ZS08rGOIV24Jf7yxNUezcuUTBcjjJzgn18O18zEz5lfh/d50TIenKWHxxa
6JETXxoF4V+eW7tRBB6HXUOtSddJo7Q7DxYL8ceVINRTD5V9eYDDcr9pRjFcWDNl0PM2yudbDQjS
guk4jvzqbQbG35tpf6fg1tjFSrgZO7iUhsS8mxekzZ/Sr+P16gHuFen2gbq6caosBPMIq5Pv/maB
t5OQDQZkuOeB431HwgCSoafTJgjeUwtkdsyP8m2M3wINdenpeuyy4HrFbjoNYM1NdpqecJt8CZ3W
G8HKkamx1sVZOcqp6dohv8ybSLS3thnFv75FyrvGGnqWsiIa3zuRLCMa++eVHPQgpV/AYU1nT7Jc
xeBh/7A65897p0r4GJF0s7v8VzkW1Wpyh9M7XCiG2zPXii0lH+Ur3y0aDlYOTsMpxMP0FOEpi3W2
NQrhp9Pll2VSHS7dJWdx0h1QqnrN0qw/sNqGuOVARDCkhvmAHCUaE6nILL9/Ca9jweQN0U5tKzzJ
D2XJaHdqXQsp1PX+qLM8aTSDiLZ01Bm8MATupxTT0s216aNRh8P6x6NaYit1dFGdhRRo3vIszjkj
C/FtU4TSuSma6Ngfhsp7g7cmOP6x1YihyH1R1nC6vJRL+P0KLdq/dtw65+Eu99tOIdO/4kX7wjms
AUTsm3EH1WIsNYCbQXHf9in/OQ4R+kSy+qeIfgVcNGPGPOTCTgOouHWTtIFgYXdYyvkC9qAs/mBt
i9uHVbaDNXKDCq+7silUptUix1hp7C+EwUzJVj9gdWpx6ble5onBrdrROxIYnspbBfHJq5XFr+7y
X+hfuCte/mdTNp0T0OwoYXvj76ZRImg27At7xN7mA+LEapJV6ZlbrjZ844sU7KAQ+MZPhEv7GLZm
G56fAgbNlaTmWMWenAeMW3x47wa1Gs0ay98SYROeoaC++77cupks22ikRdl5tzMlvhnVy0ArzjGG
v7gjIvmkVTGbJeS5THObSzkVu2cR5zQ0ydzi9EeZhK1P4gurwkDIfTHtQLhkm0K3aqxPx0SJ0WLp
dGeQsCFyxTN8Ul23CujnDcjvKbknN4H6kR/NsJyhAbGInX00/6msW6+gbcJEp9pQXg/AMuYCwSOd
gKtGIN1A8mMdHjTPTZbccHlufjHvCFa+pVtpcU4oi/KmJC+tgbUiA7u/xBiu6Dt7dge/y2mp+NKO
nvg1b8sv+/CxpKN2O2pNroNlu6VqShoCgskn55s72t/vNX9uuOnPxX03jjmpPYhCS37fXmDf0ibR
ZVTc8vWEBnTTVATKZrXL9ewarx8i/X8SLLN9qlyYVXcKfPheBDreNL41v44zaWdxZXqRbkPMi80D
d6JrxGO2MdCf8cl04vZRHSEREYt9kdYjZzmox4S9zanMTHPqSfjIuXEwURVz06Gk2b/lenuHlFWX
8BUoaTwnfqYeLwdpkw0ufm+vrRHilcXZR4EtovOhur3+A5TwH3hxlk/tCTDzsV7Nq5hqzrbaEN3i
Lm0RcNtnPaB2DlnUo9Nylkv6nm1H5fGIfB+7VWRIwnyVPfi4txPUESmuPHGqc/SUAXI3+PBTic99
itqNb05zEmYpGidK8/7YpsQU+WqIH/anlL27jSDz0HsTU0T6d1i/6F6R4NW+R27qWdhh60Y1veWT
0gVOnivanHwaaE+5rhOcGQ+GSWYznjQ8ZpyXRnokcReEdSq5x67BzBAW9Wcu9xwUouQ/RwK78kDE
KxDGWGIqXRFkwIQG+M7B8ARLrqWrSLFa0GBV6XzjMoiTbi/WXLXV/g+MCvVNsx4FLjyO2shj22yD
H8MqUMqjmdm7nI/E9XhNfoHFGj3oFzzjFRdpzQZPqWyY5/gt8SK/ueReEUTjUZOGt1s8h0fbCp8D
xI44ci31dGR6S0P4+L3qRkepxaPOdeXIoKCNgrfGZ970x9lxuRK9OFJZWr1LIbIgLcD4Sn6yptuh
ZA7OWQWdcWBWQcSWp2LXDSaD3P/uoAV1cK7Ax9iyWvlnY+S9Dh9QHY1Z8+pZiOCOLP8DEqVIxobj
Da2DkY+ncVYUKmcj2uYUU+cg+LeUMb20jZebNwwLP4mKvMq5TT3e3iKPj9z6uSOxUJqYmWBzN0LL
LvbDluM9a/KvCdrIsM6diKBAJ4B5hx999XbX9BEwa7Eki/jaVy2mZU+gcRsnzHkgohtrvZVMwFJe
7Iu5/XRkq08R9ubcykKa4SLlgxXOtlSuXTuSuR8gJmGn9fc+QskaHLjdDckgrg/sb0usTUV3BhO7
aZPWaci6Bk77I0AvwE00sgxUEAQA1nrOe+wglsgVohTIbVeKwd+uw4jTcw0a0F8WKURa0auhWCet
gq7z68Mj85TMkoCvPq4vd6KoafWMbWhdPqEg3SBzZ1XZlJx7ZNql/OnWZ2rLPynI+pIGmpRdz8e+
36fJtoJ6BOGkLgOnCbz21WPMQDFLOR0VQuLnfjJKHD+8LXfxiA7hxaK7FiLdCYwtBk5auGDoeosd
oweFsbCqVXGiBg4YC65tXz3+R/eAZCAMKhF0+s1+6xCMsSZ2uMsiLlu8BkOcGkR9HgtDEsamzNM0
Sm9/SNUAsokd//uC5NUzJQzinoyFub+/7o1tIyqVu1sVTP5dn9X97tVc0RGh2A+dkgiKaw9X8hhr
Qij3VbWAegrkWFo1QtLFeoyO3bzC98IWb+Cluqh8S62++/KFFMPGZq0nxfijpJz3v6ZrbCK3mbTC
m2EXiQtQvsXalbcZqcj1iXCt1sioFkketSvC84b3DrKPKhuUTKbC363USy6WXMea/U76+IEC8oBt
p56zLsA5r8CefiSpx/fZv3/M7xSYMAhngFsRZQN1mw7h9jBHOyvCRyVaC3xomLp7aBuo5WztwpSB
LoT3V3uYwDUCIgmT65x3yFMkI2s30Ck/e4fupPXlBmpLJLXokSqsQzedU+Xo0gS5SYeqkHhdSit6
kmxI3JPsyBeVispXJDJhtrIZctR9BXvZAMU/GusThUbI//zW39WSV6D+1m+IEUIeOGc5KvMjnZrH
ctKSvQBOwtdsvYo7Tp4AfKFeeCv8StEEwdlZLVxYArH28Bvc8TxH+jgVkhERHOYfGYAr1PutdxMA
4TjnU81LvsaOyVDiwdqLGoWXY5+Ucyr+TnZ88L2E5GfKNWNQgVx0QYrS0SFP/zjrSPC1HhkI3r/Y
1IyuCtQJ2/yLSEcUmuITGMPnUUTMtVeVVoGRIBeRyM1NuxeMa/fTlymWceLPtfF2DVx6p0Up+COi
ZtTUYKp4Oc6GrS5XlGXMwVpU1wkZThvXOlG5dealA+O3JhcGexwyLP48n79b6xbAMmzyy91eNO6M
a1KzhSxltxgflZd3FmMQdxjtzf1ZIJ3CKKNbkbqLKLb41ehpIgmiBJtZ8WmBkSVR7PROKFXzw/qk
aWyTr+88CryC7DG0X98Vp2GemQFVrEhe8IJmxrF9tocKnWjm0ESHYrC3QZIeNQRHor5tbuG0JVFE
LCrU8H4CVU4ofwlEo9uJNGuiwgpG37KeGBR5fK4esnv3STPclEJVDTbha1QkKuV2gkA4h+N6ZFHw
c8lt+bi7CBzoxseGyyRPZgt7nI29y5e8AgDi0al8l+5pMu5oH9glVhZqtlFy0WU5zmK2+gM5R88q
+ngRCe5WyqWRUN4O6c2Zvbrb0isWbmTH7Tg6gEMI3257TqIE1MPHtyt4n9Qo1PsdBSyURaa/zgo0
EgonmT1aRz+OtMdiK7bSI7RGYLiROrEXgJIdteKjXhh2BGcDP79jqYUTRNVWSR1114igBf/5TPZ6
aqiHYywQRERlTUmeTdiGidoCfsvZGUd9qH11kkmQIPbyvthUKAxJ8er3k93XKNRL5WQWpQxBUvGY
JnW2aVeX4WD0dUkNSBQ96bxhlsJuf6+7eoF49Qob0rqbDjQO3RCXasVYod37Fzy+YdLWj88HCWA8
CkPw9Woxe92so7/4Z3NKQEIBjHKvVRdJkbJP+p1KCBdHMDacgpKp7ZlUT6TjGiTCuu6ygxNWyvbN
NgWMqNGNK+6rnyAkXyKi6WsZyK7ZIy6ivcbDih4ESuUx2J7r27VjAQY672Pw2qCsXUJCTyaMBF4u
HaKBZXWlww4cPlkYrbFb4QP/ee6CNV9s7QAsFpfwHUwEuDMTZuh7jlcKdsN+aKoDAeQMmIvc5nYW
8MvZK5GJqLdWNyicSTY9OWXGRXFo77R2YmhO+B5xPOh+CRtf74bWxOA6Bo/b2E2j+5J6sX5d7FYH
tC+XpZCx1/q/C21T1zilOmmTuOYilD3p5nMWzC7LYZrabbn1Sd3x9qz06902Y1GaN98ixiyE1Bhs
coZIZT0RhAE9Jka4KsNHFxtk5KLwPTJ93bn/EmgEdCa+ETc9GCtd2Nx5KipIOOdczXFW6bLwt6IP
aY2LQLUUCLeXljCE7KMJm3WqVICUkO1dI1K0P6iRz3cp1Oj3prss1W8Wd/84Xoz/2VjlnuX8njBa
Fd5twjHPPixgd6QJ2SW5thkDU+ZAKm518492/E+k6S52vE3HLJF0zunS5wTtApL0jecSjXv0pTLP
rAhLB2aYhCMB49k1cbcd3rll315i92qYCjR9Fc9LP6/P6jhIQiNU7D3SwslC7nZ3DXlv6tGYXJMm
buRSroKRPJzMf+cQmwh5SVfGrK6rCHf67nJDrH7VFz9gniz1DS7/osikono0nXwLytgp5OYj0IJk
rPqYhQFmZ5y54cris6iW6hFLJVpU7wQdozeGqJFskQeciJv06u7vW3q9KrrnhQB6n01QkFyUAep0
ajAYB+3D0Tl1P0WhJzRsW1fspI/Yh2LRs0SiEmOS5UQF5UqkVoV9DMMbuqhMYAob+jl7yQv5AaIv
xznPfXCNnqVgD6O4KX2Y/n/kMeLY84QA/C9k93S5R3sNkt75DH4lbhUAx3mBt8XwXZo3Az+flGQu
xGasydBgdC49klUNziSuEBApLQV0BfUaX7X3yUORsM4TrDkk7syZ36REOcFFqsJIvvujSHu7jARM
HNU4rXFKOHE3NPc0/SoDJ33bb9JMhWjXQyUjfGRdMKowDAtsT2CUNBVDpHkYI7lzGglCfjlva4Es
gdJV1KOea+D9mcRcTRy2auCfzdVK7N/eCKltAkyikMPFCEQGralIoW/cq5ai3wU4N80dmmdrw3Wc
8VKY5QOlDsDDh4T4unj4cVD+J+lShcHNRyRi6PvG49Qe3CBACcNau+5fnh1F/jHWa9htQaz2VHWW
9JdYEVfdwTPXGXuEc1gXQAwuMo7nxS0dQJKQGmfuHXd2fi7MMJkDRhMvCF33lT2EKDJkk+X085nh
5Ytaw2OIkAc+s8+W9XLthkOgwN2v+HVrGFoMO5hhM5S5sfxPnDAcbIHovv9KlyCsC5KrKi1k/0jl
pLUlb8iCZM71Cc3C3rmixeTWRw1klCXmIW6sJzw37gfK+9JjT2TRxKPVat0m7x+F78dzWBx/5Y0h
y0ljVmoOdC5FeCkSU829EspfTsSfHOvRDwlucWSgORzKnuaIQ5HEiUrd8stIbDJ0KQblckZ3NqIU
kf1kW+mE0nJG8iChQk7ye+a/fTIsDZ6Aqg0DCVHnvwFFYNcXOHVsBrM6rdz+NVtCHmB/AiW0bbKy
vgYldTxfhSdC9IYtgNW6Do741o7WI6/3quIGFY4wC3lqYUonBn8ZD+tINDumVGjRHqOOJmYuCjqz
qvJM/F9sKcNxIz4CudX0zCtHjXZviOn490wViJC0Tp9ESbmNEYkh/xA8+nKk6J8h8UHpoWdrXhst
7obUffD3uCxribJOof6AZrLiQ/RALM+6kazQNbeKE11rz0KhGZIx5/s3zSOuo8MRZ5wtsER71y4m
TNxLDajnGA9rhOWV6MHfgsfh1XM4ONss2wQa+tAcRuyVvV2chOLzrA/wIqSRj2u8X1PaAwF4DDyn
F7beUAcwsBZS0yKf/T0pTXnDPef1fPCODxys2EhvnDM6jBiEeDrA7l4qaiyxV3YYzsivEW26gfC5
dLjkMGqcMAAN5kbOcv5Pof3il9Bi3xxNEzZZe0TrtNTsdTjqTgZwxU9mNe+Jhd1qtPkCAfVAalFp
8Ze/dRfRmdSqLiFoVfpZpBJLXvWbUTsFrfV712kFGATGdPIgQudET6rSYSV7Cgd16XfNzb3t/fbc
RLbJ95Ib5aTMEdmP0ymX/bKfyIX8TsZ34YhTq8LTG2huYPuRrtQYNUKxnfShSFDJIgDqjSN5PQVw
2lUB23GHfMycFDRNpqplJX3+rtMnJ/syVn/qWUfsWtssXO+66Eils84XBYOK5Pth14+pqoMzSmR2
9WAQXCr9/MfGLSO8IWmzhLjYmVInfTrzMnIFYNsNlfTCrAsqJ9htQqFl8g1Cu5WLBSNVxtkekPTd
OHVh1jHCoWHsJxOkxkxUH1PUWrfw2AkqWl4Eae2a+zovUTt2EbzEdUoivvLvuGW8p1ly+sClGvnh
3V/91TcdEjhMDb1Zamv10L7pAOuehAURnlT4ZfMSmEOzNM9ZomCj8TsFSzZLYWPzL8Ng0FUMro/M
B80ryxI4uZxbbbU3slXZtrq2a25qA2/gzT3voxjeixDFmoQRmvv9YDltJMO+muDVbp5iyv12ZCBa
0UwHXc0Is57AlrRtUhqrs0zKVqtqKBya925XdTwA3xBAj9stsEKeQwPYQfFIb37O0zMyX5Vpl6M/
8YV9mVnQgHt98JdTF8EauxApSIM1IyXQa8Yxf0YBLfZppL4QcSqJ5TYQZdni3go8hoIY64vO4n9P
rxArolHDHw0h05WrDQpwW7i2QKMdmSC8bxpvakdzQu349sC+tuJa7vQLtXkIGcGbuNU1AR/TK47j
ou21v16IAT80uFGNdjsbQlMv4GI/CzkNnvb5mlimXCpF3Y2VzK6+fVPfS1NFTtus1YkLxjj9XrHA
MeMoPk506QUi3+7j4HoKGuGKuSp5BtEJiiIPJKXaOk6BhCdInhUzECAK5jQOE/RfKkEXl2JDPX8P
XEwAh/1yhQDo8H2XiZnYdKYTtcuNyXRWhaRZdAf7mopOkz/N1V7KUr6dZ8X5UiyeniDIrnuWY8kD
lXmeljt0qvHLfFGRtDzTXCJtDTnijY+HD6ol8yLq9pDbBLh4A16f7Uze93CB9YtFIMZ6MDaZA6RU
pohaFCG1kuKnbpdAMdq3wV9kqPZxj5EmRro2eOJBt7iP9r1CX2LW//JCqkwhg2Ghgm45fft0THzH
RhysQ+/lbKlbf79SjLvUZntNqitcBvKOhF84buCnTb/R3kTVnmAZQ88fS0uORR1TPfFPpkF1ibfI
19wVNHyt7Wn22l9OdZ2zjKERxQnP/F6j4S6k6Mo21lhJDCNeADD9xELZodO0xfAhSXDKfv/7Vh5v
88r97rTul+Mv8oLolsgrQThtYhQUkkmDJ42GWK3aiPjGTSXMaxan8CU/OZezNrDscVO/DeT/ms0Y
IVTmw7zNLcEWXgF+8P4GHVxObH+pbdlpzhD4tXIppmntm7Q5YuNsbVld/EBo3eJk6+MjRekqPVcn
ShXuBYMPd9BvfRmKbll7fEluQ9ZOQj19DI8a0ygEQYSxhBt/e0QsIwko/j4irI81AK2+is7rngzn
+UUOQQYMxTK2jNhnZQA7nz88u2FtDksI7KBfJTJsCl3LHOjJAxGcCtKQi1E0Tr/a9g7ljDZNpU4s
3mgyG1+f6fkviUQNMSUoPmKTjMl26Cx9CG1Lrjh1/i9Q6sZ7QRTMAM6vMqrRfRv49aN4RFcce4bz
0exjUd9E6NP1TVn33M/t26M5JN4m0yh6EqYDfRY1rkM4SXj5XS2v2wdfj79QFVzlnKgyuH+aSwxk
TWxNp+DA/c/l8YaxDNfaW//i8QWOPI1qELT5HpS11AgEgk/OmV3KW+l1Ou23U0t7QrOBwZ26JDSf
22cUg/9Ajw7IZ1oP3Cvlski10rs7UjjhKq6/apsOEn23FQpPQEh9RPFfrKqfB69p16JwZNYSTTsn
hT6RTivK+ZiGBXXpBE6RLEKSaXxQfRTagC/P68Luvuu1SPeoUwbTSo7sqIffBMPLEWzzZlmMpqpo
ZQeP3gUKnhypRTFOiovBkCqd3J2L8XQanIm+2gq1sslZ59w6PEwJrw6flKpDoYl02tC0MHKEYfm6
7dAivGdRSzcPVFxMa8FGsk65Fnkm5+xf+29GYaR/jikD0AWCbJ23t1zLvOqO++0kD5d9SERzE2S3
iPjMaOOLhCiqsaC8+oQyqEfioPGIyZdWaw8BOpIbvksxSDMf0Kt4u7dxwKO5YI3YOrcT2unoKZ69
IpQMnGPl45NLo4poY+jDc4tjs1omfBz/1DT+4sRWQWJpDYfsr3Pj9Oo5YUmW7SAS6OhSX1T+dc+r
Ftfntd3xiwpzFdDKppPXXQVH5o0kG7NleHyc1ddqOaVr46RdILeuEqysde6E8qXO+dgQSt6s0JMG
jiVRXFIZwwxj+LyFzRmE081awaL5ld9dfQxHpjtS5j/DwFQ2GS2kzxnkU+abB0by0QtlorGLnTOF
BfxLt9BxXknA6DxL9AwtoIb7PMlOhLwXKxXpKAl13f5fDz6lnS2FYf1GuawkzgBZZ+si8aUJ3UyM
3JevUmAltbNFzf96Zi7eNE5DEzOkXVoArO3Nuve/qpZQq1EZV4JEEzAOabqllrxU+2xRmQ5wb5mb
6nYHkdoAJ4gNfyp5qTMJop082uVM9G6CDqkONOAc8gN+NqWvFPzMsSecB0zCTksFz1IefLBd4BtG
XDrctHTOvFIXFhDWHVL04c0bno+uAkB51usA0dgGPw6FLkT82X8N/S8sMHmYEkPfjoWCghf8QlXE
z5BM2N+f7UCBt4SlBOr6ucG4Ox6+wQKe3Ho7wezyvLQ5o4sWiAKEq21axQ83KCyoRUiHY1Ztpuyq
Jd6S17ei+fMmg/Wn60p7dohErEwJ4qjpVthQAy375ml1CjMVuxv46qeadzdSfQKGCdorT52Ieqgf
0bAqnEc1Mp3nNANXzRCE+0v6rpacSWmqxx94mAEwy6JOUPec03EUm+CqB+uh7jYu45jWD2ZihbTS
kC9t6pGPaeWZHb6eTmzmTrrBhs7lCdEqe6LiYKSgQacYdTqWb95yhOIjRQZ8hxrhaqi9hnNqApgH
uIvbubQ/s3irriEDah5OMgsTo8ifzNfZ+7woZ8bYoOP8hl3ztZAZZaztYm8EVctEvir245uYjdVK
9DKa89k7DbUpp4AMEmXSmZwTK2SQwHqGsluD1C7a+XJV6Ye7jM5CbfJ4iAxv1CO2L/N3loraBY0O
nxxVFJBSFgLIIJ36CUH6bd8VZbvAGHOu5OpL8ATGjEFWKG70SGDBwTQ5EdnJKBc9RngOBXT83Odb
U9hHONLsxeVVPpkMf358VDLYT54uIScno02/dH34V4PQyixqo0hqCUv5n/QqBoJC3BngsGNglNas
+B/ZgK48GNr2dMWKqjibo/DvR+Xj/3GKXCfANd7y87nh3PEfUvWvkM2zIcmMCmHB+8cMlqToWTkH
WpDuZU2+gXEU5NjPlgEWwThCvSPVnv/8dFrX33hdO/JsLZwOT4IDdo8b0ZKsc1m0wVYQ2ov68daP
YYsECAdxXV6E2oesASfoIb98g1ZEh9UbUFcQEjxsXqmM/GIfhwykMhj3Kl5C4pqJ4Eg7vs2OOq0S
03eoERKYDGtFf0IHH7Yiv7rXShs0il/II6LPuX0ngRe544gPEu/MpHT5a/XtnMeT/qAXqPWG1FWx
qVXpf+kM2NkG/y4z5Mk/KTmaCkEX5c3y+EBN74do82LeeaQ5BBg9/2lh4zC6FOlnzO9001kXuCpU
n3qA2uAViLmjfMQj/5BJYPKeBAZ2pYLZLd3yNlUIIyepRCKkc3W/tyPbzmIatR9QLd2MfvlL4L4B
D/tFxvrvOm0NRXcz6qQbA5UGKTbvmt2HAWF+Ou5mRCYCSSyaHBpSsjzTzrdv6Fr/nxJTuN/RupXZ
lpwpPtJ9ImgpgNqjc2U0T/OBJAxu+MuQg9Wv+XOCQnsiS1FJGwwbM0f4bGR/u1bUtdaHBBCQseQV
V1DuibXgZvtOp43QyvLU4XJZ4Lsug4UZTQhb11KC3NqcCmXD2mJIPgx33RHxifD4LwVeIc8/vNM0
MVWZI0iYUSZsU3zgrMjI3vFPl2do8mo3zgR/QeadumU+T7mGR4r0Klmdw719Fk+AEGRZ6OmAmfs3
YcDlstto4IJseVC9h3q6LKy/fzvtpooHEFenJIdV+DUaSTDBP/b5r1BbLo0iHL5ZqBcgEBtfZoCi
8LDs197zCOnDXNKiwQUDvnQGMxgEVxEO+oiOBaX3rrXqnkEF3MjjskmdqxMQQGIOGn6P69sqn8rh
IBJPYJl+EFaVuIEHa7Bx0SbWX6GFiNfAeCPZeTam6Xb4oUPkL6IYilwwoDLzDfF75jDH6UiuxHsK
jj1bJ0ENC/0WvrZ1zUrD7wAX3aTMoJSjBZCgRok6P3CKegAgtGbzEqVlPjLja96Nu/9TNy8ylVbO
OHEOor8AjC52Ne/7wNzQ6XPn1REpfXnYZ0SZVMb0Cls7wVxYeyzOPgtEMA5JYjXNSuyPGX9Ga8ya
DuOQRXM0OSRX/CMjQlk7wUM7Sz15ZdpGH01wU3bCha8p1KGs5yH7DjkOAs/L2uIxhCaTZ300eK4O
nxegh7tVfIE92QmbiVFQsLyQqQI9ZzL1Yq5gshEILcuzUd5nwwdQJJQMLB11FDtSDKVj4tNg5pnS
dJz90GCw/4eAyl36lhtffKyAcKXOsrNldg6b6uwmHdfAYBv15Y9TgtgZdaYIc1vdTL12iibNJqee
NBwzE+1dbffcfxBq6gafCnWze/HVHL2VKEknfs/nOUgx2+rJUxEbm6FK45HM/SyWHoyoYFU23oXw
4RHwKtoPcTwiFnDb3e/PvyVDLC5e/u63Igg4GZApQi60xJDv03/2CaMK3Ut8vZq+qbVk2nltsLLN
73aUMCkSK1+4BFGWXoYegQYByR7Zp1biq4MD81o72/iKW8VngI33L1u6X23TJmsb55IELgbSDAi6
PWTWsfx8i5ygYKnPUhNAXm00hqgDeUE5whBvxM4IDDfQsBRfxtfJ6cfkjTqeRHm5xPXp7KlTI06O
AvF69ExY9W2h/Pj0jgfEGA6h5xFJLGPnlcCuhFDrFDTW+HL+pyWnw8eCbQPv4y/k1FCqDZ1AlGjz
oiVLK7isgOuWQa85v9KT88QLtQT0yNVx9IuVPFkDqXk5yHasgvrHWOTo0j96Gn2sSupvdVzOJcz1
Z7+feg2nQoLYOVxiwh2UFQ71PaqYXRgGRI0sNNJRPzhrAG4quZP0MNytW8AQG/iF8aAcGhuSQmoq
yyccasZDCkWpL08BJhOHlvZstLUFp1pVDSCoQq9Qx0a5bvY20B9374mfE9QHxkA8+FTULwUAoD53
PQrE+ku7VpokN2qupggkSudRJ0V2ezzCmL97get0AfioPm/QZ4o244YRLmnNfiinJijinprBzUTJ
HV/lhAbkoGl+dFfrBxlzJG4QbGtsxLFczrRPibu0MYhLs+uyv3pLz9oeb3eH9gXf/cig1wIP9nZV
An5YMJe/oS7H+3Bz1HiHSZhvZPXrnTZnhT+rM9P+K0kIakbi0P3L5qSw4S5v79KL8+1DoXiS1R4U
vsljDMCXjo8NCrDheTVtRtdOQOLI/tC3mGS5HOjDe8cQqGB777eRWBgTYpbTkZ9l32CRHfvLkW4C
f/m6BAMj42l6BSoYmGebRDbLw/Rq8vcv+03ieT6TXq8ubFLnhnIqbWGr3pHvkk4eDk5Cnn7eyF7Y
5BucPo5Aa2G3G7wl7Hpq4t7NnV7B+UpjdEuaGmELb5te/JVbr0BwQw/yPpQ2bQqtcAC2GUy/syVW
dE6m3vz4KzBQbNXnVM2EQp2TmS57tVi3ASWqSXAGbPqRvVBkpFJ9ORvFrBCKBnvKN4NqIn/9oD8J
yGzlbmzQimfMgipjbL3PWBPFsfvNzpL1qydTx4yOWd4R2TQA1Siznb//P0d5BN0qAATwn6uYMvyQ
UAC3HExCxTUJRmColA2evXi9Ld7OQmkW7Kll7UxaPrgAxrpgxobggrsl+XXForMOCbe1lapGEuoM
Y7hs53JVal4nlBwMgCo8d1mMeQZ/J+5VEdf2/IxBXKPh5xrRhlJA9Q+zRIuqZeP0P5WgqdHZ5tW4
WTT2mugwOEsRDEgTCwccdjmn/19C8Ef/sbkqTebJz03ngp0AKJK1JZzUv7xYelZDl4/wa/lmPExJ
f3zBGGS2Duk0LpWj+93up9xx6VeNlfK8HdTAP5g7CDMr66P8Fz7uUKtf7hTMb1cXrICP1rNvfjH8
kKJMTqEnVf/4tA+cBJX20os0fFYBt4if60Cifqdc0VV/3j6ulHI4pvLxNb1D7XBTTlwpTii8hmLi
Ce2OQoX72MfFrmBgSIv2bu8NRrFXFDMoTM3zprujnRBJdG6+sIX9hB5+YnUnv2+jIsy1Gzu5bKRO
yBKrOeof/vsMZYLnnOl4Ulcl45cuzqPqqj2/KIIRuOfRZ5VHrsGBzsfK+XG+dSEGjJs+yRFNjScx
ZUYgVVWJa3aDQbJJbQ2MV5YLor/snGnr+45IqVyE61uUMnTWOJUXkCSFnSHVgaU33+RIuW1Gu1pV
VQh8J6wMOY4PhpzfKHG+KjZqd4st66eXIMjw+vZrgisA9V0SYDsOcNQbOJFNQerU8dFFD/CUogWR
NwMQDvVzX8PAcguZn6MiDkqx/Yrld0j2QLq3K9N532aCfnnpvxZzqeNX2n+OnFcSCM9LAQ7vq35W
epgfDSkQSoLf0UQWcsLzKNopYgnV5CNYABvIWE0lA5YKuleDuv4iBSPwdVTWDcsa2bnrepBRfl1l
HQww42/wjw1TlEVLbKpjVYp+k0M06dmlL48bd5Akhz+5OdiSBsSlZ1r+eioTwEHowUoVIpFSckKC
4kGhja9QiL8gwh0VnIB/LgJJ3XJBE/d8bViY0IHQZ3qH4eYpB+YOTlxg/C4bpPCF2Jx0sBeYs4Py
b/5bYpYka42kQVPbOEcy0ve1hTVLv0cuJ+ziJ7RP0aKbpMXvv+xuFPjXDQMTi2l7TK5xgAcc3irv
j+MWjBFmtAkUi61MNpib4mDX4hkbqxthKdWELwW16yW4HXC528/bGDwaoVWSB2ZTdSGdEDXwN7R2
uPIN2+2JLtAq0Bc9YQehFhYj41NwiuOc9K9eeFBmD5YP9xkypH1qw3MQT/yLiRoYuOgE+Bd0g4We
JxYKXyVYbB18MjzbgTH9qP0bYR/mUo7no16In6bpZVdbrQLBJRHhdXMIB41iZq2Pg+pWuTXSbPXW
uXwU0Gt6fkjuoifiTOojyKycKZov1EvIIjsi05RXHKotfxsyRC37RBz2yx/mu+1QVxN7Ocfg6JHv
oUwMR9GH7rwChej3YqLqYfF5edHL2Ytw/VD22X6lK6BJo8ZEn/jrUn41dQ2haNcZdJVyonGWgG9h
IIXEocPqjCxzNReaL3FpxQWwNNZHX67wLgwuD0IMvQ5TDEP9aus8TljUq3jnxScQffVh13VlDJVi
eOxU1wzWWGHRMGg593cz1qLwxdKJD+uu+hdmpkRaCQ22BsSB3Chsrw09F33BFtZRICLeWpeWU6d9
DH00FB8nArmfiNJYZahHVCCFwEAMKAZL4V13seRP7UaYh6svCFRtwgHI3buMqMfaPONEottxcKWX
iBUF5t4ilsz8nxjWpmMvvnPKCg68WSa7AYTRCpDe0MW7cm5K1deDypc02Ny6ljAlkEiulotDYMZn
9geKcpy2ZGzVzQNsdaJAQkhHHU6WVzK7xXedKyXLWVJDzxEriqhZJYXCZvqQUuV5qQeSugIP0LsK
Wffaca+wjAnqZKiLM5IliSvcS1t2n1r44UvI/H0whl+YNXsQFCqxrFVyxTglZypPioYbjnwXieM7
tRQ5v99rrh098DTUFm9RhsYKSi2D5X1borEFPGl/KGs73mfLTJhhRXkK58j5sZYXa/3tj9laZS8H
irnORGlCzbAMQ6S78waqniws90VjwJMYjMd3fPOvmHra98EBhw+awdtfdJAwPrsIT99XPqgzhT0I
qtflJFRwQzk1+yBE2+ya+5eneZzp+o0pD2gHEi95sXxlBnkJfqWsUIHM93wimINEftjcjhuvyxRS
QIndUQdfg2owBFAT3bvPGmTd5kbx0p6ONofgXvkXa2fTPDgyz/bnFsRoiHoRK9ZutstyMdJfr0Zp
1Ql6UN0ZnZZ8sUXIXh1jPjBi6rzepOq1o+ubTmY26EQcOoIwD2yrhRJL2yA4mMFXI1UZ3L6eC73t
Wra9LCiC2p0HZFBXsvmHg1dEczHjvW59omXKZFCIkHt/8UsaWzVYs8vt9LiPLqtItbeevud1qJl6
EHOrAH5IKrJYPCjDHd2maEDY3WdyLnGl1Oj2DY0zoIsYn6UGrrmRXXI1U521eGIMlAYgSf39Wvd1
uGTtSY2osSbsX2fRu2wbyx8YKDLHJLjUHDRramC2lnDWSOc9EMSD7cJcmEGtigyWtdWcYjnby1Wq
AUXAsEyeaRi1kWQVuRaL36avdUO0EKwXoX/P8GVuIfGtyFmfwkbnG4K3gMZtyjaXNw87SMkuwdt4
xgTL2HFEk/ud2hOXxXbpVSV0XtRMY8AJMFPpo8rbzV9AQTAjzcwyqldliUeOGn43RDbCAf1g/Xn5
NKxrvoAn1AARFClGgCOEAvt3nyZG9U9L1Alq6siTytcDU/Q6tuc/yzMoHEdUmD+km5Z4LYht3+QD
LR8kn/MV07+UrN0WMJGIucCpJaY8sA9+bWv8xdel5b7TvrRojqlFiWWjdho9lROXm/lvbKz471og
hoJ+Sesy01Lme7WqPmKNsRmrWNkTiXuA72DEv/5ULYC0ONrpw2VLgvmZDXnTOZtfmtkVyfMVt17m
/sq8bU7U3gPiPwMeqslHUrUYtidZfNSYe7+palMnNV9LkELESMupj/jag8s9Itrd+dl5b1oNB1cN
9+aLT2wtVtNisJslsvzZWmijUT5sGd2giS96FUVvrHMM3gI7tkHFQ/6I+hU3uvZUELoVEOHqbN7V
sFKgbnt/DwzBs9VHOHmccMR9pR6Ktbw3rUBowdgR6/esft5OD3xDHE7Ue1SLT632dtW9jtmCFhiu
UObQdvVf2uhRfO41wD9tNw5leLBB2moLnMgFdeQHY8kR/Sz0h1WQS0aEDHf2D4ayUg0G8xt7Mb5C
BDzYxPpsWDSagLELoJxqk3ouxkxt2WaJ1M60NcIWXk6sviDZ/Ch4quzvJajrsUtxN21XJoV8sc1K
eJJqYElyquvJxNjomP20wbFL671toFCTNgViv4pbgROX/+V8kvklp9qMmEQP57adOsXlVo1Rjd2q
e7DSNF5HFd4ek3cxAhvpS9IGIx0KvroV8lbhN3dbBHGgt6C8HXa5qfnuxBvzlRuLJ5H6qrQ/FmVS
h/gZgXq1qg5jYz/gXCpsi+F+XQ46SpQ+UpRD/N7BU9KGy/AzAGJWj2Kv7gTuMqdiXaLHsZoKJlHU
krOcfR5m0UtorGjj5KV1w2P1rFym6E88O8mvrh5hpgbsWJwSky6qU8b92I38rZDiRxeNQs2zkoHX
zSW/CmeGu0gWCxyyEKxjEM8vt3u/xirHX8sALMC/10Yjzi+5ZJFi1fToL8u8GQ9N0gh8uxcWisce
gqNOqiexmUlAKdxRO5d2eDtA5oaHr0e1pRovDTApKqi94K+Drh9TPdhR4EV5qoXSDJTNd8suFflx
fY9V/S4OuVAjZABRmvDOhSM//GZ8oE1ZPZaSLVPqqhbEV43dqXty7nyR8kXKpLLxOs7wHsd12PZS
zXJ/Kji5nMtcqvsT/CBWu37hXSRClb8X303j5yJxKQ+oodl6eC/AYm8YOqCv9ToGhl9cB5zlvpfS
JscP1nGI8FghdA9gatYTxdpgGhH89UzXG8+i7ZcATFBOrPIV8vrmRzTFZrn7ESs4Md55FHrF1zq5
EdKrTUTg3RLyRysXPuziSH2gfxzwTMbCWySZeCIZDxWR2mtvb6wZ6y35xW2kgUyeFRntk0+l+Xk+
c1UVnfCT+ebEMJXQsjgWwcXAnH3F6Pdd6++Bn0ZBVUY0ELpy4McJYyejt1JhIxj3SPuK6TukrrEh
67BKoxSrwRhodgWIoFYmPnB8fPOWR7enWn38G9ptq7YofuXvtPkFZaq+aJ88XwSzSNhBXeFc4CsK
KJvcPYPD/tU0mzD8tg1ULRJ78e1lMEGBde7Fbm085Tc+ZdAjENdHn8w6NBsQO0jmD/hD6YxTzGOm
/6shOQ/Qp6DV2gPVfHrryt+ggKXHJErFaF0FxM9VXi4Fgrd5RwOOAilcAdts9vpxz01YWodVt0ET
fHR0/Ev4UotIC9ISFPx0OgTtmO6jnZPyIhArv5Q4aeU7X7nmO+VmCyEXoDcrmzNP6TZyFNoeOnvB
brMHX+dLppfs5w3wS5w2sQ+ur+YmAh1gUdhq278j6nbIAgIBnkvX4tRLGY6eAeFUUo4+YJ5kBMRX
4rqif5iroAlk6EqvKMtCpuguTfwiIdV0svl81WW1zz+YVEt2vmy6EcKONzjgsTXTQdtQRNab4fGm
H6U7u8fNPeeuo2Jh0KPxVwaK7rAri8UMLjDBCMiFrXHcnPaVpY9Vz/cbhiQij1Ev2EXSHMt6sO4k
srXkInDKHTIyRJMtHbcZfZuVy3j+t47LemsUysM6hU3r7VPneKHCq1H8TQYEYp1Z+70Q2eVPfD3o
K2u8YNDGjWrOOOveGNOKS5q91XApxeZvR9ojlcphG4ayxoknilR8NVXxP5oyo2nP630HiLNs/ve+
1meMyBJiRuDoavDWErqr7SSZ/rW72Bz7hmEYnEImFAmu2g2efk/w6x6OAMIc/uJQ5s3RBI4FeZlf
j9Z/+/gZGuBPQHdkrntXcEsvWCG2M9sD3mJAGvx/fxNRevFRi2PYxJKuTbrcS2Cchen6Mf26fou/
0vXpfRhZLOVHyguwHB7wTN7LYscb9pOCVKxNGLuPpln80ZCl8q9pVP8YGrXbz0dYYlyhPTDxdxWw
DqvyTo0PyU4x4pJr+ErYDe63Xj3WXxql22SxLeGxiGRuepAOo5SVClvGe9ubo2+Vl+O1fsNPzt2P
P5DMRchLPtyyzReRvuIqD8SC9xGDjGAE//x07dNxlsK0IoHxFwbjTVzkV9Ocs2gR2Csdr65VfNuI
oTd/MsATSGDPk6R4OJrKg+/Pxn8jHlUvQQ2FTHsvbkx331tBS/KSItmkSXCTFJUMDK6IQMEM4/yb
9sQ9O13B/EfA1HJuI3LQ40rw/4zdtiHO1T23yOkGj6v6kC7tRzF9mivM6sFv6y86dmPPLw8Y2lGt
q1GfVNoQsJr3q41tnXAWvTUDR3BxAc6JT5yU7m3rzKt2uPQrbbCy3pgEuIj4XuE7nEXowwDAEMI2
rXaLno/vlGeEtkwEq8/40qyjicTEXvvcY0QaY5ATcSHthB539aPimrp5WIrKzuqfr8uycn1e1w65
BC3z6+BnL9hZOD5dZ2z/N1qMmh4xjTrkgIXOIFD3L28TVevqhHynCLuGw7dKnUL2VgEMfcoa9VxS
eNPCZ/6AiwKs8QIG734Fv1wCFQQ87HJYO+CXuBm4fN4dUg2SKINV8Jq23GfqaEFP8dJA8AS5S39B
otxBaQECDW6VizEFJ0MzIisvNCN0zoipnwXs8KalZWehOkG0eH0YTxJgRJs8n5R+OgDAsBB1FyvD
VzKhTrkk2yaRGC5oOuuKxxzsbjgMsD5fIt+sIPSLm1d9mld68vWppyslKVn/tZEPgWUXr7/VVzV7
/D4OGdRtFlkRMY6AsgaDbD0KTurBQpaSEdiz/bRsRfuMeoJBkFHqAIKRNCF3K9i4yCPAaIfaw9ID
rrC5hN3LAsIBrts1HIQ4tOj6nXVEi2edr9AuW8hTeclf85bFBYj8i1i7GOsbKm+BoK25e4WmtB9Y
ORXS6Tbi2Rn+EKMHsWabe3fchxUf8cwEF6G0LLtKJKeQ/1tGTmgSJwA1+GxQJ3ikd2aNK40I2HSq
Xq+jPsiuxMIFT/OPLw4IT+uvMkyPuf7TOL+rO51zbMV4fdR/wxDOK1gGolEHi1idUJcAKXsPbhIA
4OCAuOm+Lhz6ypIxcekncOmdu1jcJPkghxih4MFnHiQ/yK3MgidNvMW1rrWtSIrWbGw46rysu9tA
4wkByC6pyql7QbiKXpoj8vkl9Te+hXKa72ioxcG9tdGmN90a5BURxmr3L0yv8rzHk7rXrofnyf+e
PtmRyA6+s1fMC58pkjH0cTXT9Tp1AKIni2DsN/A7zwgGp0Wnm8ue027DXbnHNhR+cCav8rl9trDN
Qk9oMpxY+AZkLlnOvjgZYfnsbFslzi/uEP3NngXY1BMzCDfBbBtcDdYduO+Ju63b3+IX6fPDQIcN
hV6zVHVJ/3Y2imnqulzo6T27XY4tfJAFjL0KIkkM4y2FJuVACZXFJfLnOBTRmP1x8RYPNdUwANHL
B2alAFGY2JogTtT5FvL/wXoZ3hmuWEZkezraPx/gpwmrKPmHnXSjsGu/80qaldlTSOFWpfslZSoK
mFLtx9G1ZnY10PVfBfhD+dANfHZ+8WYqYZsZgT15xtWRtKcLUXyTVwutUd29WID9/fsmEuk6ycEJ
3S5rhSNgUBRHa5cy6k/N1f9MVQqAnLCY97gGg97xt9PG7E58/+Kx0fpq8lN6oEHdGIgEy8avaRk2
x/c0VsUqFDXQrd4p3+j+ID3yY/zJCgK5D15/0zAn9feLIxO58coZ69RU824buPadsJUf53QlBEgD
sSDVlroGgx2XCAq5jEEMvC00pd8oE8carU7Rdo3mE77LRZTJRzEomr9Xp1sH8I2vIpjucNvQF6OX
kjFeW0iTfPGP8VriiYl10Rstz7m9vSb6bpcjqeA634Fdd8QGyHiotwNSnNYGFMaGQ6H8BQfvpp2B
agUIYOXCNIqqHlZi9zrLjwXs/mnXRQUAU1B8KLyTCjiw0ymMYbK/VR0ULXdw9LPblEKk+LYr1BKP
YT2hnLn55jO/hdpoxETlKD0+M/A/vqivFTHMDjZQ59i9/0XVwv5JuAHhGSa096OlP9zMLMIa9ibC
wbbJGyupYvfp/65Kmt611TXnKAyhJCvPrca1VrlZpybM0HBSjfABKGvUziRt1RGWAtoidyDKjfWb
GDss6izp59RKnyfKGOMceMrzNQrnWZBHXR9/Z8SCHctdnkT7r4YSfIsGtqHGBc4UJFLsDdg8TEVN
kSaUuaWw2jKE6lq6vaMFax60C7XsXgtTsrn4Ynml1DN2WfomijTTy/PxIOvIcnwNHAwSx5rSBmKm
ga6dYOl3rFwoHOHCEmgbGVyMoZcN79hL8jxXiIhJEZsoftIUZ6NXAc28O1S7g1d0iHY1Dw1PBLAH
3pIWMba9DsJzl8b/dY0VevG5ckYhVmK94hBO12N+fogBk1ucfTkj3T4heYKepDClMuhpx98Li2wJ
KCXWt431atxuR0Mdq+EOJimSxkjDelZQs6XtrQQOllFoVS5Aosb5/RIN2M3/VD+yUagsopZt4vFS
bOC1BtXai6cRVcH8eT5p0/O3zaAZLZQspj/yyZWdG7L/T84XWME3+YOrzu1eCwIresrqwDmdPIzO
eTlWOm2EVEScDVwdl7CAbmBqAn2T1KBUVH0YJBNit4Dt2PGnnkL6Q1WFWxGcO+FQm4+PBHXesnA0
/YjPiqdGq/NTiMr35EL8XMUByI+bx0BHP+rgeKUW+vyqR0/1cq+Eg3AzeP2ThF+K3deKSvL6zLqB
xwDHdBIcnG3ksQx+fMZyruym2MtOXWnqkjgrTddKXN+UaYZxhfzQZQK/F+M+kvxnznmbBnnKtxQ2
wkq9clV5jf+mroaEqHisQcXPlM5mp4ub3cO73mpjjGRbZUP67cWldlGwFkw4IHxbPrLoepZ5l8Z1
4SNaPhq07AyZwVWDhh0d52W7Ivbi0jcU4zZ2c5gVpZ0tezaTyvBbNxdSKvGw2/7xw2oR4Yz6SB6e
4jr+flsQMNaLNJUROrQIA3lkab4E57fm8CEo6r+FqcZ19H1Mgu3Ex+cmyN7L7mDjq3wTCtVbdWks
lr4iRre59x+/qB8lnK7f76TGgKTSgCxC2PbjRIAeB8/u40nrc5WilZxvlbfvIcfGz8XDzKjkjUij
3qYZUfigZwdXNG8vXBtZ/0Uz4bTVxUKjfkGzoPtfGQ2Xjqq9D5Citco6ZJ1S3kPk7vvXy/cOHsHY
PCPii5mskpff+5KsUZpFrl/rkCSKfZw0dDDDfJ+AuRkEeIMhS0VjoP0qCNcFlXZKr2/oKkThl+DR
sRO/fT+fDvsWk5yAyxq8iZz5TMGDAAKL4WTspkKOPD5Y8oiugXTzhDvICrjcsHIlmvLoHgwtfsXH
SnbssKv+IGYfO9hFbrghTBeP+XwvyQTgqIJ1UgM3TamdxQBCt+XqqMEhaYcLFxc3DcLvs4e0XIql
zH0qEg7qZrTSkaHc/JJc0v5cCeRj2Bd/wF230/9NNLHXWXio8ehLioDy0O4zmxZMRsFNmkg+mU7A
+UMSD3+6ay/MeEsFgcUFEIlkfsFe6vSNPh1aoYglOy2YZOvAwO2GJ9TG9y4QOrJLBGDXNMY/sCUD
3mwvOjVuYgdm/xIsgGW8cQ+cPfDYk13BwJjKwqCbmiwXCqRvrlWPg7p3iOLPSyel2pF9SJNki5vq
51eltDZzgLMyL8EtUkf8L9/t130f1FK3124yIjyLgbQPyDJ12lAoC5M0YCrTd97oLe7wBLJv2m7a
KZ8fQLXZKOBYn/C7k0LWc3QjXnI24QC8j89FBq0BYwXB/NQakTqV638zUUrvZacYnrLr4GAiCncX
frzx6AB67EgsYXHytUfWj2BkJ2moPutzi2SeDA0/PAXsWVlPLk9xMvD38IdUzVdoKIqeohyOT3jr
BFwa5K84ko4qwTNZ3AHSnKRo9fIJ6F5VNRMu5Nke6EE+N5KKKd6EApAF8LEfCEc/0qGDgEclCVft
VHsdi/AoEfO5zjB1qhdmmYWlPQypX0fSMTS5jTVzgDi6Z3Q1Isn7DJrnYgNwoWfFSKlfnFOHlB3h
yUgACp7Mv2aHoiHdbLo8FsUKme5J5UVNhCF8ns08tIeFJjcd5jgYlKuKHw12VvGWQRUPHQYqenlH
LBCzaIb2xDhKblDTtaWBgg3z/A8foKnH6RtBAz80sH7FuRmcB8Uf5OwuUyCYMsa/d+8Sd6vjUGKB
BkHlME6xGgoN+UgcjyAm6xd6rEI7iZJnTCn65T8yeP52WZn0hpTBFx7ODWnyinfxkFPeF60gvo3f
l+QQRpicDYtJOyjlcxKFwX7K+D+48Z7euLxUgLf5eGgTda+swa/e5MLhUfGuynGzEZldMMoAy2k5
wtnpv3WBnGRaDrJO07xF+agJAATvN8nwYMBlxmMDK/qsqaZmvRMUp8QHnVAgpM5TIOyRtss7Z0ye
X4AFmmIHizK6am7Cl+yY+DR4DEH7tZuYu/PKjWOe4lgOS2SJXRtTiBtFpnz2U/dDSqfn0+Ae/giq
leCaupjKxVSgOU0724/dCYTKDm27A2PUVSp4V4oEpcDzvH0xk6VXOeLFIcSvgXuU57ghd53wSUri
hakzisqsrtpDQUv88osbSACHS/OsFGLYfsNcby1sPxeo7kegzv9cVxoDg7JeFlbNlTgek5coQWL0
0QM6VItAba+8qAU9TqjXca9iA7wtndkVuLV8tVMH1wMaNDof0T+lltqDvROQ10HOr6DnMFyU4bnC
R3nXGYyo0QpVXzj5ueMuboKLXdYeuz92OXZDq6Nyx2XaQpFBy3SL9zF9KkgShnc4a2xHeQUB40mx
jg+LUIZeac3mDLZqKYOSkS0NW6PZy+o0CPedsT1BmxI/BReLMDnt5sR6KuNDKb+Fm3PTVhgqknEZ
vD1uqNu/+GcLRaCa3x/apt/tyebBFGUE4v/SesR8EPpccDdSE6anIeC2UWhCn24nHqkhpFZEkdmx
MjAjGThtzkHGZZueqjOp9seCA9/hj1UI1W4u8jB8PQLH+CSvceNDiPDDuwSZOWESN0JCCth4ivLq
wK0Lin8A1NYV1NNe6iuuWQqmFJqIkQGlbvwrIcSOY/Vc0DswnXoeKc9caUpLboqLu4X9HPmGQt/Z
/YgyUoGwNoflE3+xe1rexPA19JKWewjf+pjguurECT6i1+WJzoGKo++4BrMoCeI7RGb6Z0IggM95
FjmH8vVER8sabCHlGz1VmZI97SofLJ+Hzux5eaveL76D1izgrvAyBhuUU5mVUXDgCrI/QNYTL425
tRnOu7+eaCYV8kMvjFIsBFOwOPuZOFYcR3LXjomGi6G7ZprtjjOrkOs9atqWMm5No+DwCTZNt+b7
JxGKTPVyMFHwCCZXOcoOh8mTf4vriSqAdoui5o8wjqKpy5fV/yjl/djBrJcI26B4ChxicF+XBHBe
Q8OqiIrQAd9uCRp0NYicKxlvRbf6CojS41zFscbuHDB+cuDi5BQhPBH4OXgAtLXBbxGzPM483jWL
+aza5PouXNRYHETwrTVS9vNXnSR7XLtW7ssYSFx6jhcidhS9o/bW4X554FlZt0gxSdophwIeQfVl
48NJoBSzVPVnIc9I3Ye4OAJrXslTuCLDMToHTTgmo883AUeDjgx250xPuFl0EKw5eiN7AVe3FtQN
376659TkBeDBHEPJqcI+wVKgznyHGgU4OEd2bS4WXTH549Holc2mdvBdt6j7drIL6Okq19HtLxbQ
2iF9xzJ1YcSVrtKJy7nXtHtVmBzz3fpPu+wsfkKviORxvOAvRqsIHhl9acyYPybDrGxdefYAF/as
lmAjZHnLNwJ1dUvpYPPxlsNvgUUj2SJYwYx8vvgKrk3OxsvxmKTawAp6JFxJUE/y2oyIm9XIvVn+
dw8KeYmVnBQiLr3tiail0zRegwx0HOdmydvyZDsoFGYg/LZOKCyJhaCvYwLFhsiNebYoV5brvSH1
HUyjkZX+9xNnp1CpTi39HFrpVrM+uAp4G23i/dRx5FN8wbeY66yatsoQcza8d0bLzWp9QyaaWc7f
nCh8RiT+hPIYptiK4ok6ejCYFyod8C5xZ3LKWzA8+QMis8Mm3TasMViBK5s2n7GPJKBYtobu+tEX
2+5l80pwIcuD7wmZqHlkMz3LIHTha9uFZ51nF8owIKuec0XIm6tK/LqEMsM1Z8cLjLmnPwdn21kL
zfqK3GjZxUlwPrpOg/UTq57s8D3VroWbdc/hD2ogrB/Jp/NZzZ6rSj4BYdwz6NdwHpEg9LRYDFO6
UN+KRZV7iMiDYfRDyn8AwPxpS3Ct9Vyepa1/ws3XKaUZYojTIsB1NOLtOFORntEtUqvYljA9opUG
Vxob3bMUvn8unPVwK65soZf8goSDcqc6gEBv65EF+GaTNqprtTvUNbtm6Q0FW4s+oftkKD8EyJKJ
5Xn4XXEpBWf9fWtGtDU5yv/EN14hUAvlc1uXnC09Vnyb7aOjd50ficaeSzr6Mub6L65qbLo6MRX9
0jElsgV9qlknIL/2rom9AoOvaPj/9P2t4a0j9vs0wbPpbUxQND1JsVO3q/whLH/tVFHSjXfXhlMq
c57ktvlgI6Bo1g9SvK3kYr9mKilhHTMRt+bANUqHuFbhRjCtsIMeUdsa01QPNjrGokPQRf0nc7mZ
fp/6oCQkZYVCNf4aEN/Wc+zMumfiGkL4LdTiT+65kOp/SZzz2Bu8Zz4XIgG+5Nu/k48QgRDP5gFv
UVjUR9GjfDZKTyqpnUlIqkNQL0IE1Uy0dqVXUT8S5I4es3FKYfcjprejeRzQVoue+2u12GpweJwm
z238QOAe9Dduy+kbBnka6WjtIKctRsCZ8xe324UYTT5Edvk9YJZRNRTqmOIdjICgV12UgxCuMApU
YhO/GnigSbm+EEQPofU1isvbmyZBiu0kWYLBNng+h64STg9ifs29AqzBFDxhSOOHCIYHykcJcfCy
mlSZ12p7ivnwrQv5ydmE9QqldSUDX6kVeN05v9w+4PPqDcmC3iYp4ik5w5Vrf5Z6Be6uHBHl7IYb
rnzp+dVbjD56v+ygNKZf+hgxqoEjNv1bkLkcIq4Z2SWHXhnM08CvOw5IgXSle/qjvzOV0DwqFZxB
gc+4S8cDn1lpIMsx0hCSTyaFPLAI78NaXrMoFaVAluE5H4+miArMjSGktICp0ZvcPLQRdFTw0+v2
D7InGme4fPHPDIPRA7xKmtw4rn9KGrjM48oGqBWUUzx8wBNU4kuzXaIFolfe31zr0Q2uVno9izKj
Hm178pmNgOFxIaFYHjsT8N1mbwS4UVUzKKAKWcQseF9awZYkma2JVfuE1Ulai60zPZb0sBjwUbGD
YNGR9vTCBDuizmqtpphVCiqrFAtZRPtsXmJxgDN2JXuYXB8uor8G8QsuOnTtv7eKhMIUmG+1BpFT
5O72KnPZ+7y5dsDEh9R/e5r3FRjj9F/b/9Bd2LoQCU0E1phWGLKcS5sDrx2m0787idz+eT1Qywj8
F2jVTyjYtp9AViLfi8zte40p0YYSpMuEHCeHYhE+z4gXGm9GdsGWesnnbnlg0F2VUQBNrMItxzpT
skaDV1iC/Y/JhQ2jTUQqwxRgDT590Lr65wBJ7rJ449wULYBUv9vIZJUbnPAwvMPYYQmXC5mJwd/L
/KSxRzcsCbDIkQibj7ej4KW7pq1CWsSreF1IiH6TQ7mAgFwApAqbu4e1I/UkGbopFN0kIpmotmEp
cXhVn/S00ONFW8uRLMUbAxm0jF8Migcg6PGc/bw/79axlCxjYR6H6QAI7/lYLpAsIsQ5WF+ccPRC
B99n/9fZ5dpTsfR6YkiuK+549axuilDy1h4zVVfaPbkOBC3RPoVXVmaY3fIaZgJSJaCaPzsjJROv
HcVlBunizJSbR7KZnVlNS1fnTqMKLf++wpqQ9i3xAwrBjjZftG13L5S6ayXqrCoJE4FqABB7MYnD
YXLuvg0oHAnpv94ciQmYiMRFEYnsn8aWuCvcC7uXentxdbsagT5JTo4CPZwJr7Jeka9Xnu0wz6Tv
1m1VNg7UfB2VSYxra5+nmjx2NROvHLUoweKwKYD9vrcbLaSAjzUzZJbhYflLwGivyiFnMZnpwADs
ZpNzBT/aTxoWD2z07znZuN/AWfBv965SNWxfKu3qYMU9/ZCpJFLwKCnWi3IjA9C7wfpQsBcNFX1L
j/OpDSTtl7+nhR25jW1ARzxFob5yV8xpFncS5gWFJL3s6CbEJ10AmD+SLL9DtcCjZJq+ETVmXabw
W56XchSf0q34tnBxZ8rQGAmYe8cpwM2g3+rBAlbGtXAe12iDEwhfAcBcvBjI1J6v9SRr4f+NnS6Q
wJG3cyh/6mzK/Bv4b4tQEjioTGQxAWxsdD+BoVczIUHUfJTkinFaPYzOxCNAJTp0JYcXZH8SwYoC
g9YPCDV93wLZGz52QLAEQvWspVDz/qn9jv4btfn6ZazV/Hz+fySQfAEK1hIqqRqEYyEUNX+70/U3
d8ULMkZshxa186u8siXMRJOITDGnyN3hOyKrxFHZvj1YAoeLI8gKPwMfEIBpBZ5ycSWYCC6Jj7Ov
LuODvSuC2thMkDTOGXA3nzeUB1IHZjSnISGBX2AsSo9BpOZWVbzgIOWwLeD8oY7D7AgPV8FZvZGT
wJKl2+2PUOYrhd7WLsudndqW1ORLMXWonA/RQcTEFvHlxEIU8aQMS3VhMWxHAkyLIknptuC86ojl
T566zUofJxDn+byiquvevZ+gHZZxwz3YTNATxNFCAemwR9mYs+mYJ07a6tna9aDVuYjOFbByPVCy
0C4KFsPEPYSEqI+v/FpFoEuoloQDwLxrHd6JGi4tdQtPWYQMxt6SegV20xjl9OOYwEbx3AmqodvM
APZtoLjFgOEX2pfamwPXwqkGLErs7jL5H9qReGcN+BncLMBmOhPuzqwT8nb4QMyxYzl2+H5yyfHp
XCnyMrXcVlEyDn60jN+P8GllxTZ3t40YwabB7abTKQIpXAF96ldjkpiz2r+yotAhIjgV7V1xFN20
nbkoW20zEdSY34S33N8XSfge4bPTuFWgHIMoDBdE/besi/UeLDNLQe0xjoKEcqmTte/9XYQ/br2a
FrGUnrudsuREnTPLGpcZeQnAx5+RpjRrgTaQh/TjeE2dwzUJZSmM31JNDpm7u1sdTEm3vfxxJxbT
ofiPJo/tS8YCruztcFa4ZtnoVloqPns3slgS/gRDLHAp8Ni8zB1/RgdTwf/zbhzZ7iuxmw2bF2C2
OyiMyIKYzJiBzTAjCVuHnKVdNreDOFTqzzJCURCx7jl+fzVGR5DE9YVDDxfDRzHbDZwbWT0obuwj
FP7VRLOsg4I7jU3ALjm2EHO3zoubUrbShm6QXioqk46Bij1kxb9n96gyMQQxAg65y2nfRAIVEYIC
K2JA6dtcxfDjM8nT8J1bUzfIQLvyvtKunhi8jyPhlrHxd+GPXoLigrtu8Se4jYI2MpRBaBVnXtm0
s3RpM6pvOpAtaVoQ+1LoehKJxBSaZT3cJxElAKv+BwKo8/ddhskTY05XmQHe1YlZHwe9JLxOyLyF
oN8Q/yoJappI04F3K/ltSH3CKn/FQhtCTv3L3jCny6SJaGfUh6VFH+s6FGVM+zo8vEtlAMdgSQC9
ZSl13Op0s7W3xqTBiIdAmXG9Oo6+sTXu/7X36FwsUeH3i2lTpWKM8n75g9D1ctPxe0+qNGHGejRY
J3XRpzwWkz60cD/QkugfPGqe8MPpsbnOzUzRpj1LrZE/AntJvYWrFqn1BmmIPN8qcR9kTKOnMdx0
E9YzwjTrnPIRiLjKiNjRn9eGbDVXun2FbKS3oNVQuSudeo/T7IheNZ3ZYmdJdK7VCjUVjgMabfKg
jVRzDQNG0JWAWWwDOYZ5U19j2OvJgIf9KgT5/R99oGixBONxqHIKveHkaqyYheUoEHoneGdqaRlU
ayqpy5LrBzLct67bmX+wtw8DxqrNcyhV3mUsdjGc3O1zGEo6KxfLFVMJVEnJKb2sU5Asf0hjv8gP
O/3J/dYutzbxYC/kRwSEI+/Vc/jTd9WtDJM7C9G72buQkbNp4xVFTBrJorSJF1cUzugcxEedXuNf
6hhJHTl2zDhYMp829P8U6ZVvQzuWoM7f0UTc5LrxyQvr+/aKuOzBClw9XXu6H1y4eXjqLE0gwuvj
wUXtvBVUUoCsQ5hiv5KxEbe451fDn6EQiAuaw2OqLPet72F+4AvosB/AHOh0yJH9LgisTwZALu3u
pYN3UeHXdTwsVSZA17dYSfZJ+wxqldb8kbwZQGfmRFYYJ2h4b294brXn/9hTzuDz3oozaUbgjpNF
vl1KdpzkuDYfUvrywm32ZqsnbRhqAc6PL6Tt4lbC8qhFG5dC9xQYBRSysshnKfb8xgUje3FGnXsV
t4+M+X1REL6Z2JsLNlhB+UYNGN81hHFyjh03ol1L1IbgHujEjepfgIpAyo8V8qeoYb6JyIR7D9Za
xPbD+eosxQdqSvXluD0imlZcNvIUrcRHEZP7IMXLkNfXoiLu4AjZPK9cDNbVhOFuoNHAI+NmDQd3
2Jqich/VstxEsC6pV3++NjlZ4RG/oT/F3GzT+/WDm38AB69D4l16KkWciesOCV/553SfjNAjov7R
XThvlCmFv0w5SRh+Yc6SlwLg6IpGSSFllKi3G6BRoq8QyaSQcJu6ggMSLP7+b0R2s5jLETCW3LyF
E7blqME5lp0UIDGdG1CVfKn3fO1oyIXQnkqR7egUulVBXXc4s2ti9z183MRcT1jj8LS5FNN8kXi7
Zr/72cMSM6MtSBZz5bwptnIKymeBMl33nkEexXqW85PYyVdm/oKD5TqVmZ43yr8IuZ6lO42AxWsT
3vaVl1k6hVpl5q1DjgpjZbc21g5BqBU0x8uQzWYLGLD5Ht5K/S5InGVf4uukHziKO3x4IelGAfFL
teb4mHGSCRmX1DYdnG1zs7d+GKufCqAsbBSRisW/+ORDH6eJasa6H0D42RFTVpMqx3ytZ6jWvGap
BhomTL9M3hvDnYKOXL3XMhJ06A6ru86ake6+zZYwxTBKr9NDO2F/QxBbaF2kcuzgqnGvrSFY4SzH
iIXrg2bSc0bajMeW1DprYg14UL7NoZ8mXui9zxcjq97BGtnPp5e3/8YzSOTMhlLzz3PwarvWfxNy
c3uSRwo8ht2oyygkjk+VwMRp18kmcHo7GEeIcciTQ2ETe+opq6raMUUGLbqG4b8cNlpgtISRlFrk
y2MZxnwDN3sJ7P4lCd02QLpK/Zek6cuAvhAuU2mtYK1A3J0PO9ICzBeQDjbqMb44NNn+bTGGo2K/
piNgmTuhjRGIjSV1arffQFBKbCIUFwypmIPyrUizqbPYnYBH2b7JmOSxA8xIqZ6dr2hW48QZZ0yu
2Q24DFx2DGMVQrye9vLQCvKscsxPrUi9xNCjpQ14cF89QEzDe1+RJ751vQUlnUwMsoKlye9lpiMt
M2Eyp6NLs+27Aa48mSMDgd2XPkA1hiHwMTUqmFnQ3ugWV6BLBiYLlg0AGK3CoImXT2e6Xpw/veFT
q8J6oGCi0wW9W2Y2QGUX6BD2hwxfYyiZOIk+E3ySKzk8uqHXwwhTQrfdKflRh4bACTV9zMpRozxq
VPY7baFLr7G1edFOZfTTyzxw5A6D+CJQnTeG6MYgNSopOn/rWu9Wnzl8p4cmKOueK1bG9YsgCy+u
lmXhSBBW48/vw1FHP1Pjm9RVvnQ/0LOvtJtT2LJsrtIn85r57Lq2a8p4Rk7goWnT3gdY68iPqN6b
RR0dyQaWKteYGMrgmpSyKwUbVO9i5Xtr1SalYKsn884PE/y+Ok3EDR8FeeOZgivjjgGVpQWc2UO4
msLsSeWEB4T9TxO/82huO4ToOhgdTbI+KqKQo1+6IHnoeUipJqjepO8V/Q4xOfhyo/yJ2ohunA2t
TkzuRRuTirxJMYuCqlS5rEv19IYe/gxE903zm7euG1MEVRInlJkDfxeq+cuABC0pm4XvAIzSHzNb
2IWXmhUTeNtjtrIc0Ysta7IfJbvo+Za7N56A25Jbz2xFTXMFHU2ztoA7IplXNIvIdgSunNgaik98
uHEOmEE/FKt9TtlDKMyyb+kZWY4ma4LaZrBgzdGIWfK6W1YB+9vbVqWlnFvbAETbnXrw+Ez+IeTY
kODTm1KfgRiAS0kWkDOHwGuTUOQEyA4klE5mk8yg4g5q+hAcsWNxEjrJn5nxvF9PnKlIt4/ro7uU
1t0/BCKqOBBUWMjFEeO85CKIy3XM5LS5AHo5jLCXL64YNSTNcQ26L7S8detVZvQcGw+mcFN/GW7U
mEeOgTfhvXSgv5pVJ/nErMhlumrFufz6DiXzIMVUPB67gtHKOinwcd+3OZx3cBpS7DsX+yXgbgRc
1g4n2oaR7LkhlNjSA1b7hKdbiP5ul1/ZTNLggr9vYevAv4gXHgG1BZ2uFyrdqs05HnJxVwZ28S0g
v2SbZmmGEz856kgLbNkdkKSgEiAE5+59dBbncdvF9eSTMICsUkSIfS5vAGEMB7qftOWbDk8T289n
r3vRAKSGim3wYYRr8j1mOJqRaHP7OtoNvvjYHpds5f87n31e3FPHiOSOaUqGi3uYF1NwbHMo4bsk
dPrFoV+aG11PlLatWyP0hgLgXGiuozKDJpOgdLZtrvjXBN0lc6Bo2fdyNNV3oT8JzuWITLTofL8u
s+O0Ca97ZS40N3Td9SF03QESqK8mGWLeqFtJTJClht6Zs4+BK+8DA7hxkSZLy3QTNgqniZ/y84pR
4+Sf2R5BSVNIHER5H03mr5jgvlDbLSU3KpOzQT0OTzsFVGXeVoX9Q4VdbInyZsyCpNIpd7PEm38s
0kd2zXqSfhR6q4YADBdGt5mb/cIxC1RWXAmDfRRjozZh58geJyCmRq1fl+YDQdAswIDyBFOvrjSn
XpV21o+4Zk5gx51+nDJuokAeDTUG4rDQrPuOFvolxvOM4xPGndKSL6ky2OW169y7UQzSrS+X8J/N
b1plupyA6k2XVVKOreP0ORFRB/1tTrJN6+KWB92Y/1Tt/nSL653Dy2WUNgL4FXSCnMPy/xEFIcW+
nr6zNSx3k8ezQ+Xke+CgQU4eWLzJ8umr8eMVhUmJwNC/uBmH5T7cMwLa+w/rqUy7cvAPLXMKcrY0
2lSqaagx6KMK7YomdMoJAvQmcIy0hWXvt6mH13YV6/57WyRBH1AFXQQFyfEVAtDGzMkn+KKpRNy0
EJEx+MsXbAUJRprwMCBkVdz2LRLT3jzLETnFoHq06fbgLxc+/bNVEklAOf85kKco6NXC+P1viupe
Qe9oBZh1NzQg3dzmxMXG3exa6SFfGq7j4cnJkiXQgdKh7EUmTwzZg8v4SFx9D31yWGf1sK4lv3iW
Bge3nx9QOBd2kDl+GYiKHod9IK13/h3QHEtvNJ+ySWVVoNEQyVfwAQGD++CZY3+x8XPpBCIdZy+y
e+LWKkhfv/bo2aw/uiSflull7kpfPt28i67ETscYojGcvOw8edE/KrC1GJ2ZVQ/IjthJ3dxfdjA7
3fpGB7tneMUXBtSQUWE3dcW489cWnL3WiWC+IxwTR9i/S7Cv0ddU5X48iHd6XKnkEC4ypsA3NVxp
ZveVad+GqBFIfR3emylVO5BTRy4ErXRrpHXsbudGt4RVIj/A3J9aBCa7qMLA5+IE3DMqbWRop2U5
1illvtuTlk++YOcl7k8KFSg5pTXvuzECPzfY+lHMmT9+yYrgxwzyI+CWBgsvjrO4K1lyqr1lxmuN
mVBNJVPLGoab+Vi7si5mjQg4eGLxHXIsevzVJk71zJmp2AyX9NQLVaC97TlNBLFjNP+QlWn5YPph
FuLlryMSrT8uwlC7B5NWVHs612uLr/QUCW0C8uZezLWPq47J+ulKZQNP+5SmtjqUQDix4fu+nNgY
TT+V38leoQEu5dDBguunA8tLv0qgS0bDWLbK1vuIha7Mp21qhFKQYL9chjjG/s6nxKoZyBdB1KiW
yOV4Lln45xdJTmaQgQVwx+5WTTFXQeY85IdMZM15Uk0mfG5Kxt1BTm7hnSQvf0VJx3paNL68zHop
HjDkRn5odw41ZuChSDLSLgqEhV/Vr+BoBRm6PYTNbmu+jGx2IbH52JNLlYOxdSAnfcmyiSNUbjXj
sIWK5LkQu53xAqu7LZmC5Ohtn0htlbRd5kmUPbZzzUmNnt9S490rXqq2du5Yd31ZyXmCACbL23Hx
tLYZvdYYWorNQUSEftS3Ms2GcufRInrgIt/YTHnkTkz5mW5Mp23rIjnFe//NH/chGNKBQkIbvhIF
cXe+gjmXPrWfbNWBuGqmgK86XDzOasQErV3gh+C+FWOWKZVZ0tg4B8u3sPJBLsThobbk9ea5N1A8
TW5oi8ITw+eBXYilZqFAUVgkIV2xWSsQJHKixRfA7lreTHI80sF50VzcQWSlB8WvjSJzhuOgh5ML
4a/ysb9ExJYtDvShYStimwPnZ/0c0/6R3cBBtGC6xWd+OWM2mXK1shVJpmX1aVet6gKpMQ2p2QRZ
elqfAQO/HO66e5sw1YMlJwNEdL8suV/K2vtEebsTSKTFCZHRK1lz89/lMz80AccaoVIRJHaJS3Nm
B//eJG992BwyyH1Bs4MzOiWKUrWzyANV/R7s3XQD5EcDPmr9LJrHUGz5R4G75U7taOxEUCTB0tmM
ZbxD0bphHRXeLK6a2pp55Ze//KgkSMh5SVhcmpxu8rzZPBZnnXCAp8XbI943OL/rNH4bAIdOma+d
s+t6AFRP1q6E+Qo8BEqF8T6Ntkq3MDSuLIPEWxC4YoOPCpyL+xMUgekg0TL7i4g0bhan+Uen7xfH
WNyeAVoyJ9AyhTsnnBxwXHL/YA03AFZPt+rfuTx/G2Qs8+ZOW1I+IXjfZox2bWS+2qLzr4VJUEcw
X7OOPBSXJJjd+l1dr2u3Q3FONgc427d5yV81CYB3w2LqFwPUo8mlre91qFAL+58iDH/98BlLzfQx
bnmMc2E/ehQzFSNZ9rtDN/UXJiZhPoGKUw0ZMBbj0svjUkScsGRC3CZYuPyfHL0ee5fwIEsoKZFR
9RG2BYcNpn+GuTuZBuY4ujauC3TQsj40aRrTTBprdaLqoZSEvOjNflYPWPrTZl9VBYLCPy8ZoYrm
QaImcdf5orydNKbhzhcwKQ5mqAR734g3ic+gbQtfu0FTBcv7cYl7YuWr3psvjDNWhC8/eptvNqe/
Sts5Fc0riivkd75tQ6MB0WxGg7a/ttX3FRx0PELA1K2SqFLkn+CUxfLhYHKgdpPTgbrAegy7JgRp
lNHvLO1CU0XasIja3ZVQ3gt4RyIj+QrtZqxp8mkzN4EMuT3+kudUzmtlE7Zb3HOtBv7IMbYZ3JMs
NcFra95nCiuqFFbSan9X9sW+iN9Seio7BlE7ia96DvdjygT93NFYnvyQWkxng0JIcZ1kg39mlhlC
tATSUdQYgvV/HpPZd79GqxIkZOHqDDuxhY1XFp1bZtHhOGqH8LFf2RJAeeKGUQpgBXsWOZMdMGCC
2cKA7hzSS1J++cSrjCwA1+o6mUmlKptOc5JKFiWqdRVDuiHHFjnjP4syd/vFJB0Ja78ybC+rgOad
o1MJJ5AiaO6qItFnllVrXzc+DHQA3+qryH/K9nhFCIQnvoMFHyhkuRctARrNBxu9V5PeoLer27sI
dyuUPbnzX0EDeTPnOGXlrWJLw2YsrHhZUkq3j2CGhIXLkq2P4DHPE+0KwyOGEKOZpmKip68b6STC
B+Ng7kUsHdQ0qOu03S+SUR0TzSCUZnLghG+hJJFik4XVMcWdbyPY4hmhf3bB7Gg4u/YcntN4Q+fw
nQy+uzhqqgfd2B4yYPi/WF1fRExXrpa8SRVRIYbordgS9PBzHFfCBffe1f+x/rqCaN62GNK+yTSk
JnZu5JCCRB3F3rRcCkxsnBUv8ZPRmGonenAya0KCqZti5ury/knzhVQ6EoYsWw3hL1M2gtp9FRC8
85LZ4LE7qLbuGiaw0LsCQgPYzMtWkmcuFm8dt9/iQqX0zHHeAeu0ou1uQTdD/2jmBtSibKDUaDgl
LZj2BmWBi52z9AZb++zGa/xENfpL+8ObOIgWU5yKDRlYfFua2fnA26ZbnnPVHj+jLNBIMWb5koMP
l6majZRoZFY4HWeeSvcCZqaykEjtBWE3ejCau07NSRVebOEJTO27xz5Pgz8/SI9J1V39SQ/MYQ11
cd8C9CGuw2wrJQPltJS/HpleKwPnR1Bb1YPbaAm3WFpMNmtzmwwYL63m6hU7uGp9QJXW+7ZPVxQk
hndAuICaNEzr4rMem7KHJLBKg82cdd/S50nTWM1GInI164/Lx6zd6fvBclpzXAvC4BHKg0ZUu4nE
7ATKT6FxsZIILilimKwG6xxcBngOw1EvEx6W4kxPa8U1YNEVLOgHbHHTx12cnLXlaQtsYkL6yh0z
Bu8tuc8+iPwb4hZTkA4D5IDxEXpO1EY5+2bP85Pk9BI8MBJ+w5BPftsVhG8y60Sqh+UQ7gFbcvq5
92B/WdJWx00IUf0nanNSAZLdRK4vlqyDc34Q/UvQCLaH/SABJdfeUPgWYNhzB7zUpv9hVeRbDiP6
AthsEZ6ef68qOz0YXZoCn1e+z+UUQuaGSxEkioEzoPp1uD5iK9dxOg11idyk/WTjnVKHcoP6d4HA
3DQll3Y/cP4mrX2kNq2fIu2zckKjZ2Eiznp6XCDqH5fFqWN1pdxZWTTHr0LbzbHeWwhfOzPb/hwG
na4imBv4WVthXFN9I7eqp1ukxRRsQIxximieuV68U7PRWLuxbWqCAalzlQ54OzorKxsLrNp/JqCS
hzrTxIwVB8ZzyLOksooS7Fu9UEOOVDkjbT+1nvKu7PYNl9V4PJFKebXpgo6bE+rSGLrzUgI4sBWO
AkCNnUA6ae5laa0qXxSR0UlQTp8FhG2BEZ380+QRuA6qIyLg9wEaHW2RKiAf85ZHyGPpepGwvWv1
wUjM4cbUnRYxvn2K2arOo2c8Xf+pK9d9gJdGsUph0dDN39/n/8eC+oro/gPDNdlQ0q3HJG0LDBtI
fRfa51dbWN8mkkHuZVt6k+1vkEM7LslNTG+GDQ8enRuvcZdZ9jrpftcZGgaqIygmdI5e1qqLeSJy
fOma4MaZCKC0vmVqx0uFcgdVZYF02d5RfHHASkLoU3dkH5drhxI+13ttEE2ogwASJX1ecRx6CgJV
bLK8pS30GsQaXm/YBP/Izupc0YyNkuWOmonnSB3N6AQg0bzbI5MZbXz3KPIhF7nUND2OEswBzSJ8
eS1iOF6zSHLXS9lII7kc4Tfx4HByVIYHIXrLZzndJr7QkyQI8dyizzmp7VDyk+uajIN039IERsbA
gjiKuhQrJ2Q40gIIhcEwwzd/5xbbYR5952qpmVcqwNQOqHQWjaVcEYKqWGkmlMAcpTFVL/F7hER7
SD3mgYL6upMiRpB4IzIlxI3ID2nNK9m3scvJXdlUzvZlPZNc9tR5GPk91YW+zvTZvEBldZuZnYfx
ZFR4XsQ5ohajHt4r3flhJmFDUhy2WzLlllxiI2DyXRgKC8IGLYJjjZbIvIMeV5OBx5AZydnpa4Gp
NT5ieeSRHuvU+bzeV18+I/tSHL7k1vqRaR9zVSKuU3DEN4gfHAViGI4Z4e7moewx9GrEmzdMymsH
hbWvl38/GVoD6wW8GP7gPJ4h1WMdsEskCGZT25W9OWgcys8s6IZidFtfkSIwP8QfJA2DZDrtsBvq
pSQ8lEZIU06akws6dEmg2KAVL41wySJTHK8ophBFPQwQOQvUFqivVNkFJaOz0mKqk1/wtYL0mRuW
6Z+OSvYEmrzlRlsm8UAoHSjdyNV67Deah3iFHio80n4Iv4I6VswB6heoi+q6UNaPWfeZNarffrnL
ItYDTeRFoZqYkhnHj2S3dOIUnH7wkBug5HTDESOT25r1pWcancDZuMSZK2waTqqiSyobtjIvFKu8
CN/j7TerHjV4W2D/xlaFjPOC9FDEmvtHWw2QjNAkaW5/H2lnacwstjOcr1w32GbylTBiWVEiJE1i
amw2A9HmVaUN4hfZ0YZO2ZfAWu/kc/7IF4D6bTjmN99++esgqCQ0cyG8X2GbAYAzZ7lqXh+Hs3B0
btFUD7XTdiIVnnpCStyotfg3aJO6b6vy8LxJFTmCKfkuvSelFuL4G060i4LDBFcr/eFSO3Zcq/87
Rn+NN2rGRLa/TAPMS4QdDlUqq8zB+Efb3AxcKKrKr2OF42eZ88FK4adI/SHIURi4u8SerWPWtJI7
q5vVPy0s0wMqMTj5uizkhTDv/uOpyqolyHTbPuqjHps9wb2U7Bl2LoSuUz3g7yCzQ7mGA67gdApb
4yAWqJLVMX/ONshoJU9VgJc+buYPS/mpWLQ8TykhU+zQ/+qFz5DeON8IP8AY02kDy47OTyshbd5i
AD5hmXbw2zImM8qeKTfeyMoWDVSClHweD5M/dr6HgRriap4rmUhQkQGIt4H6amnHsLI11okT1Xuy
2MO5g815+yrvJjqo6uFLVkTjOsuS1CIvMYfr/8vIqrUGo2MitjdCHD2Mori/e0hG5eo5lndLVdq9
Eqq1bTwoSHdgz6Nxy262kRshU35jpTyn4Le3yg0OuezF3miAkpQh+c06++BYNlKFlQfX/96JYSb1
5M7uZh8otDJng8bN3NSFu4/0LI+CXj3GxUWyHFF14+zE5Nsz43pauhdhaA5CVASiKMPVICw6gF2S
Xbr1Lry0cSbF7Ag2EVLcy2xr9mXLrbI4bp50dxUtQ5oWBWpovSx8lQ5bSL15HS6BOzHsr9sV5uzh
qi29haSm3x0HWx0xRI+92iaEj/DNmWuKOTOG+vgsBrdebfXgnoZNTDjluQs3XcItjXCjlq2ggUeq
+cS9VbFKt03KYkHTOJ+zRd5dxCknyvwlUxYEetSQkhOov3z0Mb3NUl/tLKtHLkcbcB9G4A1QfpLt
5HX5kzYNORKgU5AiCbhcs0zAOIiKtSglqNABErxsbvCjyaOsWrJzaAJm/2Nxcp+B9OWUenQYKyxE
gaMb0Rqk03oFNHHCO0SwkqRsBgJM+IgGNF9vBtHJxBfxzDoikUPgswZEswNba6NoR4+bCkiREVGv
oXNd7JREvqZvGTei6UrrL1sPDuZ2+qCgOTt9VY/KqMctyLOePjKthMwTnez1l/SQgNV0ZSaUYiN6
DTON6fJZQ3DcNXWNJnaGcNQbnAoSNgoVIYC1SZZRelsQ3/fDCgjXTDSWIdqVsJMhfBysnuludome
GkOBT7eyiijIluj3Qi1HoLJkxqhZqJC7zUI4AwlschEp7tRctnstPrJQyDc1kJuZFs32Vex30ZF3
fKuD9V/LIqKI9lnfhVslV6kBZ8MFqnv2mwSg5wePOvgeffTUfvQmku368nm0fSfG5uDYmWzGSf0q
Fcc6p1L+UfUjA6vwcCqBuoZWEKNZPAHIcLuF80exETFYLi4aew74yV5If52WUvKBIAzuORgh+FGB
yu9D+G8jhZEoUslRdAwRt9v/w5cPFU1VZRPQxwglsjXZkEv/gHZ3blZ8uhBHXUvbnyM/xiZLEKe/
6pTZCn/YaJF7sc/Zlwd7/Oq6gaASq9lgFXBtZXwY1u3DpJQExEDJj72hmN3byTqcy5oLOjmRLOMI
BXov4D1ofKO4OIvj17p7SaFH6TRkScrCSJd6FXl8K4CQ6SGzjPJ48yHxYVX/0EhGFoypqjYWzcu3
X6lNHBuTYh8hnB68PTXlUUl7q0K8Ovgz519pLlpf3J3FRUxBPCMxcnm+Lglj6SDkKQT4eKrryXcz
ustsKTCiVhSFlo/2g4nl8cXO/5CeiZUdaVGkBTZ1a7coJCmjnRvG9H8Zvhn4yoTrVWsFKoh034nX
ocSy5oE1N/ZKHmw4H824BBwK+kUdOR4oF/UhmiS341SurekHxgCCqBajadsSP3LB0aD26tbWSeCg
6KzfOdSW8mW6YWJDZ/3W3xA9yqVtzqmcRMsGNfZ0VsD3qC2Sxh7dmq2PL375SImffAycXiH5slr8
vI+ewKuRd1MVLOiVEAcVGaRiNJzvZFCWhEoU5I+2LjQMDRD4xAXXeXXfLzk5ephD7wfoEj+OaUA3
R9mlLKwCiDj3KHRneX7btKjQiU2k3iGiOR4n2XDRUfwbBKVaVGRScIwv2wMF8AnLgAbMcF3f9qrk
KPq1pZ97cx56H9/Pdy33pN9kdIMDjpFEXW4CadbL0MmqZ10FjsTjih3BulIST5aq2umfbuKMxLTi
jSBY/iyI03xH9Q+KtqggqsgbVabPEo0SW5qdwxR/3jsVsHmB2QESnbkbBDQbAo+B9z1U30WOlquY
OC0vd9ylhNmtSIQiQSTezbt9mls5xWN9oEzgZLI4hnHmXTc1A8j4KSUiZwSXyAbqPIK4jkQRkwYI
VXlYwgKiGfD8SWg4VyqJLySM60iF8ZQMwgZmFBjRbcCTkZ9xwgfVGqefFksbHgaaN2BO/OoCfXxc
bi9u1msP1o1jgDbaYDohCLcONmFwEFGCAlut/iVDzYxUZZ2anVwzNdRSkUnHsriZ5DKHgA7HW4qW
jrfdg7fOrT2qf+9zAGi3S9WtB63/LWr2X5I5fjtPjy37Non24czXmdax9OHb2DFEfLTtNtLyNXO7
69uByCuY3qPCAjxUV4GYs5ha+hfrGbfu9eoSotYmnZoI77aCSVNX46VX0jPJoTYJjEPKbGLqSfh+
HeCJo4UudRxrBX21lxumzGfOaX4rYR3SurqEyPWl8d7CRMJy+EfErPoMlnE10eYBj5SNWX+W2tB7
28Y+MTydk+NXAjz5Lcyjx7dsH6OM975yNMC8uklOmfsnFAqkUw4bV9pJzwub/NFkFjBc/utp1+29
yMC25sqExlw2HPsTIoWwjX8a+l4XwI/vJtXmNQRyavReNhDiz7HQvG1xXH98DE2cyFB2VOqo4pdt
dU1AaFtHha6h9XieOp1kYkA9enqHP2tLBs5nL5YLhEtI5Tedj0fj0OzfMm4VrsLHeObItNylv4eh
iO2SHHMGP9eE8R92hdh/JVnVGuvuU9B+5oSO59uTqsLKfMwjkBQJQkC09oS4SdjSIKTP6nXbou6k
Ybacn1LZpSnD2PGUrQsG36+/B/xgI3Vh1+j9nASHO+oQ4Ng/nW/Xhp1m2mJDqSp58FWrD/Q7+QxS
aKLDRaQEUbSrWuJFOfowJj1cf575+9BeXKD7q8JN3fDSY9RVZ4fvRm9LHB6kmGkXobqM53t4TkZM
gQgL9jz4fajj1TPsMqLEPFonv5BLwJqe6iMYLXmjVL0sHum2sHeCEnapkexTbc2VFgX4qa4zvf4r
4AK+L8fJCnAuRqg5ewEfqlmZ/rJcOa2Ty7veyfdeFq2ZyScIHN5Z0f/t90ZL3gXVkvwybgvqaDaP
H4a1j2QSaHy8TOJeRjxHE3ow6oIO8nZa8mBqVdG7X+XJ3+hrvqytBkIB78K2D5FkiepCSoVigGBC
MsZlq0EdpGXVFbZbEDozmUS5fYoZZ4AG0t4G9L60f4cBSGa5iUjiy667pVZVTddxDuXokkocuUpR
9JolwBaefHkY8pnsL8TLBu63LcJTRSSeVQTv0UGZf7XU5CFS2q4jbARdQ5VbHYcCkeNwvNySkPNr
BeqS62+wcfT76BKrn3L8BRP49U1nGpr8NyHvgVzNYNOOorAf1fRWORF182PGnHYSXPHak/P+KvMZ
wLwNSHEiaWyID8npRXIhCh8+7H+UrIYZi/83y0i4oe8X+CJY/bTEHvsmfScuvc9nrqQxlezxS0lR
w0ThuNoPlFDTCIdwf4Xq2HatTs1yZXCfHUoUpJgMgrhkZjS4Wy5fYOhbXjxjflQtA/VKzoaLoa/f
pa2XqTfgxPXBHA+a116S7yWDBRpTr9y3ohKXCXETX2E/TsSfFDjhVT58HhjPbVIZXOt6tUD5RCND
1/O8zFSY+mVaXFou3cYq9QYgC76DEFGzkJXmOJOWxGMyyeY/vTI+vyDbL2sQ34CKfMY78ycnrwMe
9GbBA6VxAJfB/cJIk463hvhxmV3+tSY7aTNuiaY6icqBboro9gOxCl3/H25J+kcWCHJHzKK4jrUO
ZOOq3h1ySepc1yRGm06T/jtRF9UWoqOZU4nsvofX42dGJSDGvd8GmtvjP9GwGynI93HggKdgZs0n
4F/bqi9/lwnlLL0Dl6KLVM5PHTDabmsiiPB4Emy3woRNPYuIGt/GLI7n99Z4CFNbbetH2hEYabCb
qLNNAbM4GQErFOSKsk4Do+ryryLUPNMvxnTO/fwlziQgiyyFkgH2Norwit5askvzgE1l4RRWsuui
tAgN8zNzkiqL8VbbePDC065WK9s4Q6jEUdaRvL30am7IUI93KZgnUnXmblcAcPlsqUkL1xsDQWkb
8V9v+rgPGKqfhsLsMVjzeWwTAb7DvyhRxR/i8xluG0wGQI7mQbmK9m/IN2g5muuA2iN9S/VXEZsk
gjDzzSgtQkCtNNYPoVV7uP0MZKKHalnkmIuJw5kT4/aI9dOnR/ybW333N3Y1hyD+4Vab+qnehr56
KdBN6ba/0m17rImbC3kJLTl0kJZ1HeUOA+fOA+GT/PQfjtM2K71J0t4Vy+USbnrNgBay8q2ZCQ9c
XRR6YxKjMPnzw1D8/6itrw3V4YsItyfkfd3YTbLWI5Ua8zc/8in5nqE5dmsNV7kd1Fvvkt3FWXA4
G4jfDWlg7Vu0W2dVvSlSToS+134PMoZfFui3rEsQ1RD76PMhL1T7ZWxQXd0THGpKRDEO/kAO0NYB
A5RIBgVXbfh3KbaAuCdlebNxwVAvvbesYinmvbLeB9spPzFb6AAEu7dzPOLCDYvyOt44UWPbJynn
nNaV/4eQ2PPA9x9SHo0JLAr3qzWgQdNgATT2RkB+B40NlebqlT8qhK+dsKZkIWzK9Gq7+5KI6BEl
G7AdcePWvqbQXGXWKAc8okTXevmi9T8xbmT22rNJUQi//4XSdyxvQHLz9dU/An03ek5CtHqA2BH0
tdyT+vHV5ZWnBqGZ9XtwS/RO66YdLo5SKjSlmGH16TmyYw10vuG+5TcqnmizoOjubTo7vzXrj8fC
R7CV7Kz3Vify51qrBQOlaAjgNyD0xCEbhRv1wfqF0yQAzN7cr2tBmppg2B8dNFVJCL8mYvDS80xZ
QnlQl0BQp12zUOWcfDbUYCTaQTZ80jGwVdRMly/zrZveEtCXHwfpSJ4Jt3NMYjcoizZ8Kb1ZKfBw
CMrLZt4CnFreSETTFY9ZsWa6D/+kNZdrGAwORY7GpwvJfZB50pvQAxf5GJMPefHXiuAqYZ01SSq2
dW8gXnXkIUwHyT7NTrY5dYSfOovyjPdydDmzVKiPB+yvf9DmcZ5nMMREAJDSBZSp/tK/Pxu21s2C
Bfkvss1C8SmCrRpZxRoo8alA1N9fycFMPGnWYRBLr01KX4n+ShvDSU/0zw41Z/RB0bWJCpQ94RRx
b8j2lBRfYSZjDaijIXPU/ygCulaP8MKT+rbeVb5xFa4MVfsrPO4EH7JqBVR0sJZpdoUI2KtoKlfe
n1+mHjWnyIVPI9EBBLyFDHmHo5MUJrL1/totVnWvXrOpHf4yaj7GfXBejgK6LvqTFyojWgXCG5D2
f+mrSkHCMIb0sOZ+fnPinUgQRTM6asiFOBMQSGPRXqXwslAO+Xtr5I5LjRwrfa4vY302s06xqVfE
Kool/QHfOeg6jTVc4fHHFKfG6qdRg1Vbb6eITdluscLh0wO6qZ3xv7Pw1B7vcMHisA3cMnjhRW2I
lNKmSERjAwbYXP7s+Ov7Lkfcnrn3SZYArUKKD1tvdsf87G+xWKuT5aqJWwjl8bfyEXsV98CNSP8P
DLg4tkH28VEMdoQ1/eWLIPheYoPBvEqSAU+Q+7X3N8Exf0wNNq+iWVV5VRL8Cw7YHC9CFJl3YRi3
DZo8ZU50Fbr6rj4kckuW9m/6eNpSKJwqOMDayqZJTMczOsm8hhCI+C+uaNnjzhOG/vrM9bSMkPLp
ITA6ifBfUOtdFmZ7RvuYKeIaNdFvybl52P7I0HchQU8ObagFYUt2uqXBJADWlSYPdNiUisOrmWGK
qGxAccdFxqAriiwNG82bmG1geFlUUEBOducHLcEGNi+YfgLceFfXufdSX+5WFb4R8qvcu5vYMU8g
X4eO1qYHG4e23M9lbggseDbWLSZeJa1ztFsv1KWw+Oxo+WcindYVvUD2kuraw3WwLLAi2Zipf3Bu
HDPRIKUtOiVDebOQamBm4todVaZ4NbOztxIw4zEMO60oN/KIawHjcyTZTo0K5CpjejBSJ1pyUEzK
abXdB9kAcGmTngxvD7Ozopw/7S3zU3ZVEf9lyAkPJrPo4y960bc04pWuKv+KhjSlHgHZXqVHqnTA
sqWgUQD/M/4l3XXUhVKH/gYoNA4bGJe2JuRRY05Nb7Y4LL91CorG+PdY+g242kMiJog4eBcD+V1W
gO93NCsD3VFFu03ACwhHXedrASY77R16scJLCpxsOQS+5oYMX5P9k+ptmOkhHbh5GqxxZQ2JV26n
DIvk6+GxCVez/QOPmVtvzCPp8TARTYYc/Z4OFK8hzXb5T2D2cdv3+SSZkf9KOj9q5LmBcfwxdiRO
gXInaHfe3wBM9yId7W3lnN9oZZ5K1EqdaMvHFLDVL6gqei8Uy9it8YnR9uiCHf4g7QAnE/WYsdCn
McpgdLGnwGyF3nc3puONMpj5tDHy8gI7U8sAlRKr9kNwOnJgvRglkQ0Hir+VEirlz5zFIWGw/TlJ
pnwROSRUsaeImamNgtz43qyznwvqXoC7xqvPQAqWOMXv8iQrbO4cNKnuCoosmx0EMVNce5zljMMl
BAfVnO5yzmcpoYbRbS3BPmIZxIOqnWCDpXl26X0/NpWa207iRda6eUIbpS6BgczQUXcKK8+pD3ag
wv0B2lPU/1S0KUGsVX8gNfydJtegtcVffG46DC3N7xDL0kV0+BfcpFupo9YB3BIMEdocbQqJTecR
Ll2cibteLd+HEs/Av28uT1plIImlAegBOuvFgB0sNx/5/wdao2bqXMHDxnsrmAKgKaC1H2dY5c2Z
GtNKPK76InvcQ4oBNOMc2iqq3e5Q2Vh/KPlZcxwJ3RgcQ6kbm7baNwJvfr2TfnP4JZlKz/GhPyEK
BGu089YXgG8FfQvf9PmWDWjhfT4cTaQHZlPqFPOzmgCTycqbbqQOeGbx0lIis7I7nxihQ9J8mmWu
xrFyhCYqbkk1OtQzq9dFBOIEAJ9OxV5RzC7JLgrR9rzCZiJcgndlTdVa/OLK8DxwoFxEhqCh2SoD
qZNQoFL4oo+/dpwEfIR6W+wLpzP1VVggkexlv3HGz7rHy0V+a3tS0TGjmAW/Gat5rUW1JZC8cyNO
DknsjGmeJPYY1Jd3gmc1/FqPAm0zRn1Qjqd9AQdXiMORyC85ARtWhgwZZPRP480K88QTImnlrY1T
M1+f91XFTl6RkJUAP+Xat7pulqQbfGKUMu2fZCB+XjCEVpwcdfBmqNkccmSce4KktopWeeVULuec
ILjsaoalHyaMI4c+7+MfxGfj/LeBUTeEj1n2ldKTsyzAjqAHk6HJ+g3aSx9e6pW4dXSdtjtarQBu
2+ZFRSQXNow+5waNXdgm+mBiTNvouemm6KqF0/g174u3D/WRle+wFsieY3f7mUsoIIrOIAVNjrQe
/m1pnYx9Dx7rgeefaMuJNZa5Ly6QUJum0Q+08Hx+aNaM88DF4BA0D/1c/csoEaIYVPVSjM6Oiu2r
XLCSa4EPhCcgQXjQRBQEIpkax+Ngx25C/HGMtApXy7Pc2y1464zjfNcy/IaYl/Fkccdl8eDvJ33z
bif5a/so/W0GHts0+Y1a1Gi9x5k4vzm1U5L0ZMSKniaDNUwfVmDV8NJdB8p39q6h8p033kuNnYHm
T/Ia9uTDnPi09fGb7OOIFxasI2zazKKzURkcBBJEdqi6glGgFhIM31oW6Yj5nIZrvV9pvl4Bl8Qd
pcatCZjks15Tl9lUTwdqPZqd0unH5IE0Fq+uEBv3HLjExwlx/Yku86TdNATrLeSXnsT3cJ57L0pg
7O11+e71Ufm8Ii9Jz4wm6v9wHkOSVzp01dO9eMPbqNHKAyK84Clgs2LERDaB2LBqZdk10diQ/8U2
3FcszNxkwAeHQCZW2HoHeVakRicFXDuJDzOq30SnSPDNL/WFPPHNQTGwZkrMr3wysw3B+1pm4J4y
Trdew8DIk6XPX8N1HTVnpeX/gCP9ki1bEk2XysZCcIgoqBVm2SSHbgRXXjwoyS+8jHcu7DK5Pckj
CUX6JSO6z9hg022bApLX/ZJJK1jcXLS5CftsI5hZxgJRps/f3TmlMz4JwimsILdFebf4ovVMgF2F
2nxAxntXPQjcJh/Vxb9SIJd48uPmnTegoDjOuG++hkTv+q1LhlnnfyBcCYLCz50hk7egydmO68JF
VGwxPOlo69KGb7DbdatUDCUl7XOfow68KFdvKHLQi6KncSwp6Bi3Td/GTxEjueNtYi5MCLDYDiqx
Y0RCbIYkx9XPnvsytAbOnztOTK/XA+0eGgqZLi4vqZaN/K+0BEp+bomhBF0vyUGQlCZq9slkrBjd
eKwlZTFKcKTVYJoynJGAZYs6gMqWcZDSq0HDZ2fec1nNRN9yvxEwnJrK+lsdPF5bwjQ6Cy03hqkz
kvDLX8fNS6kmV8rxgotYhckS12kLLSJ/Ge2xOEA4GfUQeCmce863yySHrBY+rhnbrNj3D5csm3dN
s35mVi7J0b9T997bFqS2NOu+jfdBdmTSVjY/+dvlkTtjg/Zr+tkhePbcbzpw2jILoYjuZ4VlyWe3
n5LweeskacqrBAtepx2eNYzrghbsAdGokc87OqGusRiGBWF1W47MIQCZegV5lcc9UMICZyV17AzJ
hlO+yZtAhmzsB7dRyfSWw04rPCNsqWLlJLV1WeqINmx4DiYpfJpIQewDJyPN1Ii0CqdG42GIp+AS
b5Pov/oPjLuhMouusx1Xez5WFeHuPTXBRQDbIlRLupi9Or/xozDf7MGtmqae7eRL+fU2M3v2QwLq
OBqcdDqgYiuNIyD3Ozh53QhuC0Sfil/1480wbXupX7peb5lFc1wLPoPEbPVQEn1QdWevqPb+F1Xx
Rrlp8agGqPe4QCV2Rm+lyfBcShd2NsrXkU6Iaik/ah43zGCVe8nIdUGi6dBM1TdgkR/6c8XF8yf/
ubtwMhTPQza1nVECmAMlAPUgaLpGc2Zqubwxhh6vb8O2Bxj5DeqIiPYO6tjOXmZ6oE90QJcutIMD
x8deYAcgeDm6Oteih5uf0o57F/t2EZqYPb3CTWypjW29kR+9M1AjRG1dMwPAUbNA1ojdRrnImAYO
YCaLHFVpuOYkq13a3EUq6KYXqkycSviVv1OPqvY1pm4c5HdlOhWn0+b+SwINFaDBpl7NWQBVH7p7
arhuTFOhtYPnD55EQy5rDTaZyFVKycwsUUZP50BIHFQSYdfNY+lDoNeWnm9XtUs+Afb1gDl69/Y0
dfhBkOGkiv3j9pno2icnlE7zQpI8TA+OXMj0AURsMUDMXJOkzkAou8V9Zr/dQNkjPTSMVUHbnBXg
7SH0LTrfbKpXbKEXtOo4nubqtXoajG1AIPQMrbBbueGAys3xNWTl5HuIkq2uWWTRTrS4oDZ434O2
UwMMPZReoUw74c4S92KnMBcy5Ph55Ay89SMFsWVJhBjALG9c7mfkhKpTrYR9GqXJlPd7TMkdB6/L
RlKoE0bOcfuJe2QmRADHV3aPMzOzXF6dcgYclawVElth/OlhyPC3JGoZ92qbVc3Gau8M4KdPsZfT
Tb+75kuH6eUo/rHQjU36cvaA4gqsAkip3U60Bh+ZDN8AlW+s/x1E6SPd2ZGC7jjK5UNkSji0TR4R
KaO8T87h4csYjqDOkFC2CjMKgYAXNwhLC6qwdGMkVcNetRp8vySTFTrU0ywYHPrRv+yJZ29KOKb9
WXk6B0QOiVheTIs2kpf0AeRGcGRQcWdcEPRaJGmQ5ZhrSGXNseLdMU5OO+63qJZ5vwSBLZgu0yHh
qLtz2gi/UEV+b4gUTFWUciAh5om587bVwrOuxRlizsX+b0sZvR810TtHVD73YMMkuGpu6cZ+TATB
FvNFxFaLrNz8ZtXVbC+B8s/Fba3IZ79vjKwdBoWh9boi+C4/H9GhP4kZEk2HrnfCsND+Jlq4Ypsz
S01th/4wOiUofN9KlQxIIxSiL4qz4v1ZKfH/01maVZjkiWYOkl9S7T+PP97PxP/sFAC/90X5vDH5
UaSOUr7y+Ty5B8w+kJJE2fIuJfEzWOQp4nbg5amnIGXbBsP4isLfN4p6J8dru+bCBnz9ekKa/kIP
i5I8udZEEUOLGkKAYLPcBPZiBO2CRGsJE0cDzcI0udrfpfDwzSqcwSfjqc9xwhPCk/Cce1H5tL5V
qhPcc/NIKavJ+3F0a7H1gKWD2C5JRBQWX+ejjF2/XJzzFQ5xNqB7kMbdgjIX1269fOgzQ5IIILJV
p97+hzwowa3K1tybrqodvhXCTINTf+xw8Q+x8imJWiskYiuLR5Ei/HZ003yM1aTg5TLQdPxjFHSX
hCiW23shChnQbcCeKxeKnIxa8Mc4/a4jCKi5hblcLRDMzwJgVLrvPFdgo+77r9xQ/rGTMQftHD4H
QzAt9URLAxiibZSKbKXQbqUQx+w2T9unUq2pEvN9V+/rBQhYDYRxtcEVbA8ay1sovpXUfL7cV304
o/xQc7DniPelxRP2dfcnAhoDjT+xj5n5WX6P8Ay+0Bjo2IHOB0nWfiJHWgGxJnJbgxCyKHOUnuz3
XqGDb6EMt928tytlnSVj/j7Yd3pk52L07TIAVCe4kn40sjtHemE8nH2xAtPW5xDWBKP5wxiz92dv
gpZAx0E96nJNYwMZmGkHvoMaNuNX+KOWkNb4Hx+E24r0r7HT8yyOkV1ZhFu/+esl92Ae4f8/MFCn
pJuKmPC2Su8YfR6EEGKJrXtP7oPDU8x1K5f2nQwZtRB/VemRDQGJn7+0B4KLxDpsBmNR8KImKFJW
kwJ3lSbrw2Yp3UZzwXBgHs/XTMzy26xD5k3xVWyxjAcX4Vkv8f6znNSan34NWp3+XotzEOyYUPjg
jcK5m9gbJ/NlBwUAsZeNctaXfxQRyxJa9xVicNn/u45QIgfj5rhi6blSqu1/MrgdjT850lmOzY6w
CI/wuBKDS+TsrbOgsHl6csRlpZVW1nt+wNDmpPWKhd1WpUDkO7mRn5wopEKK1sIjTUKN2Yu+IIaO
dGqSbRLKvzjPHb8v4XCocARgto+HhhSGoyVpwXi/hvt4h5SFUdePrcu2oG/DC10kT/YCZyUP+0DJ
R4Gua8qd2kIt7HShQdJHnaaqrJKoSFMHiaiX0lmX3/8rZU108D4C94HAjUg6vT6ZQ1XwVJUukPg9
zrHdbpJPgMNfsEDGJDoaZ/DSFVCUxFBdpA4rBYZFJ2funOofOeg+Evu35m7bpBn2Cd9pBaa07yJB
0GrVjE97v1EsfQie7ZKQyTvU7+l6lBQgXuJEuyYeTNZwF3dFCFrMg7aVcGf8wEL6LhgWZtG6ntTx
NDcfW+cpl6WDxMt5kazjvcoYtf7ol1YNs4Au5cM8AENfEm02qUgCfbtdlCcPsUzjQJ6w6KKKRc9Y
DIWCrrJCfVoKdsMgZbJVUg1w+5PK3c3m95KLvDYtAfsAzswcsaJyDP4j06+UhSykUIQg5Ktk/iPN
QKUK4ECjcEgaCpBsDllBuu3X5m2e8xG+gRcMgBcQe4wktNBrbByXm4O4LfTyxQfoaz8GL4u/4gJT
02LAHE31R2ga698lMexCLfsniTM3jIDHKVm/0EJOPyrIFsza6gWrSg1qbAqAayxIyLEAWzlopJPS
ua3FqQgYpioKUqM0nnbNXAWNduD2GgsjwHpy81ob1tw6sTRHxWxVTsEm4RoeYiYqb73FDJrW6Nps
/Pp/zp7lsnsRLlsRnAULXUs72l+Pp9+sQWXyjgY0rEiMycu6TNQm+VZyRjWlWOJVykdLeMQuDdnp
L6S3CnWo/zzjtTdsMOHa0mRqvuy4a2+mziwUbG+H2lkta7LaedVbLbP5J7XTF9gY69W6pHxJ31js
TEc9KagEyyMHEHM+ryd/dZuZ0QHCxxLMeYuiL3r6q0xMbEOJA7+Mq0HH8imYgia/ALWOz+t8CeL5
VHdfY6LsQhvwbTlSego/TwTwophcAAb9mQY8oU3kEedkY859/EYwt0m0w2jJFuiWGdkYF5km3J3x
dTNHhPEs5kOpbTUQFftE9idXMAuP8tjcDrg7q2iGz23gRVpaeUPfdhxGDWKAsxZsa32he+5wu8XZ
e6ZZfeh75YTYK3fJsGcxY7KPyqAM/0Rdbo5ZErDsReGtVApEYPFK276NUAXWFVixiztVVxSRhgJG
k4ykHcHm33IX7I74Oq2/WXN1dlgJJQbCZIn8weCtGDHfuzDOmTnz1T2T+PYaQXXXn2GlbW5qJl1a
5/l8+VTCx/k/s60x82TPzhpFl1eEV/Z18cK1jnQv2H/X8atFQMbKgpBb2BxS96eZI3kpeybX16mY
K6JVpQ6PKAX3aW6hUarM6QsA4sY3xl9Kn8dkCW//DjD5VjNwiyehyjGn79QPvdkBEqaiQWKcJf17
VT3Ri1Bv7DkEqa9r13SKefBx38vHsz+Hs2WLCwGxlpAPaaUvK47IqT5sI77SS6JUeXWhVpMnaqR/
CasHjtPj3/R/jCpv8a/O9cLUa325FaXGuCBYkT8R216fga2uZnul5N+bY3WU37seoAHCFwX50MOP
misYzsaD7LFepvUNxNvs4fxA8bE+h+OSVP896omQ3fdOdyGT0hfDa4Fq1KsH/uH9D09BfPa9tQM8
wqub5M7y38woTgh2Q7LRnkEVbICa+zjSY9rF+D8kgODox8tlSAKcthlcBjfgLk13Hi2QV6wAQn2K
3qsbuEoRl+RUa7m+oGxHi0VRvAi+o2y+x5zIlGNw1JPzm+xDr4oxlhvNlNlvuEoDb8VlE/ZnYQvO
mYY1yDcE1ZjCC0OUSv67FA3yA00GhBDxO2J4GQOEJCKtHNLJRDY601NShe5hjXSXWGWoIE0PdZWv
YEVc2RwePp2XEIM74axKd0+BpS/BtsQWLaOqRAeSfXEvI8YgyjzJ3dMbXDdxjRB33L6r87OCHQN4
EybtZ+fFfZ2BG3I12ei+kdnh/Si9QGvfanGJuj2Kg4cQ/jQAbHCnPw7Cn37L7NaqjfrSoO7fGPCw
4chzq1yqJqHpVIGSaicNAKEbOCCd2tSNXGrJ4GrPGXpNUgInS+xNeFWsnM7gMtRK9c/BjBhmLzZp
JSKq7lqn5K20c5MEdf4YVAbF/yZ9AH1nO3qu7uR03NDZt07Tntba0VqOGFntNCk0pg4cRRtBRBUP
qeWq9rbto6qEcLZcrK4HUqeDRKc+tzfbTYP07rQXXxuK2NIl3cLIXaNRBTJ+QDett1LS8LYN1BcJ
OsoCR7w85WH4oA2tPNWUPUx4xzb5cwAk/tzbNtBawMxWAi/aF//JvxwnpSQHRCwGSp7rlFamf/nM
J5FRGk1+z3swF02HcHvvVmgPxbXMDZ3Qt41yKFzgPb08LgPIluwfnh6dSelGNZsB0o6g9V/D/jru
jbRP0AdFWOlGUxDmRiFE3GKiq8Ob5OBmxyVWVGB+qKq2fKGeUKaarxXVDR1f16vM7ko6ktGPXdG6
J3mx1MEA2eVWVxKl5DWlDEql4lh43xaNZmqPmrSQdQ+jsC05zteIluSmUX7ItMSXB5WmVSHDcu/t
NxWKTlaN17oM8IV385Xutws+sLWEP7K3ZRNMKefWgIu4eOKh9Q1DLG7xdP2YXdbyHYMGijsFvG7P
mAcHcHwFXAX8YXFvv9ds0qr5Z2OHV6++Xsb9nuJb+abWxpMyV0DqEMoP7JrKgEVAn0GNj8ksdy7e
6+blGufKc5zQVLkAJzwlRbo36WQ6OvQu/MEgSG75ZSOkC2IabPOHZjLISUvcB/xNXXNUvuxcQPPM
hjwCJvu/2sDD6J7BHbYKEMFkPDkaUQ2GPEK6g/qJg4FRoIEDdgb+c4WdVcCdKlxiemICwczB9Ln/
ME7KWLEv1FB+Ewjfv9N6BoAt0DbMaNdB3FQsdE2yShq/vhY9bznyn4Og0EeViQVRHmHXD6+JbKYZ
u3qmCUExRQp78S9u5SoMAFztxEJT+MQkMJUwirBa5jmI92d/7FVJRbIL+7Z8K4q4x0GhJNgmVJyn
0aEqr0riq9bkxm0/bZVRj01+Uflqdwy29ud5aqWP1YPKLfUoBWjKj56L91vD1qc9FU5iIieLEaX+
mUPsmLpujkJG0WDwUfihcUXE42Z6I8njwxAM8CKrglEPlhzyXnLRK1bO7qUeV9maqOI2YT4RU8aE
NOP7tx8hd3tCN7PzNyV4mfpidoZI1azS7QgYcBVJBFAAC8ifsjg9e35PM2thdgcEHPzvElir3jkW
Snqg25PkjhSeTnZdIgNVYGgpzQlhI+8N9zKnv4hTv69WeG1lF+ZL5Dvu+BBceA6cWusuXL7IUkOO
TystXcc4G5pnXIVJFQ/any9fbVMnT7G3NjIXOaFfzoUUWbPDqvBELyuGZxGnYmDqZkz6mxjjz+dE
5vKID9CdUJsGkzLebq0DsJWApKNskXr1YxbEjwAFqP5EW3ZSSDE0YreEtTv1EGulW5AujQxaHH1u
9RkJfruCIMU5CVbX/qYuu41wTu2/mIA/vUP21EhmhnGGS1DNiOvO7uwf+/LA7OWYcgste+Ea9SAJ
Z8U5KtkGbguDz9l5zVJZnIV7/OuDKnJF2XytaBRf8booN9M2+wnCdXVlxRhMf/yuRwHKqNPidelR
HVvJuNrmHfB+avXfATo5u3gL/+GpdUEpVtkOd+ynDzHR7vLs6EMd67ayKeJQbPDvQwF4Q1/bdWw0
HiqZ8vUCZDhnk4xqERi3CehgNyWZSNQ+2/elR2sTtRYFE1j03sgRWcnvXtSn2yRpkAEWVmQPlFUr
j9eJNSfhOVEAd2tFHCwPk8dbN/nkpDBR3QBWPkWGhSJpdjbxpYcHVsTHnCQhhE34C79UKqVq7Iae
IRlxIy5GstEaVMxO2KXRb9dXJyFs8QqMP3kkb2JwVJEUoaMk2YgSm0+rco39MS2Z+Vdf+32c3zsB
P2cVSa3tWeXfZ081R+QQUBS0eAJs3asSa5GoCIkMBG2O2yNpAqmTnECNOHr6Qoa5T90Rc+vLYOWl
zJYfXzn0C5rvQ4IPwM00xStZYDm2/RmL+a8X/31IoS+pu7YfgUYNvUlpM5CkxYVmbdbpmclz5RXR
U1QKRF0Lz00VRyCHv3yKeLpQiKiRltHdCgtNGTQIEocAHuIcaAQHdwmgXnVj6RUJShnBDrzgblkS
1uegiqy4DFQgD7rlhd9Qc4Hd0LwuZWOdLTp/N2BBxakoi3H/XUMO43xLK4GITvBiAE0+ba0xN1k3
ie6ZT2+dROZpKkeFi8UbI3FYCwxJQFCANww7XkDL7E+c29B6eaBxO87L4tCGQZh91Sb8dCADRzmL
nSMhGBDDbHbQfa5xHCU/4nAtpFfBjANNW0UUfUw7q91/J5R4pPuUsTlcwGstF9sSxUYknnuy9BfF
JTUgTrGtyIJSbvQEf4Nl2efK4PRNoa7eqxpL6v557wy3kBF69/P0EGjQxrxFtQuJ9lXDLB7Urty2
Mzr/S+vv4OmztdPe9NgBXWbDou8QDYWUp8DSgJltWkFg/lehMj0YRaajyRZCZTMYN1SkZqm3Nh37
Jx6t8keWlUTgXFxNhNqTdkHXg08m3EKjwkTqBj7tBMuhUTZi3kHlOLkiak//AousEUUSFtLLqiKH
T6IB4zc4NkG1Is8UG8FMXyjukkVU6jFx1FETuuetxMDF506bHhhwGj/wlE2MAt617q/7RSfR6fmN
N3905svj29dG4j5ezcxC7Rq8BeaJGNQvnIsh7oSzQQmXuHkspCno/Swd4tmJ3DHJillWZpJWLw6Y
5bAQcd1088HUE15GQxDUlf1+LEBFhuN/ra5tLM2508k6nw4T2CySeBJYs6oviUmdaWTELqygq7KO
eLZmIatsmCFOIhotNaY82o6GPF9dPSQ6ekz6f6/sZPgYkHQwaFBjUIgwdiSiDZHB38E5nbyige2F
dMofQ7D98L3vEPNeuuSdVg59K5pa9hm/B2bzlWqO9POjpRzWLOZX4qpjpJsrvANWTDYKdp+8xABD
6pGLX0mvdNm8okPiDA2cVemShTsjSSTKyYjncH0DErYbPisXAL5vaX5Yt/tv3y/D+Fv+R7RN4+JK
xvz6oLWFR/5yf0XvErert86fYVfF13koWV+EmPRYB131CRJat3Lw7GMMml9z7cS8M6XsFzjkH/lZ
6vUGswEAqfrsmoRzCHhvDbl/klG6CfRVH4AHuuHqlwN1S+vvVgT3HgkXEa+NQMTJj3BFEj5AejGO
Y77huyoiyK0oRgEOFkZ90w4DAjBHS0l/d9NMaPi5ITPKnJYRVtAbAp5ctb/WaRNqNGaVMoEjJekF
ucTNG6TYpcdU/5L3ax8ajPkCt2YSyC1W5xJwWDHHA3llcMDGtyTcAQ1NrgQdSEMobJy9jbdj6rqa
NcFb/IFFXN/WTOdc3O4R0HgvcoP8EhE/HsAWUpdgljLew17J+fD2+0YgD5F+wRVSiHyvdEzT7aqA
zUhgGTg1zGLRPWv4eQnIzxNPeYMT8qv29rmWyn3KN7SZr51CZt+1CrL4h1hI0JsWnc60aCdLV4XN
YlDnr+bPhXMIbi6IyEckvZuxngeGb2RHW2FGSOkqr704ktswbabZTadFVeF2nACvhrAWshPeR6Lv
BGtFiRmej/lhd450Wlbs4HM/DdMp0YjHxJ+66g/xtWHP1WdTPmYPm+wQlJ4q81iel9orJAfG5dN2
Eu/rykEbBlDAtNHM1TFFq99v0bTTy/o/oDslV0sWqO1DnhhKZkeIJ7KRr3ZE6OnMaSRalzFcrbD+
kQwblBfflY5HKr7IdUnF45u8qjSEEEx3Q1qLdEcVlRtfRxYzI9+zMs0Hh7NgED0XlKxCRrRI1Ahf
Hg4xrKueN7RSWRd65GVTtR6TQU03YazWyW8ENGwmBKxgzs8o7aDrzl6tBFRQCwNC3orURGhHMqfJ
rINMKRMbtYBPHOailYRdpDx4Mea/p98h1E3MPJMqQXKNv/uRC1ocFATh+GhmRvP3o3gcPrxDOtQE
6D2TuCg02lOV1SxQK7v4yXBpsMW+UJPdwhw8OX76zFhXHoKBhDgNSzv9TwhV6AfAdBYaBJtftL7R
C6PLr3C/sr8DFETBy9w5h5MszDzZd5bdBgR6USN0FLQ9+iiM9Ew53vdGU6ZurFFQT1WuoW0XA3TC
Ktuw1psB/e4X3i6YL57Wb4YpFzCcFDGd0aqj6OhLfmjiz1KQKQ3lQeFoyBZm7I7CQtjmrG/Rtn2z
z01Ln1Z9eDpI+TqwM6bIIqpOfGXG0J5BOZLDPqFLShQA+183Kxhi4bKeCDNHOAtxVZUqJssV9xnj
sg+RVHnFoOgy0ZavCLY+qqChUkvke4juNPS8p2cYMQqwkLIirC5kzDtfR86gXc6wEMNhOfe6c3AO
sA62rZisNJXm1Cl2WNMXyZwDVHoSKKRTZDd0UHF4jWZixnQbUyPw6TD5w0JhteS5g0ZS4iE2sbll
ab/1FNBef6JkbfOcCGEi6K00VGWbKLg+yQv9my+PWhDB7FyDUYPThCM+lSTeTF8mh1Wbz8+8sFtj
cMlcI/CUR9g25FiI7l829D85a4pSjXJXRY5Mj2zXPA8Rg5kYlqzOr/ROY6PwQlaHtehvH4t4Ibtk
H5MzjqbBWpR44t0EsB1/94+LOl7AJCUlbJSsoEFIFV54PlXFfDYoS4o/CTF43pFYmaxs1l9X5bph
MNDTHBI6aFpU6m6Jfgq3CJi0M0U1hZ7EhChhd0yd9q26R79mmC1n/LXp1TNemSCnLXGebFfQukdg
HNaHj2NS3kilVTjrcV5tLloWZCHG9ku9fS0cSPAHGRQ40/P+4oeu2bJ6xIMTd1tK+1YJd+Zrn+c4
PG34HIeuSleglwphZKMKfyQGN8AGgp+GN/nmajUA/8aUCUYbbNGAuEu77YSqWBXOPd/Qdf1e77fi
C+XBGHs3hhgiCOlGX7xWfbHC/xe9BcnJWEE0SK9Z19+EKwvxIgiT7uUJrwf4qVlyuQYlyfH2AKX1
MIJymeWUKEKiGjLIC892kalHaPmPjsNUrtOWfyfy9A2c5KGmtkqVmh22h8mkEzRWTv9odWiKXKOv
gt4nLGh6HqFF/WHu6T/VRUu1WGwvkiOFdpW8epFIjgBAdTAUi2Haxk5z2jaoDE85V5K13UKwU+bU
7Wb6Ax8Uj/i+iOQqn60U8NxfLJjp6F5bC+YmyxF4V9qmG3qfLU4OsEIquybJPqvr7bDyDn1D4qIX
cGSrat93FRbV1chdl7HLE69t97engznEAJpQDxZmPBVzqa2o5iEFiYdouT+2GTv0MfII1GE4aOZ1
oPlR/q4tqqovRfWvtzwsgTuG+Bxu6A+k08LideFzstC8IlyDG/4dVykYowWzYghyQx+SZxSC5CQ+
r9IGYHkuBJG2ZX4rxoFrgjfeIpQr1HioiaQh51hjpT8uIZp0eMKUDJcMTCqZwQOoItU209ZY17S5
V2pdGj+3LB/wmVvbpw96+4NtAgbuJkOH6+RwZ16reFr3xgeNFWrnxWTcrrP6tQEiFx52kYgPIzjt
Z/tmvysHVw6GZ6r71au8OLrBuu5ILe6QZMeU57BIcCVjHfUNLItWEkTpwcnnX8sdUMXhrI1wBdeo
Ehbr8q+5d5H//hgIylST/HQnBpuOuy6m4OcRWdC4CLP9uRFUF2l82rbxBJWSUFK8XQoBI/c713K6
n82484D9wPo0MlmmEQenVcDQY9B13bzmoz0l2QdeSZzay9d/ckwG0KyOx7pUkV6E5TFvTyIaqvT1
KnodBlctfnkWxewHWWZm4ZqqAJQMU6rYm9bCaCce/8ztNrSW2vYbyW1cu4WduVFxdmIC1WZ7wdTM
/0tqZVLdiRpeDGMiRDrqqUTn+dLrZqVbC5VE2w6Y7EW/Wd2q3wZ/rxbfGdy0FAixN8JBGropu/5o
XRzGU44DY0WDAxJ1KCpZyb5WRZVdlCDuwvD9ploewY1ddRQcEjSBoOkTnCrjE182EzqrRk8iR+IB
82hOxVvfLZuU2BxgALgj1+Ly7LGopEJTBnieERhCgXF4jG7AHgzAPdws43dMExfnafe527Nz0+UX
h43imvoHhyiB+Xgr6+V2gFZypUHwRVbLLLGMiq9pi05xs7Mhwt39d0MXipYLu0f2VmUHYsEI0rJ1
acQpcGJSAEcTYtFyB2f4NyLBG0uS3ycNFTwW/Z2eJjXBRbkxJqvrXFkALBOb7EZJOadMCYjk3FyB
UwmK4Q1OHlLVfg4SvCHMuN3T1ZfL0NxKIo14j6Wl6wCF0z/FGG+y9EHQ0MJ47J7WM8zEZp94Uy9m
2N17U+1HoAWBY+B+OxNLQ39uoZm8aHG9R/vuCZmi19gXxiUi41df5Beoxq+m43l8DN4miuTXVPPT
6YIO3NMkPZYZ3j5wJCAquQXElkoSLZPdPRliW8peg7fB42xw5Jgot53di62jgZ3PlcZ1h3grtVEO
GL6QWrzJyWqqcV9PchXYPk/X5i0PnPHtkIcecMIBw8SqyQR8oWOBkwww7uv6u2EbBzkwqLymx/1Y
eccbVV2CqxCN9kFN0UsVm5xdfSsQhEsAF6dP0flE7zXepojAla+TVpU6UGS/BIrMGlcyK4DMhFMI
FgI+beKud4BQK+m3XVtYqrxD+jcrnDvYmt9ow8xBGxHqUqCLidUOyolnm3Ug5BD/r3ZSD2x6VImR
UVZk0KjHybGIWxNkhBMPmRpDf+yNBx/g+NOowiqaJuViFNEu0F8V4Ml3TTlmrAod6fhQ+zdqUD+t
2HF1xw2orsM69+NUl6WuNTIWTewlPAT6xmOWeXsUA7PnkwkpTfuUf9PTgjJ0Ehttfj1R2yjPY0GG
81a9Hr9ui9YNAxf/5ob3i7i6stXvu4sPWCF0pEgJNH5KI9w8Lnx99dmgAPsEB4KHi8G43k+u5QM9
yhhgEg1yNTxD+xI2FslgDinyUM2rM20OD8z8RJMQnVp2JDnObv88n/KHjQpY2/M7yw+aqze2wrqK
nb9q6ECfx2Plfvdcb6opYM5K/slaHkxROWw2yGKsemQwSq2RVGh8aFnBCJzHmv0rGpYEwDFzZE5d
QLH8YQyYC1jzzhAddVwiGOjrm7ZkPhAzMLHodP1XtDs6RN939fnpeFjyXSGGQoTd5R/EtlY2iXQQ
xwq6keheGt35ek5DzZVEh/mF5ZuIJNFenuYCHOcak3BwBOQDxjNbO8/zaLOEcXRLe/GspVNn7ApY
vPJZleQtqqwdpDKUgyjWWhbQoIUB8QTEtRc6TqdiEswdCxFdlTeJoMD8+XuUckG5CoOgmhTpyClO
q5AiFB85qW3S5QZL+eZ+q1EEk9ryC/yxjoBadkoSJ66sbZQoL7ZAT9AGin1YmVcvTuGlw4sFHT3Q
n5/7nBsZ/LFW/zqJ7aq4m/ZICRaGZJqUjP5bDdIzMwm8IwAjD9GssJSAVl0/nlJRr21t0+V3vWeS
VpsPJ+lNpnd8xwk0E4EruR+G/pVQZ9br4I2Mt3BkSXUkanhKoXESlhNw6MjbHH0SHnVh3J1SThmR
KkDdtbKJK9gw9rfAz83i4PWiBTj/RtyBvYwM5B8FX57xkGS7dmu7ByllkactjDyQCvKyrCJGGwLu
IzF10aWjDOrR/h7I9yOcOCVwNKtu+y/XX3mo8f7Q1Q6geW4DnllNO+q+ajil8c5ZK5yEVj1ewwar
aZIXZWsN78gKGHvE2FjTyjZuRAuaZNdRdTZJB91V6O6YZN/wlw7n0FPxfyT+z+hd1fPKYJggaanK
Hds1L//JlvzjzXt+gcq87p7XexIWhdlxC8+Gdnk5G3yeQjNhI3bVdDmOyvtM7lynxOMLqfC1x7v6
3xJz12RQOEj/LIcc3Aa9tnld7itKYB3JctdcVydpVCmZG1ys8nfBfAGWrEgNF6aJvIJuxfaATwkp
9bVc9nNnZn8WIp2e0nTkBeOkCccL/sMpGgHE+g/7yAluTY03/1VUN//5bXSepzEzFP6kFePqVbi8
CrxTizQoVde6FWuK8oEKp2Di2CBPIlMYM8C+GMqaaTkoj5Gs9gWDr0axRyci4+X/DuOwHxpTkHdx
8ymb6ljvA55XUJWghomb+0v4GjGCKYbXxs7g93MNx5c5WZ92FnWr3yowTj3WQj5+SJWDqu/6b4yV
I1HUkP3Gb+I2BA86vCXMeTn/+R4CcMmMJ8oxkYV1mFOEtrKxSKe8bFiTbrPKPPMm3XRH2sqxACb2
xq0pypbs/ZJ1zjBPIOC4Fw8z/VLKEDcso9KcAIsrAZYSoHMDMjF6O16PzU5qzYor4zY8iMOgayYP
5vtBPHi6xZqI/OfSWdiKyDz+dlZsIMFOfDgQC851XJDMPGxWhnFd64kQjLfmzCFxrffpfahlCGdy
//zb2WUwqzNGjB/tjUV0czvwnniP/6DCWTS9FlFru86HRv+WgUHntoz9AkPxUOFzMsIbICZ8VGpk
iqW4lGhZWQD/h0togCS1BszbynC3NVtslYAlKiaVCYzvLx5A/51/jAJ3+Io54khyzCnvWTlaTwN3
Xb7oU8K17H09RxlaJoTKAV1kwu/S8goVqwldMrVKMQqA1mfnv8aeRJWkk3LFE9Wf1XbVg1xBR5y4
mI8Ql6F+WPd9bVxo9t3af8iGanXLfSl/tJ19EZ5knuO6I4r+WGLqMfwzAvnxBizbTTGtbQpQD18X
JZ1J4npufbs9s2iGU5pFqhLyOt5IGcsaInt2NAU3b3wVHRQaxq5Tvr5ILL65wI3UQ6rrCj00DUjX
6xvAEi1vQM2GE/J+CdOyqUQahkSUWP0Jl4pgX6B403J5tdqvTHrPANTLgm+xvEpmN2zdOoPnA83Y
J2pdb7hc6ZO1qjpw37PnkpjvTIJpGx2YppwhvBe2fCkfgYgi24MyCxhz9ajhRNyPRWXXHxbxGuVE
W+TnJXPraz02JbArPoA53TsFIc1PGY5xGybV5fegapzFWvRR9S4z1KxJy0C4HnHlEMbqPts91YkS
vdOxOdpMjibQB1JxweBz+RmgRVbBpw1Nxo8PMLWFpifx1LIpSpOMT7tq0fLejmsjju3qA+Vx9rX+
ZRBfr3eE8O1wzPLWe2ZpW5r3R45EVfJoCaqVBt938OQLuF3KsQ04EnFMNrP9Mk/GG6StLAJKYoXG
PYgb/4fbTL4qEj2eS004UDUC2q4XvfhT7WBGndWjHKuigkfVDy2uvYmygEn+6vV7lxZWg7YhKEDs
wEvkLGf7DKWWkQWWjiViNTEKd2dGGp2rilWDuG239Pof4cy+OeMY6RgkuPFgBEjEy5AnpcFll9eS
4XtX7FYNWEvUUXZPH9nXJjq3Aoxac0siNIuulPw3fjhlmws6Oge89xQLntAduU5V/jQBuTvZS4wT
+thn6qednjACf0JlRdhIcW9tQHpVVpo9JZzwZ8xJNQk9Sd5wlTuuF09IKlCtoOPxYWvWcfnHN2wA
tyPuZW2N9rKQg3KNqk/Ux3RRWU9tE+KoBeLXSHgQQotkookAFEEaBqm1w7BOqxGze6DOgl3Vlyo7
omACV7rcWYDxvN6oGU5mi2/14IZZjmruKCKQMPOAog785OFr8ObPvL7EO9yphpW4A8E2B4veuSAM
hahK61mCSUkgkcJO3fWJ233PnUV9nvxqb6d4HTNAPNXEwI4qS+LZJMRRIy2DI1kQ7p1HO1sfiwbF
j6He10Xo4uWKj81KQaUkTzuLqn39n8geD2dp4Nk09FK8zJHIwS4YshB5LUrz5b/97pEKFb7YkRkd
Ry5pRPMsMlNwE5jN8gJB70w/SruKJsh+K64nVDQy9ImOQKnBJ1X3Qgqdm1r1gMDdJAYNu7znJNY+
GfXCqvwCOn3Lr1SAdbeBJ0moTbPdjrKrdGhbztlxzQBDAkuLzOWMKn1cBEft9CMH7YYUAC/i6Pmg
fTwSG2+aNlJKAmleWuxvrEpl2ec8TJzLRfckZEWqzWDjeR3ZayWsm2RYl6shcOokqotQudBjZWNv
KHc3qnOLEn6RFoDXxZnkzzxHE1O1dnOJ23d8SlH32FkXXWiaAp366v1TifRpkz8vWLVXM4NfjMzy
iAHTyy3dE+03R1F59J4XpXXTcuI+aCb/0KViH+Ws/04S74hWuF4wtexpGhHWXZg/xTPUuxcr1IIi
LiBvIGtpaJ07V42WtWlm5d8kgSitzqcE/M2jpYpehdej6QXLlh4J5bgYReGgvS/Y3Y1WLCkORepA
dYGEgnJfK3cWpHk4trA4IethDcePnRtVKy4vsDjfbxC928qSQ0IXDWY7YLYgBxlelRYVCfgCgTJ7
B4vIuXXHAvHC4dh9D1JVrFjvSMWupHuDew0BSHbJs+g7jkMsTBtPgUm77qSVIqXR9MynvA/K3SIb
QG9mGTs3GfvrmYv8GwPIV6h7pedacBFxMkEaH8lWPHAyTsoCRIQOvPBSkVWP6buqgoRfGLdkEQrP
vpt+t81KlMcjTIt7O8sMmfzEa0CXJKa8FxhGfgVPC/i/2/g+hV/jbl/iO3ezhbF24OCVgt1fPMNv
Q1OryCMv5WdLLjb9y5EGAxIfl4ld0DKdZrWEhXLKpb4pEiF8NAoqJ4AEzKn42iW9TVrdeC7Ub+En
TO3CDNz+Nms+Qzm/B1Frfd9syMXT7lwg+VIp9UN0UPM9UClNqRNO00hei/7W6PAXdCUltI014lGr
6XZkEkMKmVDGkXIgNVGqi6KklxmvzGf7d5L/onob2TJr+xnBqAQ8DXeA1WdD6V54A+LvN0fmHfmZ
1VEAr+MJDIrz1EiYWZbUTIjC4M8hWDt8Zj0E15C0d+A/ErQtjg4wMCRubmZRCMHoj2TpPm7niTF3
52KYNnWNeTvTChgOd3HkhmkpXhQsmvi2neDqHPiMsJURY6KQxVtO4CFoe/ErwL5H+7+V2argbFnA
Tk2LBZvNYjMSFvBGFy6dw9hx4ju8sKeS0ymTUXlbX89oEeeUOSr3eTYUt/zOzgDv8TCnyH4qNyl1
G3TLU3nIQPo+A3njS2HcLvFG/KIw/4sxLWknY0Rh6MkeLuXR3/uzbiE0g9oTKM6aEJpmJMlgVreu
euk3OSFpzV5SNYzA9nqDr1ZxSWJ1xcX0jxftP9f1PDeARck0YMPax0/7Mzr3xPme8iLx+Irw8B4q
JhHyqr4H/sxM+jVrt5sfHqWJDz2ooz5SmMT/txk0GAiyLi19Uot0M/JOVzVkU2kEMmHK++gyqZhw
dOuzX8XM7QKXdU5A3JwzBWhx05ZWPtJ7MzE+iaXoBv9mhpHilEcZgSSs4pn8Qd80m3ugzORgD31q
l9QUToPkTvntH6bh0swgllYZoWWSnX97/aTLlVEb9A2CIBM4rQ4rK6O2JmIvMfJfza/360UltWr9
HtbWmXOOkq2QqRZ0HyXsRGwQOWLtM43CDRP5odzwsMZhGqYBvrg3ATSKGdAbxI3ZQ/xTJsCstj2K
5So7z9ez/g4KdEQD87V1YRsZercZC0D3nSfCWt+4HW/oF7LMJ+0Zwqz+Oebtg9Bd8uEf2iPZov48
mwyH4kaUBwXUJhDdB/1cKXW4pj5Kk8ZMRfWsd0vwVGdAKr8PXxmz+eZmiWWrTCgxKCURXEHW6gfU
SCd8gpurZVOmOvSD5asgpprbSphZHVqv9mzUCsoYZ6CPchEDq7c8v1NlFuTFfdhEA59LGgR/r8rM
6XddFhbxjRmqTTZGaaMJmGsbKjtT/tD8sd5wfKpKFe9pzMgmwtlU+ILPqRsXGcOhran3MCjkRxp+
/QNBoPVQbFHAzd7USz8L3l3G44PVgjiVVFMW32Br9UxnidXHNIcpiOtZkytEudHzlcEYF8sNw/mG
STZL0s0SKUtYKvu44nDpfHUrS409hbg92fLECqQccdvv3qmyZrJoxr/D46OrHVZg1XHNP1htD4Op
r6FY2g+KRTE2lA0+5JT2avS+7mnq+cazVbrhE83dqXa67sn27TQWpjvUnUw6ZxC7/+j4qEPw4es2
EwXmbrey6MKjXQElhgQfj2xjnZZtVIf1YKgrpk9Csv3NgKgCbYSnHmC9W5GlYdwE9Xx+HdMKwthj
eZ4/lrq7els7kFyfBocOWeenAtiJcWk7mivEneex9aM8i8G3b7PyMv9HXGQNZUFv4mST31tRehsP
HxZsuDx7nTuEMnZzv85EjEu8tn6sD0jbewcmsQ6Oj09VynhyrTsvBUwVDsjabJSxIFxCTfvd6Zq5
Qmxw2Xw38lSFdtiqVVMzCwvp9sAv8Al+joT8En+8iMsAzlJSQCaLTqm9Lg62zO662Pv2T+7M33qP
nNZQUUc4kxawkcxfYHmRdiQ9moMQBNy6icqvWNyaN8KeUKjA0/avOctuclwLGF2qdq+E4cJXCyNk
GP6KR+plzt8cYGtE6FRuU2+x9JgEpX1PhUuL4858f7ClozERHwNjtdTT9j/MS1u7QNIUEVt7TARx
h3C4tHhyY7tpVobz8AiI+G7+m5tNUbAKTJQ4C8a76lB+mHeI0bngv1WlI4t9Uexcdx+g9hSMqwf1
cx5JnPCr35Er1iqj4PbwZ2QKgLXPeDVWbUujfiCqM10OY5hJ8Qx4ScvS/EIpW1RtZ/ZyKwPUtvPF
pBpvvNA3cjmxvwBHhlqyvWmgtnuuasQroYSDLNQhgEjCxbzRTg2OUaLfB4ztoGSMyJMf+p9gfozq
e7xzQqp1yBccLuqLDlgcPTyfQcb/w4dCrj9L5Qk3xAeB2YdYcCB7m20zPm4IuvFLWZnznR0ubc3P
k8K5hGuKmXyWefbQ4eDKUdFIujukK2sE2o6m371SzDZSyKpelsYBr+eipI/apOS/FxY7/ikdhK/n
4R2axrb8tnocZHmGExlJbgQPLEoz5BYZA6ctdKU9bG7kqFETAdiddOqUCr8QhPlc2k+VdNMcu3+t
gZtTynEEOrUeVYXhCXFGpAinUrredGrnhttQC5EF1YezhCpVBU65HzCBBOtJJJkAbK+GsikAoXqf
13QgXgYOXcb1PeU4IfsA56blr7DCF3Bii+VGtSh5tEebOXgUaN0DCWZtiK4PuPC2YvAASNbVtO+k
Kj9Si37YkqsO5z87Bl1oHTbp5c5UMyYUMAffUkEgqGcS6ZhcxzRMMpWQ0rUF4HumfD3WLY1MSrca
r56RrS3X5j6Aq7pKNLfsMxOHJhMw5RkwqOcylDbICmewqnu++Atmc6ERnmT1AHh5x/q2tPE1F3AE
Ez08ytLxti+Toz/cDdTN7VTQGf40yODf9d+6kk6ydIallMsG3hj9tm30Pw43ljqDcVd0m5RXkReq
TYbPz8n1Q0ebShU4tNQtI5sOL913A3A2MFRtRHiToKeEL2l6eblDjSrnBAXE0pwrcQdMhXF9Ktha
grgB1XsAt+E+75LyeFca3QOXAgvQ26kfrlTyUOnewwr54TP8ZJPN433Q3cJRGWScVzB+mSCI/Mv9
8BiPSlIA5r4TaIo5UX4HARoFIRxWWwYeKbJZ7S0AgKakRiDmMK9a83/QBt5l91bMPJ2URbLiBZIB
YqXj1U6157gEsyvvIalF/ts6X2s6ZLvwS5Gg+d9Pik3g4gEFNVylrQ8aNoIkLxTrr8/F5vjIIdZG
A+4EKp/ocZgdndMxmSRt3gdEjrczChjXH4jBNgRw6dHUqxsl1TjfV2sZgd+Fr+mpKK3kNVi+Oin6
LiNDtm84VWk2aJAGSqRoE9MAj9JtV3xh/K9dXmKkabGJ4eM0uy4hvG7KnNF9x0Kh4EhQ7RxtLXMy
bHm9GcX2s2lVEF7SfvnJG7A2RuThNVZCVi1FpvOhxsvA8itu00xxNvJQACaWn11IxQ+tjYITnfjL
cxE3bUJDloOqvBhs//ZBRRlyZ3o9XRI3d18A8/iwGS6QJK21p719qk2N0s20dGi6QZWR7yFAEKHv
hSEw2pPeyyg9HOsdafmCYlkI5HG7ydb/8QIDeeivH86S9/bDoOUWYyHFKcqNzR1fakD8EeqjEimZ
BaU6p89I+7anj7HjvJ19f6XWIEmV0876hLDlfriSnNz6DMSe/MtRlgnbnFS1L6dglABPVcqMhGve
W47ny7btnRpect7VO1BH01QKgKV0N6c6lzuVCf7d/veqRn5EolfHCWylFf7MqM5sRwk1hnTM+1Ut
erT7byXqawK4sZXMIwa1NEoFFM92gYkB243If+O1PlruovQjRRnqQL1bMxEEf4ciQAbTyFBVLf1o
ZNeUI2Deif7pGo/8IIRcK4byM0DAil3RjGPKR5ut0+lXW82V169u9e2uCzoHy+eWPUKB9fDmwYxk
yv4mUuJiaDhVCvqaRp+Cfu5JC3miHMXa1PIXr8bxq9qDV2jqG1C560G56kZ3FkCUKt5nCs/1T/OS
lTIyroluhzPRAhOeL0cxRGgfw0e2BKC+4/hhOb9qVhRhieyAHhCPepLjJWvQoOmZ+33pEdo6WNTJ
+BxwE1oXLMtTJ3pqMw6k9Adhqm0oWZUpjK1aeD8n/vECWQEOErcrqy+SS8Unpe3uXwYKBQwBRou8
xMlkuxKatNUTpG4L5M9U+lh5Zcrg6yMJbISS6URvGVxMDHAQQnLCOoWMxcarhw+iWO/YxEs/50Mm
/bgwd1vV3xNC8mSbF+iMrnGl47F7Iwogr0fY3YWj1Bwn0RlfmENGUxSKd/wj1OcCgYakpn8m2nVD
m3sYCc8H+UB1QgNbTSplzPMxwGRN4uzeqinFxmakaj+tthIe3dOX64HrGAX+7VV0x3JMnMQikihA
nw+6vYA/d/sviIrRoxsxQ5xNKf8QaQMybNELh0IYdW5gXiugrHctThFlkqNj7JE6fl4GMCF2c8L9
IsYEKeVMRLeHy6nd2ElD9qu0gP0wJhqXEo4ONClvQmaAu/mjfe09AJ7dSkE3W5FXctkVJEKuVW5W
1cpH2Dq0opScSEoK4qJg2cCXBjedhNqfHvA8JZV+fUSq+G07DGX6TFLxhcpWunXRm+R7mAsvgumS
Ov+BkvRI9l/gBqIadcqxNcWDL+5+dlASikr4pGwX2fCA1lwEpsSo5Dnep+kzlDjx4eiwV/2Lym71
VpBHX0cZOSiy4OHTdhuvm4v0HE4Xd6aRSRzo8AmZW8F1wyXxaVRixs9jR8TzrzlQjZO65YW0APQb
ubEGQwKtHX58q8x1B2lUgDK1FOjS/TLPH9EP5uuHsy1FIs4QJIX684N0HgiSJ9CUx30neKAXYR58
aNqE8CAxQo/CBESb+wQHqWXtPyTROsssdKfwyDn+ozoszGH/GVIoReFP0pWmdk1FKG6k3gKfbRpr
YWhfjI6I6MbYC2oM4Hr8/zd7dH5J2yYkD5a//ErSc0OMfjd5Yr3I47xPl5SevK9f2NxgGlGXyK73
ogfzk3ZFejTzTuGFrWYzwuTv67Lvow0LuOA/hRZn/NusHOfRK4oOLrp9uDOfNncCVo7VtSx6EZ+G
Q/gOTTd3odenRqT5+Tf5APEN84v2eKvqPktk5Ofvc0atiUsq5t+ZD0eDECpcgpfWUVG9UZ2ksdMQ
wsqS0RismRjIU7dPCPK87ec8VL4SkWY6FB6r8G5+3XBqmFIP+BtSE9kD5hurAiR/G7CMSrtjiRMx
jwRlPZNQQEPASqFyUExekVA7il7o8tVOxm1P18sWEi1tmXsKR9Sa2/mG53HBOTzmb1RcXKFEdafv
NwFqBOls/8ZnFrQ26Fd8P5QkwLHLxXgBIYkdsELX3pQD+czZ7niRyqdP6pzsgQ8ghQyW5Z+cNmOh
XGUhlLfl2slHCRzrR/P1a3VDc1RSQJiuZxfdaPs4HgKABRMNYVinytcWYCWIihA8TRRA9DTLmCre
B34zJO/zBdsiMMEPUVxSSrF97dHiws80yDePX31Ptotksxv+4wZTQmBBR7PTq5WbhgCZ/yk7taY+
Z7Ahf4wSpn+MalFd+SRf0wXGbC/hzn5uM5Y9SJTIPnAydLWNkP5k4VShrMaPMPmN19zt9YtdP6Ej
FgYi7y5r1MeRSsH1rWAVI0YRnaODkgT/6XD9K9Y53UKkesy+nSKDaykWoeSTj3lj/wu4KtGgE/jc
m9lVAXPPjpixLAum/rd2BZeUGHhRP6NydEOWEWmY+QmIZjKX5IIoV7DiHXQAL+IrmV5WMjJSOi+m
XfcPNV/4Ich/hcPqbMNshurcpVvHjIZXm7gdRS0ze5VVAt4SBTL9gAxGPqLMC1/rpPClU5Ozad3P
lnzQxaxkFOpKb2d4w9pnswX2496SOjs+vWWsk/PApPKGsKJHoMnyGqp7i5xX7YUGoHMpxED1AuFT
pxnNu/zzphBxpnC9giOXfl9hcmJeEAJCQu2B46qd8fziu8V7QUk90aJaEqG5Tt8lLsBJ84Y81UlV
gpr2dk9ZPkRLR8EpzdLZPpErD8URta0Fb44QvsiLRuNDRBF1gcyd5kliE4uvgBjTMexj6wDukVAS
P7epiTicXIp1HHTWYxy6EEM3PObMXTwmtN/g+/hZvr1miYLi4Ag2lgv5XmkFTwFQzSa6DTPPzsu7
njn+dDLvtx1+Lq7sJTOKxJogu3CIdjXoVdUbfVx9OvwYfTlarNAY1KaoA1h+/wlDG22pI+sbgkss
aEezXv2y7gZaT6AS6/ejfoYHlDSrd/xKJNF3m0kdJDug753PZmhOIfZ7B7Cm0qPPEgnu5qZ7AzDV
znM7jzQRKWtqsy7KeIBWpgxGvcASwvWNuAF7gvwviRpaCVBfiEvF1DDjDg2WYdFLCQz/GPMss0QV
IWbSLrY4ZURcotHkgiCa2doLm/4ncUegoFzbM31td6FtpzUksLrKTzD/r01ue+d/p7sEGV837kPn
qve3zTcoKif8bW7/WnMeLEDiOwCuqEWJ7O558LYpqPlqHDZy01UoBZKDvFkGztoFcaTXrR/NV7mu
6gc2zZ4CGv8sLtjsRHWeH5dH+5Jf0FL6voqtbBjDsqxNlMc6YY1+6OshCar86NuOhVsdl5k8nGp7
9wkf7q4tv1TzpJkD0mxX0N3s0KvulbiShflnaaAggNPTlZQBX4hdfqZo50BfFLBejEyiN+XMzhmJ
QUVBlMuoB+myyg6mp0O9CvdhZZ8rGoimICtKH0kbU50XP9MYGmco9T6Ub/T/r53Zi4HETw5h+YUj
nAKlcOhyjtJwc/EV1ZHiQSJJ2O2gvaaYnCm8tZoqiFiFj7j3k0SZgMFdjjkDTW7ZRUjmhgF/U6FR
ctm1X5v5bmcUpx8MM9isfKphIJ3GsZBelCGs+GlbqYiwMlm5EIdj8KaG3LZUSB6J8tGXKh/f+xNJ
giZFyBfReJeO8hofODimq+/As9HASzEar2pAQWiUE48hxLBrxfzsERY1j13S5o2TfjtGCUzfUyDW
zGc08OPcEFx8UdAPPfnq6JiqNSG3Awh2/KGE++QImmrfAr9ANoOsm6jjc8O6TF4wXBhZC4i6TQYF
ZslyrUEb9NK2ZMJBnW2S/c0JQMnKsfG56uyjkadNJPUY0XCZagqM8mRyTOOhNt1p4cvmrZHtpn7w
kUh+Pyn8jP+buE15RpKk7533qI0eA5Hqx/a8zRj0aBb2t5aqhdk/7rIuKQBP7nxKLM9tC7oGUqTu
5/IQjp9H9ciUYvX4SpqFwpvcvoejmb6gXpPSRnQlTdLbQyr+nayoBnQHmMI8n+QwBgRGH9xQj2A/
r6DHC8oVDdO/MPhbCp3AvTMI2XskqfZB1AkG0alonhC5vt+f5qJUWwqks4BnPgKQtmOPOYpvvWUQ
Oc+WSSLsVlmrr0voM/PJ0eCMUHhA3e44HYnixWNO2QZI+QiaoRQgHG2/1JNIjnPljaphzrrmmbXU
VpKv9/FGPvPGLiu0VpRleHGBzvLy4tQfpRKQ2tkM6MY7L8lM5piLsm+ZNmGCfpHa8iXr4OjBhv8n
n9NxdzGvZi77adXu4oXDd0ZKbPUiDCGW/5vLQ8976RmQgK74BO+Ew4PG1n8vViModw1XDOSyKByc
Y2XFcHxOPNV0+2SpGg+OnWorqtwFDUf4KyeGam2Wb4mQdaoTZnkAvUnB/vD0vb88vuIv+2jYc8Zo
RjdzR06Ro/C8UFwAE1dQsaBWtZpyXrskctsyNPtZxTZt13tSuDdxpdWjBaVEKoWFRypNEbmVR/sd
gPod31o2Ke7LVh/XA5bM+zI9+dNI58PWsRJ6e9tqZ8Sz1Y+QuCNeuG/b2J4UK1TWCDIbKVyl1c2m
Hc7/jubClfADI7v0ipNBcdBr49EGUCF/OzFeunMDDy+t31OaUe7CCc/NKKZvMoUuCNLDVWcH5z7R
3h2jRHqv0eCOVu45HhkdxZ/vbDJxbDT19FuS9fSZshelFPHR2Fsvpy1fAujaaF9jV6u6IUTktmVT
8e5bvtHwxsOFAopvalIHzphoXyrp+NGeIx2TaopegK6jRjsJ+Ujn+djnCEoXiIpOjW+9nVCVDij8
+PmFD4px7I8aSOgSsnY1DLxj6cSFfCn/hLFA+P3iOlnoHhfvGL0JFF0KXozZkGTLRtxabPAu6wWu
7ffhZDI2HpYjcgA2oFWkpm8sX7HU6JFO31rYVtiLjaUueWGO2NXzYRiJdxXYyJ6YgGgFv1Ol4tR/
CHg2cvQ1ubab6+P/M0RpNtjnVZlLpv/Tj5OoG9Cybr1wj2wiHkLnDRQrMvY1dn0yUX3uJDUIB6uT
gaArHX0OY48l9viGfzXt1JX3DzRplrnp+8izLCe2jBQlNsyTdZYvbvi7eIEoo0rlD4RAfOQXiHv8
7fXBvrtYrPsqAmsYUR8SJCUfOMoA0opR39ptJaYp3zTH2geOivawxiGSVJ1npV+6oQLAL/DQJ7C1
HVRjLypCRAyMIfeow+YzuMVsr45OHTP1N5a+De2lvX51j9obdPrV2pOiYZo+4WcmEDfjHaNc2GjP
c8twKSZDsWTPNlhah9Fyw+antYv9JR8VocDrN97caKEHOb7n+6Aj+ffoDwphfBGwMTd1OXn+WLr6
FNn+s3olFaXA7sZNx0MILXPiiJGd7e1d2s/fntLlNVusd+33OQxNIcjAOXzo02p4G1VWA79t0feE
VXEZ1HoI7EA/1kTYj9lbOmNx5G8xVifv2njdaN7XGRLeOnQmMaVKDs2fX+K1OExWBNkxfbJ+9YoJ
jzhIWsoVDq+PFkdeVN9xtgrM8vqG1x/rk0ly4dQhHtbv6gqEp1MYAdbkLb4yf/mokN625rWaaMyy
uXizSmJErJsZuRGkuBdPHkaxYvJnl6OBbsMC1iLbHIKZhpzFEfLRWlKMu32XsSmJibcVd8ZbjmKT
hZ+z0vrEKQ4AsHWQ1s++0/1hxRAborX06KSdKoK8hzrhp+43RoJ5HInFCbpyEZtUD9+XKV77TAET
/ylcK4p5/xZgaKDRMv6r3sjspCRP3vc93c4ukxqOIZbZWqX0wuRipe6Jtye87J1QQuaR1GluIuhG
a5ikzpDKHw6AJ0f+4hi2zVm/UtZTMKTjTRjqwg9LcPVsYzEGvShWh0o4a8tvS8om3xi0vNBgUEIy
HlDukaGPBjv9KiamS4bPCihsG8UlCVLxgDRh9g6dGe8CdeSk231bwX6/iUVFpi4m0L0Eh+jSo518
XLGzlj1Db5znh/wJIu3UGCsjXCR0/O23l38WJAP12zyG+mSf7CoNrGU1SwFyTKUg/m/S+S+t8/Q/
7AtLPaqv/E1Q9x699qJojhXZPklFExcHAW+ZdcUYP7HQWpS8DGhX5lMXmHZ1wIir1llmMkhczI+G
dkYRf7yjyrPUay3tPep4ypbVMEV/1wxNsE8n1BL1KcmLK7rKjOyYuVdHvVyc/gRZwaW883IPz+cR
HvRBxDvyUpNiaf/5EkfjIEeiFTjaZa+sHMTEuNfYPNNKmLYT5VfO6iLmpJv7iJ4tiScYV7einphD
W9ZmRXQ/ndE5Z5M9lochSOWB0pcIR+aBEBOOnLniFNEXjjshJr0Qk5Iex4xZt+eka02i9KeH4UIo
K9rsz67cShKNYMmAyB3eZLg7eiWr6dbmFdYuQhHi3WympUkA6cVzW+01kxzdeXLP6z1IOpdv6TAm
lviLli2DDyT6StqMcpRdscxZXuhkF/8tNrBEKO4o0/pfGo2Ib2iZb31yDJCNBzCe044iYYaKnLnh
jy1Xs9J62mrWelVVLJN9VjRDA6t2bLbWKiFz38NtlvaxuOrWE6N9vEuTneXSYuytnS69KUh5JMIl
7j+uV4yvXks+AkDdqEZnf6xUNocxDdE8X287Hw2UT1kh8BAn+vvBMKdt7A26swn8g4Tvn5Ddag35
v+UaYA+xcWb7f3+3bPj5bLpBwh1nO4toBSnPBgpyNX2nandkB76n0oNWWfpZJTbr+io9XiIQn9Kp
cNvzFV5P5q1ruiaXZKg8FqZVWltbQVDsJZfBPnyx0SDI+/1hSve21J6JyovlbvLDTsltQ5vmINrB
Dj3qrZlfm0cNHkj82tFtUhSAViOVMLHfPibcWCJtnjqgkVZpbRINeYwRt1BureiyFQ/ndCPwXXR2
vbd2dWVOVi0puCbSU0ylW9HzIw4GlfDlFw0uus3WXftPBcROwU4SNa8IfxhZjQsAL34lSf+W6usv
P/8F0nyEYxLMGDg27asJww16oX1H/t82e2uFsVxj9bXEV7NytSRm6M3w4ln6kcIhHLjmsjuE1AHI
rC11xCpbBize+wMu8quRC23hes5YB8TmjahsUCutnpRgZ30wN5KTmpzeyZU4ZHY9pX9AVQOSQQUa
wU16uLhQ1UcHJ0FhCxcgZ7KrGAy5s1A7LBHUqGzt0o3lQXFQ2hIuEHSdGMa5Sl3n4a7cly3gS6j3
hJaajTSVSIZTd8MY9OfqqrSaE5+U/pbQXvhD/EsJ91bonwe0uhjctKobp4MilDGCVC4YHVEUs8+b
wchhYDxv/4QFuiOPxPf/3B1E5lEvzN1jNwnCbh9dpKRndFf90Mwz2xklP5El51gPB6Lv9KlobeS/
oENMfUPkVGqK16YEILEmLPDhGMg6e8OBWkjZ4fGeTU14EA8yno6T1JqrjW0vR8Xjqs/fDa48jKHQ
Y8V6Pa6ghCp5U03gGcgHqplpxvoaGUbBhsZPbJWYUJXYMk+11yw3Zi70pc6Q9VwjophJU8l5b5C1
F888OTMnvjflGXFH702HPJqUGtgWqDNyVYNwAqIEaDUsDrhpOY4aXtdy06mvWuTwlZdD/PYnfk94
u3WOyvU7k509rH8/1N2IPJFQkcrzdUR+CxNZsaQMQvPJjSlCFBLByjdIgq8mtTZeAX8ay3NknY7p
5mxqu2Z1q5/l3K8amlpWGwEsgeJB164Zd4FMhLuKVQRH/AJIIKZyv7/iB1rkRA1PPKcSQTGTmxxQ
KOrHAnr9VycZ09tLDq/3N9yOVSmZXURH1t4z3H2bZHCsNjtnVdBFjenXor3+rA+4UjSGBSecCPyK
TcgbEFe/ZT6dqxBXOYNwKCMx29RmAIVVYmcfHKRJ2YRaUE6tbY3aQoUxcsjZtgWI/MukShFtZItE
erpatQg8OfhK2OYKFU5Bg0n8Id4XchZ/ao3jdowCEg3oVlaCH3AAr6ZTbXQE9reWPaR3I6Ezt4U0
zCOsP4Q2dxbyqzhGHXBLqHcPfshnByG6S2NUWsg3RPu+cU0RUUs96zafrdKjkHkRd0dGiEmNmYbe
oaUhH059gEooi5xbu89qOOw8OlTl39K+TU0qxx7PP2DJ5/9/eLaAcMTa5gw55FX/qktU5i+m4Mhp
eoeXQNMK6BhRYHItPMZ60d4zMFvRNcqRj+ish+hVRc27dhIhZOlDpKKeE3OCTmMFwX9CAZ6zUeDF
Rai5VPLgw64BFB5bCGd4zpvZyqaV/DjWYguTFfRO3ldnp2q4DKOI+/gM56owC2DJs9zTbJF4h5iQ
X0ELXQKeZh6/Ex2OkBz/XVk/l4kiNKXKyT9bN/3viy3V3cOyRrkcFdp6rxCrkZ4fS7wXTU0JkNCM
1ij4goaypLrX0pbHr/jWqIZmmldj46oQ+VuWudN7pePzEDA4ZQ3Ajkk8tfDCsOOpGke9847MIdkO
OqJCjWpYz6K52UXqAKrmz17mAmmc1ZtETaRbTgBw/nNqA/8m/2TW47+4bcVXKD0eahnQyy7xS/+W
x0JeR0pEpurYRBJ656bUKrXMPArjzVbminJyHEXVZsEpWElB24BEHF5xiJfQwYr93boTGka28NUg
vxQf/qiGm0WAP3UUf/aXiaVq4tSmLwwk8XzBzEvmaJh4VvKO200hOeWrJ5n58xDVJIaLyOhKgCTA
JNUQFeapjQzhbJ/jB497QNsGthoxTppdGBsPdiKj09vVu59e57WlX/rA32QGKLpFDaSCX02mYcRA
QZgRSm++gKXu+wMcAP5Qzh0Q3r6J9ZPIlgm32xAei5R/fZLr1huiuLy5OwLDinB5j5c44iRZ1P/c
LINISyeSX5ud51OXHdzKgqfh0HWVNuIjEqdBtbXFpA35UxbbPhv1/J7SsNxIsMxm8oM7mmK+tazd
j54EYiiSB9shyLCLhsIGnMyf1vJZNJZBFjvHlOBLwbMpgXhd7hP6kuxro5jH/28bObTGjMy6Ynah
6ZHmiEv8NigQ95+c1CMajkdu0orCLy2lWTnxUcnYCzX4n/EDxVXW2FVvuHQSnPhPff+ZLBmnyUsn
j/fuDQGhKfVZJba8UZKeZhJAvAkiP1fmoRf1kRojgdL39lEGhS2+MRgEIqL5GhAVN9KPEFf25BVc
9HyOy4tO4xbzl3HPSDbPk4CdZYah5fDjyOQGUL+C29NeFgAdpSlwj+4c6rmhIsGDHoSpNKSqBoDy
oYbxllT6uJoHzAw9xxVYNwBnZal0+kdQWftrRzZgQWFBoP3/whRVLi47p7RUkatvTpuKpQ/AXjGl
YJ3ryn74Ao9JAZ8GxqpqbS2pdpK6sXAYjKkpxooLXIJZ3pRQbyKkajTIc7tHGXhZ7nwQhPcvEcwB
nGiWdBpOzj9d2qRBeM/MgfbZimggmiQLLgQVUP8Sp5fhcRF/k7yiVEvl9yctx0iEcSY30+kPdPgF
CeT46S0plWxYQn0b1JT1pfgRtjOW6v9oiULloFiESLrvXeWTHs5+DoSU39lhY0pimtFuUTZFCcAW
LDhZLcetkqzqFKXvwFpOxciCPMXNSSjQWk1zLDTQrBtpq5EtgraAY8j4Zm71VJJqFCgIFPpH4Itz
5krXl2hZoMOS53KdSI1OF1M1jHwkYWV/+AsIa59ZoJZr8Y+12O+u6vQDM0BonOuIWNE6pcpez7UH
plpke1neXKLhlsTe+2PaFLVHpiQ7G6/d9LNG44VJt82QFurSkBSOBlZTVtGxGDehdDytAw6KK+XT
+LN6J6X8/d9+hLPxMt5m0iqrC4THf3TK5jTxiPoLKrRO4gobMj4RYYFQ0nZw3UU4TCZoMZAv8Iei
c1BDH1GjxrtFhp3+BhKF9HRcBo+HnC057tW1PcziPnuefS+uOnSyfTOGK0nxsOJKKWeRFS4Fwlon
515KW7hmJervc7LbAUSuSFOjKCZmlzvI94oNNvHYCs5VprMn6k8ISyaRMUc4W1g28x0SN5d8kA7O
sJdCsFxhMDijbZTgRsquO60oVTHVKUP8uG8UB3F7i+F6oaMw9a2K+g+B9r37Kpp0FvvPnpckvnTE
FmFs9tJMRsUGVhCh+S7kOJmSZM7BGfePcSEkEno9azmu27c/w1sgIL5K7vsHgA/kg8E1XdMn+uaU
rEk2byntl+ZbZ3F9gmYoKWR4k06zIXxFngDED8ndrnyxsSzCZZvyeV9PlK16Wvk4roHJZmKPSmUl
BWCRyqxNLr4JXRNQ/AyL+zGB+dCb+YSxD2EnhkgF4kwG46OhQPUblwym5h29AnPi1SeDfIwRTtoH
mDwpAE48K15Y2FcIu2tPw97pCOML+KV1LJIp/ytNZ21vTXx1Hf8iC2pAZdiN0+ECcwh1+4v+ASox
RBgLGFNTb5ZPcgY6A9+5djlsmM1dw+zmc9Z3VQP2u5KYvNbd4be7gjfeAtNHMAvYRTWcxqU7kgmX
87qLno2KmO2RNrhYn/Ot2nQUlawijbqlbCdexDLk7jcWI8+j1CwD9KlL3mqVSosMx+z9LYDcCpgL
rPMTsyAG3WxkHtVg49TUflTvLqBUu/oJvxUQd31fvO1ox5Nrea/O55OqcQr0VU2NE9xmUvPtBQg4
TZwXhMvuOMi/ncZF+ULknVXB6VNMCGmaFoF79+P19M8ZIouGW+rcynvjvqvHgsRf1qOBpLSA8TRX
Wy2oHdwwrZpOMN8qgbHJnm24xYemuu4b+0zlrwCci0bt6rCdbNNKR7GKgp7m80ZchOFdg2A0zH6Y
qzTXAGWeM5kU03b85uxNlx/xRum5ojAc55eghPIPSMeOslli+fbyuhzUNoyb+B3fVPyxWdfa13dV
2+ISV+2qMS/uAwEsf/h3hT1NuGeUdcenV8WEeut3SUT0RjGYHRxm+PRDRPrPSREgAaFfTMx582Kn
ebMpjEP3MZhsEG6BRwRDYE4hh4ZxafMaJijh533ggLSyqleqRlAinbcj9BY0hYrIK8JITL4XwjHv
77FIWem7pF4WxcPzdgxOwzZezUd+Ro6vLiEzQTUdr4cF2V40kI3auGgw3kCH4Cfn/Z4bpuXf+JG8
ZdMGE6mLTa6GYwrvSAvR4jVCE6BVxWMW5uc69RZaEjxcOmtIXXTQScuO3IdysCXl0p4/MB0afVmB
/Hw0VIth6CVtqWTslcGULD1U5e/Ox2FEg//YzN0fkUlO1pgfl2ZjDdjhptuOpGvckkpKo5x90TJK
Eob2GhgSQSre5Cp55GlLPKzqiudus/cP8byE9JPH4ZJJ2tkwSG/ziEIpmmCnbd/szG3usXdRWmbx
DqQhzpXbsgi4dGufLCghjCtF3fLItPsUZYYOFLU7aa26VboB8aDpNHucjHx2JRPYH84/jnMiCOnu
zFK1+1XVATn7FyAKEJcQYiM8farDgA5KZRZ9+9D3O4VVqwG8YNWRlBgmhyoSd+WqZu6aZAT8BK7J
MdKkT3QnuJasCghoxd+rZbYRjF+dcUe/AbudAfzyWH/ESxSOfMFlHRES+fnMi54L6ym32oFPgfug
GP2NVz+3aYjSIVmAyBgeUDRFzq6vJ5DMAFVF+TQRAIe217YjwjGpqlTfRnVMl/84IkfNKS3jI6B5
Zp/FzlkBxKf3hPNQk0kv5a9VNX2o9o/r+kd+pdzeBz4eyhJcRdeLkxXFSZNIuv+rlen9a2phHmMk
ELcFLgEdOHxTyJFPTcVM9nodNsdpdbY5W6q1mz6Fh9/y+/EDMTx9T6vD6cJ0IZgnNqjsJPQorSY3
doQvbXUnfbAn/Fa3xLGmWO7quQSf5ZXirbZzCCMc0pdmkWVf55MBMd9aRzXbmaDFycpYP0OIJ/F9
F/6R2kR8T4kIw4SL4zg3pw3Ol+3NWaOw7GIiJfME6wJwJ8wu3Y9nwaZfItFHD5QGYGSma43b9iMf
4EUp65HiGuFKxwBdgJfqVVoj+zImbZbGQ98aDhfrA0mTJwun29eTDjZrNLN6HwHYmYB+evttxk5D
ai8y7TqKqV8jU+btYHtnmvqghx9hk1v13QS7h7kppdM9s6F05Rnry45fmxOWNBeWabJhzCnzwCd3
+Get891ZPU71FjGbfWY9M5Cb8sMdynp2Ukt//Qy23SBpTv8gUpHz2aMjnVK+NjqvlNVna9oEKIR4
L/TLl288AXaSG688EuFagBUR/3FkgrFVW67BKY/Juv7vbt+QeHJl/i4+WvE1CC/DADWgMo/3K+uC
CVZOeMUVu6KDOoSad9MjS56SkJoLzDbsgqftlws15bpK/dY9gw6UPXu+FHuDTfP8OP2MNocv8yQA
XbUqTS6aUI7YC6sJEh334V8GP2NeFDvePpktS876vsMlBUjRh4SHhsMZp31WBisnrtlUCw49FBvK
Pr60J6noWJPpCHjxbeCo5fVsTZtXhUvRFlGpL4dkgOsZ8LXDJk/lgxg6DU8bqZ6/lqZj2BSJs09/
p7v7/552PNG+EXHvkc25AZyHiiOhbi0IVu/0dbOcleTcF6vhgt333GOq/G+NdltiV+z5WTa9UNMI
/8Qm5kHAE+wUax/nu8fl7arCApLs75C1ZXMQbl0UnDUCvi8SCoAiRqlgJaXNu5S+z/znl9QMJUSt
xAoFbqf7wzGdAuL8F9W7QvsWrBAUUQOWGLEMMBqj7NixoM2xO3n5aa+7ePMxiC70J7RK4ClnmfYI
6Xr3CJ9mpqAep4oCWCpzmIH0ocBR4daYP2WBuzjvfdVdOZuUyzyQrtgI2WUBDERXjoHzLrMJ8MSo
nsRgbkf9Ae6VcMyJvOZz1bne1kuVW8x+eFtUdRJ75nuQtX2bWisP/NREamHgGfSgwkOeBilyPTX6
Zx2A6y0PS2WV+9sJ80hiPiZC/XEkPxbjigvnpnUsF1iYMdJq/bWjSJbOND6X0Km1qtf98w4Dbb0u
lguzuN2b8mUG0qb7jouOTjdnptJlnjhBoqV2vngF31EQUdcHtGE39K21Gy7svyX8Ci6VrsVxmuD4
EoR1gEnCcg6rTym7R+dh2+mJsfUGowup47RTyWO2vDo01iIfdQ1geBkDkvsqw6ZMZwcbmYM+LT/s
H5qP2jQZtdWXnaGd6FVSB7a1YAVhYDjn4BOiZQdvbcuYyqxdJQt+v6saVMnSY33VXq37eK8jfJBu
h4zGWPo8mneOMw+KRZZg2FTKkDneAHU6g4sQgf2AWuqsOkVslAyI1wq1wL4fvwcV6mIwNdts0Y2P
2U2xu1/czZ1d5KT+VgCL5P4pZ5ZBLqxO5i4safhAZ60TDM4p5RQ8DGt04ThrXsNdWIJlnDmX1OIn
H36oNpvjC6xd9rVSL89tPnR/eiNUqwoFFJFQ/3qN30PTYfehf2unn2iBd45+vd5itQLJchhhO54a
mkBNRTdx4M7qDhGTN0aTrlYZ3N4OBMBRBK+ApaoVMTuZh1RUXUjy1L0aRTNHL3pinZzmO3g6lLRG
z6GeQ1U2DAnXsoPSTmHHI9D1ekqhwgOQ8K1GT1fhsrxlPU+iwKUpkiXpg7q0+hLQg1PNMxhxy/V7
IjdbCOfmpVnotxn9gYFTeDf++NVNzuYuknF6e3Q8Nn6U47UsY0mrKoHJyXe0VnQDsjHIhFB//eOi
RCIGUzudgfQtZEVaB4iys2B0+aZspy5oMPDRQVNGQ+QU51+UsA4V+gswKQcqi4Os2bZKbE8FgZxT
SvAZSAnsSSige4EByw+CJXj2pmqGJWTnN9nTWlpoLfzltjiJuE8srVMg2E1+qgRU8qFq71uYxtVz
sokptWWG3Ds16Qumwowj5kPoEiKC99DnxOOMoO44A4aMrjmA/4pWn8jA81hb/mHQCcNfz4ASaQGe
6olCOkH7jsQuLRWgwQKye/XcLY008ioDOzQpBUhxxmb0xOSDB28ORzzxR+UoRPz2K79Ic0u5wPFZ
2WgmQbwZP7ajv0EjleNfKEwQ70hEoNF65cGsUnYcv9rQ8q4PiSfhIBZzak4AOF+rl53jVTkU6fDg
WS4I0PmC16wWPS6LmsO1JioblX2Xy2iDb+0rAQVslF4Q0wAKWpql5Pnt0xKjh6jym4rqYbNSehjS
6qkmdxjl09fceDrWE82/Qsu6a01zJ9yvm2DqdVQPDeNuZ+QlWfD1J+pBhkj2RudWIuxg/a2nR5Ir
xYLbNR1jUX9uifexHAxcU4sdUyZBsuqpmhq6NUwparZFfJDqU0vweGWLVE+2JsXg75tKEIB4YPgZ
iC2ylws93ehDOFDiZIEdba7hEOXgJkPM4gcHaCjLtaEEmKDcS/q4bH3a1Uo3Z8NBaD64VXdkeijx
OPUDDnFHjeKf1vgZ/CSCefykJsjuBM+B/jNpLY6sckv/vCBz3LkPUSqnXarDEd4rQQkguyJ7nVSQ
6cNG9f7yrlXPs+dLys5sUOVWGO7a2tuvvjny2pH28BXxsnYLzCM3V0wvtg6/P4QT5/k0cws3HXA1
MD0de25GO9onyCG3S7KLEbblhvWt+v//7JDS1aRMaRBNzULj4ZRUhomehY7WfYeLeEhZdoFSKYZN
vAqNTJkmD5+b/VvupwnQwi1zD6MtFrFQP+ljM50tp76nSX+fREpqWoDxOh89ZucEQn9WoVexAl99
TAC/aZKJ5uIr8ezkOeD10lCST4ItbqvVfn674TDARqCjyG7BEiBQtSCkl8qkkI6j56BX174lD2Aw
OukpOV1/RfjQYIeajpVUTqBcQo4xggcl3ZASin0JNPynrfj+I5ZNRyDTtYZjWDi5bQ0uWAQ7RaWx
zvPiuIAV7tM0qntlI25R15EFq+sZkcOeVNlx0WODhXwLyC8MPn8o5xCIwh7Esr9AUQkT4GxNDMb3
RZkhL0HyN8Wp8d9W/jt0FAbNeWwUEYy8CXIa+u8WQRiQ0/GTGRZA/efGvl8wGgF/XVLJlDvXtJAl
keBi/QkgNk+4QuXU5rjM0gqm/L2yXaSd/G2Ce5BsbHck2zPA/DaGxTPyZwpmQ9ZCvbLm0g57zQHD
naiBA5+7aJCXQgG8k6nPsI0TMZdjZam1JmQFof7Tkj8WGHGjEAFI5Xe2xEDzGuwihkxZ44Cqwqlb
uC4qmT61dnJ07eo1eeYGk20A2/mnUQUnZkWWc+86iGFuGFT6fTR9dgumx6MK4r0duF/UzeZyPKXx
CfVHzMQq7HbFRsLkoIzPmVVQWDERfx3xUYSY7DOS7Jz7Romk4sdPvgoWitEbU/Boshi2/qAUzHDM
LaIp3mmpPT5jgGFOF7tew1vm5V50JGkWs5C+54c2Ev9kHGFaI2C2m3LYQ0UzTT9ptDPob1gX13kH
mAI3tEhpdF3n/27pI+SpSNTzFLii9KU9hSgzDSk7eumQclsrYkSQm7wb1g67U5bME5+pcId4yOO5
njeLQcdRSWzjH7hu25OdTsGKv1FA+vETNWuQ9Ce+DirxorOwzJcB1WZpnNsHn81lz7FOluw0vgcm
lvqdeoUwFXm9N7hKRzDd89XgVGepMrGmKcAENZAtHqGLDterfv2p2e87Yaf6401yH/2AG45yXVdL
Z7x3xGJsEjyx01VgQndVbJqAHylaYPRtTtUdbJBTAOTCUrZfFtYAr6Gy0AhJaCLe6RTnB5cmIHwo
hajR3VuN4ZorPAi/Kmb2GhRz8Yo/mkhf0xzaIc7o4bF7dP19HGMb9B2lP9yh3ffDX9TPTZBr1Nf0
t8Vqq87csRf30a2wn2G9ZkZj7Jz8aBrk232H8oRs8J8FcHL4NPs9LCa5nr9eM5hcPl3hr1cVAmwB
bLq1R+iZYHy2gPhdhl9as9m17lW2Wq27ANtUdJmRWgBdAoiONVEuvffyhCaY8CzKw5OEx6iDELwp
ws9guLmQKYskgC7OaoPXe94sMbH40YqmsfZvlyACY13/YfmhG+42vBWhFHjOvx3gUCjiODFn3+2i
MC8Jrbcu7a1+V/l3EXWyFfdinHexG0Kk0G5kf0ws4JTdbAAdiTAuV6+oKtxTvNOhL1TFn6AL5cGn
tpN/ZJL5LZ3Hcju7eE4zuWIIXFLil1T7pkPHchYleasHp8qRwgkoC4puB7YiCgcfNBbmWKAKq4/D
axR75VI38zvEgEIl1hPpqf2FUCVgb2l4fLltZuSMrav+K4Mnnn1lcP3sRVNLEJ7nDAFtQ0GYRy/3
BPsvuY76Ww0GoJo6M4DxQNDVeZb2OKwbuzGZyEoHKlMzHJ3ogxmZYx2tGGbDmBUL6IxtCnrfEtlU
9z95ZXNsNkirhCXuplF3iGeqHUrNAzxUTtpsL2JNa81MKvjcSZ6/YYP05AE7d7BJ0vHIu6uDLM3j
Jlid+glSNizWfyNsdpgMJteIls0Bp6LdOj+RQiJZHkt85v4H2p5D3Om4Y0k9p5kD2fMnq8v1WNVw
7i1IWo0kzQ6SYF0bly2c+4baF9g99+aZjhZvGNPie3Z7l5gRURAtGkvE3zZ7+5KOcs8FSYAWUcnf
x58YpLY/VIiqO8whgYkJihnrGvk2lZHduj8Z8wKQoIrGEpLYvDUx4kjO4E0e63zgmlfkjw+vDiMV
WZST9hYO9Ogxg2nkfTa9ihWq0Evj1dtMr4BUh+5AzKmkW68s8qmcVxQdfX/8UrZ0WXgsLEisjUax
UQVXg2C1wScYCnAt7dJN/qdGe4l/hbGMiYKmcw/atoyrmOaQKZhmR7nIKx8FCsnhhMxOarytqA3z
ubGa29Dqj201cocZf6ivw85Fs7LGNZZL5C6bDaMKucXLs1I3Jajys/jgEgw7mwLjQcC4HNp5gOYG
iGYQa0AZCN0ggTdzBok5TU/b4l2W/Pdo0pXfcdry+2LuAAs0GJvI1xGYZiv0pq5WkI8MWgo4IqTv
7TuPCKFK4gfDgsZNwlqoecgDzp6llG51R5/ZpI7CfvnqCGm4Gb34OxsGl6zVQda9fEmE3pnrGLsC
kZANME+F8s6YTAEgQo8CsrqA285JTADESUYY1TipLX1eFyLeF/D/y7KOANFcemDyCSfHuaLoI+Vt
FVN6WOZAOc45QQcmPqeJFyM3Xf0i+svFzCYE2B/lQvISlNjArW5Yf67Iy5xRNF+I+3J+1OOF+qNT
ga7htEzdhRuxGhQ2Dl2mTJ3Bvd1PyhY80StYdqSrW+6wiGMM2oPaNevcEFU4ifYh97yVzlo91f1F
h26BTzjoUioQDd1Ii68rynUxSAGfcp9Y1C+kFSrNnpsq+f7N4Rcmy+1BfD/hleiun/t92BOkLu5Q
bSxS4/R0Rh6rBhhDooQLruo+G4TLLrngdVpaEPqxJ8HCZqSs9OyXXbGmQwT1dMFDpoN7LDF9EMi4
53sI4OcA45wnQm918ZutacAQRV2RTee8ODk2OTWbOa4kRCq47Q0qNkoqqfBBrmTwtvkjZd9hpMYe
Nvw0QtNwOtwTFddLORjmh6wsgMHTFiSW76YO/Lld9yTX6mDEkjBLwrh4+tuUSLY7OiIYam3ObjOx
ylwJuUcCyIKAd5Scz67oJ/ijcxPGegENzMqXS5B0oknN6iky9G+V1kdfVd+GDICZo63owGgRHOVd
J1N0fb2zPoB4/oRydZdQ4t+iiJpTtlzUWBRW6l4Gi7Fc409GAt1RD+KIqKJp62ML52SdJsu1z+lT
HShFMdFOB7JjSNcgG5BI+m6G+zEuoD8B5LoPizd6+vWk8FdJmAGcqKmXTpWdi2poPRXaEoihFS7W
4hLT83hVBiQIBVXDUCq2H/nQYBkze5h6ThZGZBX59RVsHUxH5NGdXE2Qk6KbENGZMNE/us41tMhq
lp9Q9bVeWO8QrIBRriyvz0SFba+w2aJXS4PWH6bdrMAqNVvSZXG4XgMe0J1QM49JUlhSwemLE+fe
dtBlNB/NtSFjSZF0IC3Z56PBDHVTzJnzhRmHcunKpXMm8FXTdZWMaSx0qWlRn/UnV7FCkV/5Ue/k
Mv43hhBqoJjVQsMTLj6g4N51gWD47f4QzkbFYKsmEdBLUA1swlTTmH8zb0uQaf7oEwmMqOodteWh
0Knd2ipBl22a27fj+SkrnEuA0zWsk6edjoS6bMv/jF65FAjSnC9aZJ+UkReZHZ4tz2iM7ckvUezf
f+de4KL/92zmK0qup0hDLfDLF/skX6KkSrt/25xq6UIQnMe9zcyByK+mFfjMg50lWA25FH5tWNDn
CnCWKKtPVbCHv2gAuzULJ2FgRhTueVtCpZjGbOlxpJ89aZrTigOor6aepYOlgyi/Oa0HNQiin9KO
h2FsUj0G08xLAJbCmFoHtQ+Nmk+oflCZ6cl6bOnhup61nCDdvUnBxTD9Ufd1MaKXiyM6o+657tty
PwZKYrMkpW0WX9yPVSuusSEUhBHJsWfGQjSKEs+26zrFsber+O7yXGDvPOjSOkLJIKGj9PauI3PB
IPmMPUteEJFBlwyIJ5o5GJ/X+B4IBGTl56kCyWfL90J6FANUVzcf8OnS0DOa+g+VaO8QnWTodp2M
e3qbZm4cWxN6yMf0AbDpWcFaBC3zC41b10xUfLK/gFRemhUGp+6IrAQZJQln7nKRxvbSpks5+9lV
EydAioPQZEtqaLqG5DHirdTWBHYE0XctajfpqvNun7QQykGkMVXSE5m7NSDbXDPpSaunPEb+kvxm
DKwb+7JkN1wN0/oVPYhgUWIWexLUZNrCJNYW2+tkdS5IMd4vYeyp74+BeAg+eGemvV6zYZShcqco
h7YWsKFfoeoVx9oODebODjbg8sKwgEsLK1p8fvddB0B7Ge30+I3rvMcUSiR7wGuYDE2L7iBnDBoy
NyGde5j826mZ22h2EpK4M45VxyN7UTkfUJ/wzDCciLq8ZcoPHJpnn3EUdKyXXED2x0o8t4S1cdNl
fu9aLsRGnFqf3Qbo292zjONZvNcHKOiSEkBVW/VetEoWy9zPZCYYaxszcoD4cbwm0IDOL4P0X45q
jOxP91/OVc6Xqcm/0+DDvhQehi822LjcbWUeqtWfYSCaK8e7iBb9ARndf82jgDrFSwxDC2TS/RPW
fL5iuTQTYIG0JASFi2A0gNQr3Be3qhDQIN3iWk+66dn3no7vOBfsUIooMxdtWPnpnfR64nxMrWvP
9raPKtIZ6nqnnfIoIMKm/rk/g1iuysibfmAiS2XF28H5+5whxXU6IfXGFzToeCiLwefqrbP9gipy
dO7YJGMr2Ag9lIf8fY2BW+W5Ef9vIhsLxiKoBA4hVqjzY7N2dRLwPs2pQR085DXIu/nEn/FtU1XY
FQj/Fh55nuWAdn890sObgB8/T9wB7abvfPj1hiDKRYGO3DKrXOSa/bvwfgmwKV9YRuCCD+DcJJBt
5g6JWxGp5f/zmvoikOGjLGsjIN5T7OWI9Q/25vs6AOipsuFVnjzfeSax5dEVNtH77IrQpqPUgPEk
gWTaFuy/2HyaUlBLLDY9A/UwgWzhoISiTtBvFsbtzacbu/8v2QUufHa+4S1J74ESg2d+Va8sc62s
leHegg0L5idhrWQ10x91Bp8YKIkOLODYXnMmuS6LocAKHFgKLw39P2pnQ9HNUOn4tX6P7fu03yld
h4rGBAY2Za7t/QQuEn2pt2PVAt/w1ebHxuoBE4vzssrVXRrraMdIzUBl6i+RGj8KwtM9WsP3Aacb
MuMW71Da2nlgqkAQirGvC5bWmqk1sdqI5YnPhYp47Ne6Sgljyqj4AaHiB5lZJNOT5Ghs7wPmVnNa
isyB63KxbgOHY4+rY51rHK+80EHKztd59P7iJaQ2OsR8dIgmh4Z5YJUPd7wJQqAjnP5+IPpAzGeL
kh57RmBStsRZIjxIPGaPXEgJF/FzvKhgukDVuMYVNzC/o8zzqaSDk1KQ/TVeTzfICERqeGaRi7Gq
CiwE6h1SXu37Lqz1lPerSloWQX4dcgreN5Unxw3lceeNDkijpIjLgivdGZb4VITnmbc/cXgVpmNG
eem5AwUUsWiNXs0LkjDhKl5gZQ6OB21emK7FWNQoKqZttaeOGlFLkVpnw/5Uyq+5Od9/fIRomOjn
l1sXd3uMH12nnc5G6+hwInFMt1+LMr/vXNm0R7HLQeUJazROwfa4lLTJMwkiLGI9/KAt0CLVKUPW
j87R1oe0OAXmGm7HApSTJlk94mNVT7L88cmnPmeTlksferXTC0Q+/l1iWk3c9q9RIY/+fK7oSp08
cPlZs4SHcJDvpudY3amJWI+K4eUDF3/mfvVol97qUgnuHpCJ8HPUSLsyGfO8eaOr4j0wSepds/uu
uBEL1uHUIeLLlsNeygVtWMKpQNeRRidOiRiLO58RAUAc1LjmS7xlYtUjKY3saCitrflFyzavhByx
5lsnF0/1FFb8MY/YRui+BkLpBhE1uJCtDk2dOuwgBRpF2dqIt9B4I1WQo8Fyfjt/FkbFThuzuzZV
MYpZ4meFYRblng5F2rFPHCCBT0Wu7KlL25YicLVco9Fa0hzVEIAfRuHXNdPwqsJYKgj6oJtN/Suu
fFGyBM8J/BUOESmYe+lin57wSlZrqBUMHM1TB2WlgfkgBdtr8mK+iFvWF5b3QJ8bPQFYP7bhFsp/
wN9dbBry4F0/NYCoG0vBk2BmEXHNY/R+8PG+sAPPYdD2lrRumGfCIqzJJUI9qVuIl5VARuRh6ezS
513crhh5SEN4KyUXoSmaMGrJaWN2fS83V1PpxWFZhFatVd/+N8c036yDZUbc3gTHVn4xC4ib1rD8
ekST/+4nXHV8IjCNPaR9ZARTHaVna3QBsE8PGe27NNBpp0qC4UTbFVJ5tVcDdQZ8X7mPrz1oLcl8
u6KiIBShRW1OHjNlmkuG3rWGWx2xOdC85rO5oJ4koXVkgyaN+7g1lSheBsyM6TUfwIhXZTaDUg8p
xWA+b2iMfwOTIAx4X57S0Vhs/5T2NWRgnb98EzeCnq7ZTXg2QdgKuRxc5ZAGlrI2dxuDgLYWiUCE
c0Z9NcCwZoj8DJOroajI+IUDB9lP4Gczo0v3q1uSG1doWASnKjd3Cr4X1lhizV8LQmf2fcaHxuL/
btdSD8ueM8YQSrpbiUxGm1Jbqeh1vKZVa0EHOrueMF9gpZp19J+lSL+zcaEMs7DxC7g9m6GigDpf
um0en1iM5pE2aHaEEMqWR2Cz3rzo5WJBgWiWBKHJPfGELX3zp2/ozbiJ5tN0cTuwZSAkA7uWI6FG
zM4xHqoOGpRPHtcy/F9Zs17CKta4lqTJn6sBitzkLinq/N2np3wwRKojye7/9bEcvDZY4Rh7ZtkB
wcTd1UXP4fD3+xbD+6FZClxok7NQl8c6kMqZII57Xfogs07WHSdzc+p4NJgmfOZeGlMo9qzWXwZB
TDG2T11Z6tYCgtVrwsfsxJkpcwIieGlFu0pQFNZZRZtDsr7VfdFiKwrN2lQMxO2yG57azPkEMblw
9asK8Y5XXc3AYBTef4aW3D2GtTjvYb6gaDZhIcW/dXJARPAZbYZ6vlIYm+VaBXaoIU0l7TF/eyZU
2HywyQy7EOb+SADkh5YqTcKkMJHst55gbMOUMX+5Y8L6r+KmErLqZlG9hWBq8J2vS47o4Abj3LmH
7YIqQ7RoG81V5KB6jeXPuSIuMKcfeeUwnwAq263zuffyAQ+BapYpfCM3iVQz4hHaiUtvp5w22ueO
8PzVhzHxuItbIGvMzO32wvW5iB2o/I4RAfqpMeBryLIaAufkeRyGKzaHr794viDcGIg0B5Tb/ddG
bFCFwV5NugdOfYlVvouq9VHXM0NC0CE0wJouYzg2cnscv30J1ixQ9Waf4QQxVWCJHA9Nlusl0Qkm
DpbHCMdPrIlFmuOcK//hlwvl4vds7Eu+YxWurFziJRZoQGVKlbv9PHYD0A8lflH6h/Ikq5h2Xly1
2WV5iPIsH6O0XOV/sEPgHT1zFBvzMFjj3I9Z8Mm2YoQ7xt6LcfkqWKirAe7voyfbRddCi9XBTWz1
K8xw+OiaQrHeH7Opp7h5KeXDx7ElOWzxgJW4Dp9f9OSyqTO+gyrpMchygldhFshlXYdJZFyT9LNw
c+64BEB9PqVesytV6AKv586NTKOMgA+smJScNSiw9gPr5wOTuY4ZPrBni27bn0cpI7PCdonjN69m
dkYK8Tkw2gdri8KlQkYEhQPRntRIt+LMPB8jawHCXdA5594m+aarK1V3YpQJwh9Y1fz6qdXRtH/1
WV8qJfF59+mDxtQugVeRqeXuzt9Kyg9gPdRlUgc0bHf9GswuJ7kA3at7apN9+6WZvvnzraN9fpoE
zhG3+y7t+6CW/uDsz6BXsQaoH2VHHjivI5GHjjSjeSmWLouiaqsG2h0MgtYZ22c+Pm6h+qj+fHq2
5COn3QziKLsSUrrhBzwKyFdGprJLJKiO0eKvzpO+ASJgTCbOZ5WewgSILNEJseaUqXmLBfzvb6Rs
DEfDt93U1dEf/InFa8h1HUPjCh78mDFxjCsIHJryptv3yfn4RC+2vbnK3Q8sgHfrKbpoyiV5HX/u
mvKKos2Z+55auTQ/EcRbXunTyxa2zQZdXu9ZrLbg6iLXCZH9a4cv14E6gfoG9GAQtpvW+sFls5/Q
GpyXQQ8chrWrBa689YLlzuFb4eEJ7ZuQiZpPuiJvcBO2510EuO+vE3ksA50/My/nsPTTavVH51q6
0z3Zno7+Cs2wntMkcjJheKiYpGR0/omXBQ+vHsqoTIpxIvZXVxM1S1KbeB/FU33QWaEYJIXf42UL
hh7RBj6uMC9aK4BNz6v2l00jXqxjYsOWib6wIdMfZ5nt/HYKXK0xEXfEGKnp7qvLkCmQaGio039U
dgHGJYOKF0JcJZW+jPIiCRLo3g3li+zH+2XZ/IHPKgSMLbkCZdStALviN/5AaoBfnm0VXutdGZoF
W4SzT2q7VXq9THeCVlhUMg7Vt8VUxk5xztHWR0Yfh0jOVk8WjllhafrsyWLgAuHrU/1FL8UrZKhO
oUOXw7sYnd/dWNAZhz0Rp32wA7S7NTagl4s8T2nwO+eENhBgoYXivOdY+GkgPFBXft3cK5oJluub
7B0369ragFe/dsYvoxlEbIG2LSpchrG0SIRHcfoEXrI6zmEHUwo65gtZXyEO5gTRxg4jmeMApWe4
t52PA5c7DS6aIMILgjxay0gMM0SG/02DJ5U0BDbtmz2a8P+vqQPFTorQXDGOp7zeQFumUDa2XqIy
DYZEGxcMXMDCSsAldtje9TsvDiFPJ//ZJb45uvI+kNSicilqNeCwOMM5aTBNZ6in0rbBQyyz2Wxk
vm2BSU3iBNfggOU7Ytexd7jSGq6/tKLcWHaXj8q99I6QAdurQ0BJAnkqZn9xgy8tifQCYMoEVE21
WO+/LUw5YURcSOwa/0K3aR7E6L760Cv5yTT683VB84kPyfCLZL5fuAEIEAQT6jnYz9NaBH6GCJ9x
r1x37kjGAXOCYaFgw8APUvGWHEH4ewS4mxTWl5w75JLoLXklZTby0/b93JYPfeLF1YaQlPAAJBxW
qsmN+0Eyum6Ht45Onrb2jiC9bgEQ+cJgGDPowV9q7YgY9paJQ66UTdf+GWw5U3u5VPT3C8HL8Oc2
uhpeJADkBSCZXcdfcqBP4SVNmUIEPsuadREv7Vg7tRJW9nEV4qzTcdE0ER/x6SCtfAKLgQ5Ba3gz
uYjm9+CFGFBKyUAd9uPnumv5YazkKHhMFik9m9YPzj6h9FxtNSkgYFfHjx5kVnpIWNLkUSe7I1fP
CfB9AhnUunsdqJ0pPtYOuP87gdx88DaJ7p+n7oj4tcNDBXUcGaUBstPvoosiuzKaDicScQXx8iIy
OH5Yktt03wrQk39ezuRBBFv4rnw0v4dXEfrS3NSTc2BiLWzrAb+Tbm5X+Z9oBBirWieGHdCFaRB7
r3YPWqWSZvcOOyMAMA7FFiboknz1YlbHFEdKwHg2tXyOafAkYTXyP0Kk7PVx/QgqD6UJmmapuBxG
khuk1DoMe+8Ih5rLyLML1iUpZsHx5SQ61jpyI+ii30Jj84HhZ/h4eYHnUxa8gK1m9CTY4Wj+fYZN
qZBvI9bnbAPMg1aTkcalD4UtovOekJ5rN4dvSDcDl5RhCRqwRzKyRHyOBYvJhoAUj+c+V2jJiMhZ
BZUQs6izyesFLeXbNdo8/josjLHRYDXv84EPL+xEArbnxokvfyKTYaQiCzhp6ISAK/0OT+Z8peLU
X6TdUwvv+tznRmy8ad/7M0P/4SV2Zvss2e0Kgrww3eeiXTetYU9Whp9I3Mw+atmEDhdJ/bmYZvRW
SgvwVanrq+yQyBiRzOwaPRXLINpwr+jX+RPZ2VfQJ2wINmRKXT2/KQ7FRnlXkBEe0JAH+LhJczWh
ZN/ZmKYZyuabRltqE7uvv54o64sYk5WbDHpqcWgAugaqd/MHMMQ7Bos5+lsmvkek6T46m+RZCIJe
CiHtJwRFO3rsPt4ncWUDwAsHwJkRLWR681Reau9121JU9tjmbKdYCMHWkR57lHjOEp3upWaoDoyb
HRYYRyTKKQhKPwHWt27PM2a+ulgdTjVHqNIEL8sDxfG0V31B5w49Oj3fN8mCMW2/gGndxf2jnyi+
PFe8dKhJQF6WmcLcYCzPUeLky9F6k2upkZHlBfnCq0IYaCWV6i6ADgipEOIEZ6mBsBnPTSQ8/K6F
NKfPZoX/Xh15VFwUi7YKZG7e9TdffPsvl07KT+iPWemS9frRnb1mR/CP40ieBAfkTZf7sN0ljqIh
rHRklIJ2fzCpungiWlkabeb/5LF+aFqd8bpsaEpRIjSy93YCa73JJvWCi1Rd8oXPLD/tgWOfzh4o
mw867ba4dnaUOedHgH6If1tQ81hZADFhltIE+fyYqV+cyen+MREIrOKBK/XqbUFRxQRiacDA0YTx
oQcni3o0atfsRKAYTmFxu+DmRbt67Fh/Yv0hwWAobM3BJ57grSNirqfMXA0mpXo7Oa1bufGV4kdu
nRdQqgtaB6Mp3cpwuWdBHBZuyj3mGunX2PQGV4Esh5QZgaHVQpfyCmG0nYPEomkDWkYGuA1HpnYa
0hzzgwOWrOnxtpiFCp3v8+x5umJD+kUgarAOv8EkZo2iLtliEusvM3CeLt+26x3VYdHcI20rUZ9g
7T4JvwdqxMCoIRRVRTWpj1cEVOq55JRWlGp0VEcCCMRpbI0rddInRhohT5Z+gKR2RhMRlYVfcTBP
vAc7ruHdDAUngOr6nuCydhnthYp62oONpcusq2evX7tGRitslYzx+Mf4bB8wqSSRPn/iBGubiOdy
Q1lWlEOILH5ujbkqKayimbr4dLx5uOCldbFncDPtMO5sK5GlWEFnUYXJrov3UDTckU7HbplG2L2D
gJtMR8pU3evo0E0ozixPRNgDr9DbEuGut18/oiNVXAaSeDUXEXJNQjCd7PXqWuzgV7FCjNqPhDr+
YyKBfdyME5a6jnsuA+Q9vRB/d/f7dbuUYiTpinIEiMws0MxW7aTDRpL1tihkICoNe9y/lfq4k07l
LbjXGd+F+/ZGPlqIaD9yGZvC0ITofLo7tomjylqi//oLHuh4HRd6qUYy3T2JlsRaMWz5Kleag8zU
gh9aplmC0Kx2atHnOknQYP/yme32UEJj1gxFeBlg2iBStJwBhPVApR9G4N59VcPXxEaICtduANc6
6avXznWG2qFTNVPoAMW+BHi7AEGL/lsdV2WUCjs9w6b6h9e5bVKLsiX/e+CEQuKinCV06xibtH5e
lZmiTqChof1dsq9Bu0CRPumI8ZM8X/mZw8zo63TZC668E00LJqwCNI/s46jX9CMRA+r49CZKBnfS
KAtqlZV8VLO1wMrYYRptV7RDt+hONl7NzMLf6MhWmK/5hkvRFH/4iP1fdVQ4xp2SRdB6Q64FyrzG
3wrcFjJ6cLTCowpnHJH8v15O/ESv4ibO7dSDfbghv5RZc/xGea2y3FB11gBHB38nNofdoYqhlfuw
7/kFktgLiIQJWb6jMz6nALfhs6qq/NUF+ce++r1uZ4ZXtmsklIKJ/Y/hzRdNTo116Z+H7iyMsETL
UIuox9XK1SbXolWYg1g2h58SlaDnXEV2IaouLqbmHdFaQ4Qk7YfGBow+/sZeozDWjrWW7x+HVgnM
FCOK4rkO1lRXM0TMzK8mduq36LvUO9fSMI1BjdpejV1vGl5JHcgaDd2SX/z0XVvVT2tTKcXt6XHr
iQfkgPg8bT+/Nv99PLt7Y/x3Yc6b83QHjGiX/DljdBkLCnJLrGA8YSwuoJZuN6Prde564vcXSGWE
N6bEKhu+5TXP3H9GDZTgna1h0boQ7qVhrZQp1XAVSZ+VoR9+IAYUCyJtbphkTaJM2PvYLCHJ5zIi
pa9iiObuoNV5knm962LdjtDSqlOReS53CG1R7CVU2OMxIqw1ZMa+mg1CmhMZxUv2Vi4NabImBDwb
GMMCeAOAdquqOZTL/5IxWxPvqiD4c8hHWQlrFNuomNyCUrrWL9ccJDZoiz3sqppAtf4heYZuS7Rs
Nm90n2NVFv2uq9zHpLIYj1/SehrLjJg2XSNtV/W5Pz7nMvLm6JYbwIjkyLt7UqgIKXF3L+1/IH9n
+QdghhJ3xhRKr1Ue8s0ww8HYOKt+pwPKHBjVqqt3RhHwWg7RZQedEjln9J3pTDmuRuKQJl3YwzGU
f4cB781p73TuRVnAvQFZ9WKqPnDYRAHt0cUl2uz3t5LxxpYqCVkSHd5vkIFE/SQxjmgVchBQvHlh
M/UvUFhRRf18D1t00RCoYQRIGX16qZV+dAM9fnHdowPprIRu5KgMvYj1ek4I210zUxRVDJpUaR7X
6Ku+4ctfr9Bq6sq6r5ySfbxciMCoMkAGHBCl4RF1hTfZo6331RhJ75q89/WWyjt0hP1llQyQnaqD
WLtXHC4a0ukB1bnU/ACYccqidbCwV3FoYkdjhPG7G547CwzPqpuEO43j9bttpmUQE3+FXQSanbEW
H7SHWRTfzrKNBtYgrOdJm9vUNClCANMS5CEGq+NHXYTS2KMZxR2t9KqX5+qbmLOUa6gWICiucYhw
6DrUaQ1J2e3phSSgGKXCP+WJ7z754VFCPbwGfaEnwymuBX/5Y1QZinGxj8EbnEfuxQJgW7+NOVuP
CKuaUop0ewAzk40Bbj53mmZOyfRRH+DWLxrQAY3d2fR039X7c9NElBLMjTY5c9KOjDTlFmJgFFj1
7qbNJVbn3mIjCRXPfQdy/rAnm1w0bXgCgwj0c6ljAnp1xZaWiypH228gMY++c7RasaJSH1HIaHBx
NaBC57coAPQyA/rw/ChGai9Ryg+SjgrTeEwS9zmLIRhL4TvxtoWekVcnomsWeHCaX8wudna9Xjb9
y+3UI4vVuv0JLP/ZKcDROMqRbthoPEnNueYMtpvZDE2PiPzsuRVtAIWV9L1O0zsTjIoy7sT8vkPu
0jri3TYcj+yo40+eD2U3GSVfCxd684fhGH8CARJGmdhBmGX116djstuTxN/WHyo0JZShPAk685xW
ibSnoSakQwE8T6yeyn6fh3sMtOIA0L3NjCgm2mUKG8feCMBzs7Bk219VPn9yxMd1WtU7/GTmjQKw
fpAEvbgqj/em8upE/ca1ClROAKNl+iVRcg0Ee2ZNTez9HtPHSMbGh4PR0M9Wxf88AUNzgLMDUtki
nQflC9kIxxO99lUUC4egdsEjpsDCi4HPWfZhpadR8zE3wy8f/MYoocjceO2YHgyUKfZYPVciMxr8
tCz5DV1AL7ZWePIUS45XZDyGd4Q0bVogndWkXfCt1t+mCT6J51lfkKRarQkxZZI+3lTGUybIky0Q
OrG86jL9+h3dc/RsmifSw9jRWO7dDLfBWhSSxQkajyBUNhvTDr3DKX/Z+Fg0VANIT3lajGBskls3
M3Nn7ZxRqQx1AdI5O3qZ9R6WBqzbDjlhR3jWAUfwLDdwbJok9HF6d6XtDdq2o1s29NfWxsNq6wpo
YuSNivMosb32Rw9LT4ABtG211qqlO1Vv0fKRkzQHogRS/KJmQEzlLDa8VqRT2FahK743y5ZYArd+
9HM/Ndvn/BmJPJ4sirxBaf88RzM7HF3UzrRN//lF4ENbLxOnFnJ0Up65jCZwriSZY5ZWG/Jl3Uf7
TagVwCWUXgGseGjoMyf0qu+Hnj77Aec2A7tjLCgN/dejchXNXNciv3DqvwBlBcPdRZG62lrwvDez
nOxMmRj3RQj+idTGQgNUL3qc8CnfdoXEghG/NflJ/YU29corHMNsktOhJyhlUGxBhVaJcJODKj3t
q1KPRra0O+KG4OJJKIPg6TZ4uHO0W4pAYaPBKhuzx5/WC4Oxvfmeq45dxAb+NM4NTEQJWDsE9K7R
WRcTpb77yAFmzmooZ2Le03Ciq4TfQMp3R0Pjh5SeQzYvQ+YIlcBG5sbknIFgOouDmOLTNWxeZI5m
7EnjELfH8oc6dAt0CF7Wj/ItJBk/6XbjBbxUCTsCifeSCgimBKgmCpiMSmT3epOMeYNo7a8Td9Kf
FD5Rojvsoyvt4/ql7jLj4PsFcqF86x32VXd9t+BzFqAPE5VwPssKf0kYwMwpokKq8g4hzwXkeQqj
FGGeuDy/J8hrz2yqIks9uyGm5vjU6k5fuEJB55TppM/69Li4hR/9jfevEn/Lk2oZVUELdlhG9BZ2
yz1T40t4cHMKNsgHKfL0Zf87Itn8t9DGT9ewSCTsxrvbpjeTu8QHiREIQmgXR8w1PRUVJcv0/xWE
W2RMiCTq6onGIl5MNGh9tU5fMqkk1JNo1ogTJKUzPM6iLjAaHuUrwu+mbUXFB3DW4uT9EJcv/R2l
eKcsmC5AK+e87XzPaJNpC9scuXDTIh8iIpVDTjsQNFNUaOzPIexuqziFSBlFNpaD35LT4xOTPhSd
sZ/WeN6nRRE7nv4zM8Nt7ZiRVQPA+EAz5U+LxELv0YZF9y0jZhpyaxdrSdRMY8DezDubXuS0n1ps
C/NJzuZvQdKhj+GPp/OpthW7vhUxhEURhV4O2AfnvLT0UXvg8I40Wf3EH00ghTzwIE3x1+59xs0X
iE1Fb+RovHXypoEhLnDcQY3Pn2pBLZQjhZj1a2VJQZFXTvBQMs0sO4aiXuEx5EeVB2pEWITUJxe9
McBApi7usD8qxz2HHnaJovdLeuEVfmttWyqHUi29Dqvzbn2FJLFV11VZF0dRG7n5kS4W1CB6KME2
te5GBO2LyGV43T//G/+yMRWW0rm4HEGXbgXc6G8iKZnz3zsLuVj2Cks8oQaYHHC4TFOWEOxeCPe9
vjq0vxkw3XVL1rRr7l7apevz2uaof1U+YiQN1QMo39QLnPPm7SqddhcA/WWWCNmO66K5GX8Gg/Rg
8IyoEwFKS7Um4P5u6g1NX5BRUYXPJMBD17TNuwXqTltF2+A1VY0+0tqYMjS+v5cMXqcQ5tVfMnU4
E73ItGl02AC927bJaFDrnp/wlAaZZal/FAs933LrdbhCOISdKa4COhsrQplKxLm996NakEcAjO+x
be1gm3F8/mKQJetU7e/iatqlkoMWatkC53Stbm9JKUWcAdyTcXwuN/UFiha9UF9H1eqk2l16cHa1
vUnmM3FbUCRWpCM5Ct9vDgEhpIcZq6kPiiIPd6tQcv+SiQfCX9q3FdIPsz57drBP7Z7dPAi/HMkl
odj3FxAKNKFkmL2V4MpZQvzhH+rLZLF6cZZOHYyY5vgJpgqhT5Uq1XE882EHanuRy9XuGftKCkGP
/9aiu6WcvC/JP//VrVn0Mfe2ktNxZBIeIg55M4iQQbrJyMnsIheIMXW0Z4BzmF5k4SKqN2RRXFPO
hVas8WvIOQP0LlNYCdkHGcov2fpSgzXRpt+IjnwWonsimq3WnAjbQcrFj6ZNe+Y/tKwCfpwFliEW
6QWtQtoh01k0UwR5ZEGaQvt32JsBmfF4E+XYmyzn+XHmcrP70LYV1JiG9zEUg+1uEiVgwvhqTAaM
vD5TaP06Kz3hcko/7QicTwaVyMU6h4Y01hPKrlK/NNDTJ87XH25l+w0eOFJVrEO0vZH/t/0N+iIr
ApTQUPYN4g8T4rASpDAImZFyO+aZOQNBiVpBBvqbJVkpw/xp8evWNlykglh97mfA/2MJzoid+kvd
2TVYizzhfqDq2rYre15ZbRdhDmHmgnOgzahFNNz7rb9onln/KOGTKu9qRP/zqH/PuT45ccDQ6Q42
pSuPLI577JZ48Y7wJizk4djJWAI8+58vEURhMW8YR8DdsucK+NiaT8eFokvCBkJv4f9vMC5QbOYL
rljLSdbiHN4//JnnavdualuQdr3BgZKY5p8P+qzuNrD9ykNPcn6RLGj99tBk9pqGPG5hIIn3n/7K
BfmBeZQol5DoLsS84WzfR/oKqDPNWFw2b/dBuwbYQwRbmJSqXFUwXFSzBXtpUCBqulXIxZUV9X+N
ranswzNRRqYwFRoo/iji0/ByOLat71YkwCJnx73j4yjTcGdjH8XBP4SfDVrF9i3Bfc4kX36oaNeP
iObAg5ivDE9MaCq64mrAtUeZrWL+JHpETX1hWIGj9ksAD8YB5JllgDQJ+XR63zRrlpCuULEYOv7d
yPDFRLMcqmTEnV/WiXiIg5x9bz1+pcmBMssMgwtHkG1+StGbvCktbLKqz4hSWlq9pWrboJOZ8WFL
eQOjRj9kkgMo1+8Ur0+ePZzOVjBxxAET7AShk7Cm0IOXkDrTclGzC5Wec1Qb2CgV1QV4klPDU0Za
8Qr/CTF5Sw1Au0QMoiN5VT/NeiPII2sI4fyfPaVlNdI1+2BbjxrpR6oDQywbGIzDYGmWAqB9C+RZ
2KeXfILAolKgWTbanZNeNAdqNCldKHCHTIzJekXgf6fmTvj4FS5LTfUbyp5hLm+PK1kiny0mm7Fi
ddsTpa0b6ERlO15tsa5k8BqiKV8ECx7Pu5pzyRf7SI/yVz2oTxWyXVUzyNOHPycXVyB3bNOXzu6h
cArWSCBRNiS/+Ok5u4yWJ6QxOiMdeBJdvX7giAnNJoSvNm6UzMKRXgNQHwaY6HdOqMo0PgjBZ0Df
wFnJjCWO4cJkJF/zJTGYFf4dNjrIjw7c69nKoeqiaLk2iytNy1vy1kBozu64OkewdLhlVEa9U3ff
+7o068s6V9n9HciJZ22NxvxCl5BjPLHudlm1Z/otA2KRb+qK9i/NmsGBSuGcvOt6L6OiWLRMWop5
mba947qYKGSnJsQr+GffbcilSX9GT+vGQDCjY6b5OoGDcDnmYdnIQED2qc7mYxy1w+yQjqAH5+96
gJx6RYfNaeYIQSRljV/EUJNU4r39OIkkpRz2fhCo3DX/oTsk2500ncUdbeXCMgfurVGaercOF1K4
hAvLSOUca0Um4H1wWT+3HoNtUQI1sD58k8e1lWmWT934bBYifFFOysfuo7d5f56bmjzoHsaC05tF
nU7qRvpI4TFsGZnUm+yFN4CEkKDweEUs3YI38KXYl9bZtkFCVskOpEt6OqbMA3/wLHTVm/ZnYVLE
Jc5YKTmBNug3OzXDL4zFX3ad+UnxD9cb2LfWe3cap2HJ8SQ8n5eiLdJhyTSrX3QLYhgeY+AyYMU9
hoVdB2Ha35wlJB6ci2md+hvPTayiJ53bFahFE5EzHjh/dttScpLhCr0Y6be/p13NXWtEBFzot1+H
dbJvLxRGoF35caWK62tRwjmwXXTgV0puTYjBKDgenLVIGf1+Trj6Jspyi65ppWNcHLaknCHg4h7G
ydO1bQRdo0WdZ7wLXxEifR00oKyfw8BSHDQZ//6gbUPaRbfTgThg1LJZz4R+2Zc3UjnmIs7ok3SK
NUDZOYg7h4JNVXrX6nybwhGn6ImAk26178lPsxDzJEiCfmwUAeZtqRVqWtVJhCuTV0KX00gC3SX1
cACelZuLXrVdbU1ezGiU07TIBA3YFsgdeMGjZm6OUq28OYq+8aGDrP2XOAwEzxUXmbdlL1w+IEsj
2CT79Rt4u6cTTFS0p9BrNJSoOf73hmF+2v3KQ+kn4ZAKCGMKdRBGvhAvZN7Swttkutn/Fkr/t31r
gqSrbq6dnNNww8n6T5adjVxPglZc5kA7yS1j6SvFr7RQOb/0rMBZxrKM1ZZnoxCsxLtWFXNf9w5Z
zNEAG7q/CU214L2dZ3YMG15gOmgKA+Ktt/C6rqee7Httf6meNvP7XM0Y9HAKOt5Z+EhyCQYrUD/F
FCZ+EDa2GyhYGdFyXItdsRgo+85Cx30Dr59EIccCZyPnpGxnHDTCTzqIZP9/dWrSynD0kiYn9Pwd
V1BB7IH1rlcfkzz0G60y/wIIPJf+4SercH+InOG0Cc++aXigOXkpri4eyfmIA9TPKE/MBsxydJOX
MNQg3MoYn7n/SMuEAUQWQmhe65S033dNNT53RyYOcQpXDGAJv8SogxVp69LRdmGqn9Z23+tGazVj
Jvxf2LAxZBkrTRSwxJ9R2nMiMgnyOiisNQtnJn9IDgyFnQBd12XzadzZDiiPjJHmF9r9YBr7yRYw
H9crQKo4ZusxohkYwRMZjElGwHpBXALW6aifUlmdDoHBJH1Zq0VQzodntk9Sjo0skXJZCEkFaPkx
p0ABOiFheKvaLB5a0/81WDLpdrBtJZRBLwsvSqJIFmf1sTdYS90Hls2lggiy+fOlkleuVlTCS5VK
soe4rUebkW+32m8LIQIS9VeduBNZhjmNCjyaajraZl7246IoB1wkDbWkBuGC2TAkdn/iyh1R1oNs
Jlb1clvV1lzQ2MbqEUOlM39EqtMp4HW7xnNdVc3aa9lTksOgwBTk3XtdNLO6NOtd0/kcxssYLCTX
+rTr1i9ub1Sj92AnWuvSxCcdv6Ve78YExCn3/9vLn3Lw1GgFq8bDBWQnagUy7yxc9JJK5hnokb1A
6Gpv8QtDDpnlVhR9IKcOMl2BMAZsaAVnW5yC1owh8QaXAiBpi1Ww/arU5uU+5TdTynN/9QJab2UO
op6Hk4QwX9inUeNx7jeQAaHtUZsZkImXKlrcJ9DoYjd2cenUoMPrTXRJDQl0RMnv7VGZyPqkCpp7
IUvltmRo8Q3/aZ3E/gGIXg7JF0YgqtOUn+pLJRmuVQrsKW8KQW18nD7vh7vyfdG+oBMP+SlsfuAW
7Q5sGE40BE0nWJ3FQU6mtMY8aeKt2V6t+sSlpWYm+k2LgoWB+vCa/Z7TN+KrAUdiILYfOnqJ+MLV
0j3z2yzpNlL/Nb2w3OdQDFw83SSyKcwM/vrQAs3c5IK6yy+V0WdgUfcrPVWqgotxEWdjDgusyVai
jPHfNd8Up7e5bw5ozPQ2BjMIx4c8OpJ+hofyWh4MS9lKl/rChz3i6ozDtUMqhgDz/+E04tAnY1C/
YYB5Hyw4GPNzuuvBYo4+sePs0qs0BxO/9kZJACubPLV+kzKx/pG38F6bWagzskZZqal15q6n9jvN
AzoR3QXz0KIZxbUEo6djZQj92w5sINDDaFpwMYCYQb1uDRTViBOMs0fg7PVPo1EMcFvy9SL5tIxd
A+qgYEgeUpp7Rnj9vI+kgzmXxMhdcWzgChRmohkyfQuEAu1H1hFSFNoh7XGOwModVJtmbvJ40Wyi
+hQcqjksqgPJAZu1RLC9uYnhGGqR7oM5ig+Km+nZ8XKukO6tT61fZmrOJ9uVg9elKxXcfWFRjt4K
EqXAMMwrxhxOdPEcn08IYVUEMp4gMLvIiJ2n9kpqM4PYBbllRm5V9yu7PRkT/PfjtEusqSLTf4kM
IgxEGDLC4YGuW3s6JBl4cE3hKKuFzo8F3rVgoMk2uA1ZcQTE2cL5Q4RXvuqdUWCY676GDk7SRqfh
FZI/DYSqKlnngey9jVHj6VKQ7xcrOJeXE2GIZwrbNdOtDBcqZTOCdQqRxHqXWYxWFjcWA20qnr/U
ZalNXtWrpjIq6MvUntGcjgq6U1wBSe4xg5V0tO3b6mU0X1HSRDnFCNOT3KOoSGY/a+FxDeJJbXMp
oJHo8ATN1IXZgve1aGP+qAQF4jd4q7oNh3fBN4imWoByatoKtAtA17kwWyLh7MxOUDJ0R500w0nb
K18vaB3bqN+jWx7lSFkrg0W6VWXal1GOUEt1Jgk3R1kiAHhfNpQraiHLIeKnRg2DGC38MNw5Zij0
0+xOOr5Ht9JVnwkRuOtljz7w9p+PWT1AF/UP5RCy3v6gqe0TQWrBpjssw+Bsyra/f1wpDQymP0nx
lUglTEUf+iLsIH74H8PcMHBx0RqDv6Wk2HKkuwxvUIB9CfDflGnFeHfGutwm2FZNMO0JlAY2SfJK
eUTX7syw+G7XbLWyj9CgWkqcS6KTRZIXRztbsUWc+AuQfgYdY8XhzFHjIvE+kAQQ6KkWnqzefy2S
mnFVMA+V0rGCdMgBOc6eJZ/mu/3UUU6ictLNasLiAU0s31h4jQZCUhdNpUROGPnhLlq6JSMpzy2h
xwAJPNp5SvnSZk6zxySYdZTydYw2dFD6cteb1KXQreuQ0RI6bM2DdkCdWnTGOh5uPovsQL3NuzjB
PdFzFiuSThSjh4b6Piq+dDVoVYu3Wbz/JsYYbZlrPB7f7ZOOPh/5eTxxsVQgoTqqnRE+Y3uOJqd3
+Qjt13ZMMITzlr/q29RmWJiUnNVso6tg867o9qkZwmNa0PDTBToAhCQ332kjUDTXISbYBoy1PweY
tGxr1Sv37uY51zRdXUOWEPacWCfsUAh31XrRZXbCS/lZkk5vBur4o7/PZ0XozRWthyHretY7dIkN
Re7LJ8ZJiSjKviKXIL72SJyaeVTMH1Rj8nA7bvwioeMSueYObzF2uVdKYuWDMXXvpUzH8HVsQws2
wBFNgWAJzSzSH6Poavyhk7kAd1l6LDt09CvNN0zY6Qqci28TGJRwYPukcehksKgSTP42gC2r4Qvp
t8ZkkkpANRHpOf5rij63hAPQx8OXhksCmMOdAblkpL/JrJB92QYYTlsURiXCfGf202Oz46zaGcLh
tee2dIqWDTAX1gGQ3AWCWjeGhAxiBjeMoi+2snHIadOfggOwFgWbFhaaAbjxtgvNtYPvmGNqFPMD
op84w6TpfVHrSYhkNsWFdIAIZWsAugLJCJLE3r2WgHQkr5nJPPQ54LoibCtAEXVmqszgJtHkXjPd
Qw1iw94Y0/7XarTQRxRccE9cX52bDtzv0jZj917y8T8m5jOxOoFOOpV6OrjADst2FftJd+Oty1tD
xZv9EbZWgIeyju2uNKIm8mLeHxbJ7LWTd3vR6HkN+7KYP1MuBRga3Jii+IwbyMCTixMlKx1AvRKg
UZSR5hSMCl+msVOadJOWuTZIecV6o9J8JCi3ikBI4jDQrIwshQTB2fnn6x2InQ4M88l7O4Vtohh1
8a8LTa/WzU23KpZwd0GHQzcMfnXrNjdZdW4+DB0emd9EdIT0yB/CvkVTeqD/IJwyw+cJR9oZKXOi
oT0yY6RJUiRHiFUR3SxHn1sMkVBXCxbKYvqmrOv14lIzqvi5H2RoArlCuG5YbPqoR4SyZoCMVYHt
sYm+g8hZN85VOX7pnOCKc1PG7egUZZaEMCVfdXX2/Hb0ce1mPtQ3Fnid6diue5yDJQfV8uoe7VCf
JHV8OHYa9nrvShq1qEAmw4kkFaA5E8j3rWtC3tcD+IxeOXYNekl5+qhtWkzEypogKnBm7OVe2Njm
zrIM+uAn11a5BQoQp3dxT+829JQI81cMJir0EcrlRTxXByLjisaKYbCnjNvT4TQ/VGAH2adDfJac
m4Xmh0SnEXO65hC8hf5BNfpRfDEpglGGCn6ht3s8N/bvj2y0SqDE/B8he+Zp4Wnc49sVgP15+bN1
g2ma1xzs0VMfbM84R+cZwRd3JzJ0lUPs0IJQ7bhj7m7BMEM1zDNwbRuTPj2xnPI8YsDagVN3bHok
YwPJljSsN8XXSrvfMB7t1yzMsigEH2EMuBnNvAhJpig2IxYRZ3xnN/jvVMdaaZVFkUhYaC2oXymz
b0ZrlfSUmVOZ2I4sVjJNMI8XZ4pkHUsZd/rdcyH1VDP60MzevpxEZeFR8HtUxtiAuEUif7QSc8vd
Hs6QewHYkdMXxh7xh9PBEBePSohm+mxwdpLJI8GX2sJzKSM4pG6UaLyQ56cKKbQJP/BUuAD7n/Uw
G+d7Hfyd93qYc9oUWWAMRNEed6YQz2GTUd6Mvh+p38ByeYXXqwc26S6kcqynoqPhDkhI3Fd5EIdq
MAPxmSQ1Hk1oDHZyXhjQJeZWOUmwj1plCIVnancM+iTERTtVZvVjDR6PFLs5Yp42dUSB5NOWOJVk
PGfosSjsKGzqboXAm+Fxqm1Eu04UM0EW9ToFRLxH2sd4mZoAoXnzj7JrouN2aHjELTHjCSILkVAn
4JrUqh2NpEhFTrFmrRmu9cSi6iwMFwR0nmLGl63cjrqxgnjdJ+mDGkgOajitxJPSxStbKXD2waeh
1SV9kGi4iQQDL2iJEQKxatzJSGPamJ8RjpIVAfHSDNvJ/KUormpxGeo0jw4BzCnTLbEpU0ZhCFZg
3ZUEcO5s49TQDpoDtpUISFUGbP7kgQIK6n2dTK6x5m3k/d1ent7Rh41D30MkBlNopSlHmhPvnmDi
jVNNHyNmB/gE/zO3kjum68NRDI4KNz6dq49qsJVK/hH9oJ4Xl+E93Zv8u0mGjIIwI9UCJiM/i+5d
i8yjd3JguYfghXDJO6WEwwAGEpgA8t6CTolRyIFFwzm+hPZ0WiXPspU+AeM8WHdaAw0szzzPyVAL
Xk09dxFc/W8WT8h2siVlwmjEs7duR+lTRcK2N4c6vZY8IqJxatqxeHC1CQRG/kDdN+Yh6kyhF3mU
z8VJwbe6UQP+s6B08f5t77uhHrksVP77SkZkET0vJI2qUUnRhyXy6TOnXyox8ESHvzN82noDnYqB
T8nOT3sUqBcRAR188gGE+YfdriDMO6i2/nbtiu7SddgLHTJDHv+Fa0prIqgNrdcabG1ukC2q3JqX
SzamMu+pLv+fZqoaR9upIwIYXUVh6vOoLILon542Qk36R/ramIWa4/jnpdzQ4kl3EsZ4miXqYE/Y
Et9Dhc8XwAhBhcozTVqKmKtHJ+LbvO3e4EH9xX4IiFOH8fNKh406Q7ls6Fv3nf4nvr9O1g+zokHQ
PqwmgIv0aoGIPqRTvyWZ5B5Vs/dVX87bcmLeKxa2BxS5CaZoAParIk6Vu430OCfOkNEiHzLXZh7/
44UKepegwiZm8EogWEASPoqhkA1SSZ5uSa8EPwjsHN6lNonSDEHP1LtUerYoeDRRtKmx9VodUw2k
VRYP8vpwevlKl5jDzInb1wpZitV0AQlqXLvbHTe5q+KUPZhwATJXc1QHsde/4FaBGwdhE8CieOcg
NpEyFJbeua9V9inkXT6i0V1N7Mk3a+DNuN39QEqrbR4OEz9QcnPoL3ydiQ1n33QKYGGqc9ZTsEP/
TW5NhcauXnVUlaG2b2+9BbMFV9yc3rKe1kHCFo9+zaw+eWupP6S6MF5nSliopljwCGXlTTaZYymq
qtaSs3nIXq1wHtj0MGqe9C+CKJ0TU3BjDJ2o9Jlric/Mvv1LFOZIfZ3qTWzqkg2FRK0cvRWmQsW0
bTMXwhPl9aolaQCMbKAJErHH9RlhDEduWmhlmWU91G8m1SvTwVI8DD+WMxNL33mBk0KkssfgE8vM
b/Nu3TguJfarzHbg4O077tNqeGM9oZxf20dcP5SdurH7UUFJt7J28xrPnwhbPB0n39eEJPiPNDHx
Ybpuu3fsvza9GBnDItV1YsrK8M+4Ka3R41xuoXLzBWYL9NAcc7cNrkRdGKnP48U3bnBTfxQxLG0r
WVjjCAmRkMKntFMz1Iqa42pG5haN4utGjKF47OD34KoaNdzKBWvuDO7ehlQ+Y3RgQ7CDPbNtelRH
ytID86PUTFhhCtvSztInesNVDfHURcJ/bye2wQAdMISwvSkazI9+jHrB1g56XsDMwVNt1qY+r0jN
OgKtx2cPAv6q3r5e3+xiVZHkZhydpAmTGzu4lcW6Pz9feF2A0uh2jdyN+k+NZMM6W6Rr8i91Qp4u
CFm/yCcEb0ML+pHkhM4sgcOg1bmk7WrbajVXd7VGOAm/Mx3Xzdxr/WgjmyFi7vnsSXwIccgQOgT7
VOtBrk9WADuy1ciwijZewopFInz+JgKE0UuuRjgUEFiqPPyX6z0ceMnfkkcQeNCE/M+qvBIIlNnr
LkmioAos5BDG6sVtemj65tLLN2kjE5dX7OTqweEV497HPonZMrzWVSlh0S4LPvoIcDu3VeVaGx/A
vZK9eTgnwQj6FnoFVjIvsNd1RGvyXtrkjLLBDof9MtjqLbFKDSC0wOoW9Mi3ONIXVPXbZp7jIabO
c6JMyvhDr8xHLsXlU+UtCPaVirOObzAP+keF4By4JvtLnGmYOYnAZYd6sVY707g1NP/3CKGoWrdQ
IgUZ9V3PSLYYHINnGYqbgufNQy7L/8B87tNtYrwbi2U+frzakS32CubjNTG5gIjly+YbAnH6zzYn
aH+qep1qzv9NIKdv8hlypYly5ek3RD3mrhwPSI8C/t7L3sAxT3zTdsjyWmQlQem0DLiyXulUn2hF
YVFWWMKOkQJpsi0Z82bF3YrM+tmY+szZu+EOwxWVHw11l/UWhp2xtmryUCdcO74Jg3cIrTJUFWIn
MixD4/Zn8tfJVvmdjlvrdsLjD0NQ3zzh1+tejWK8U2ZWnzAINnpyFYVBTAI4WAX48blzzM2BPWWy
znxyOrTwbVaBTRB+RnAVe532Ny+UG5XYpMp6YIaJwklRkbI99LZmsTxB/UG88UI+PIWmRWYysNH0
gUNPNNhZZxQC5wRX9xdA0Rmgizuam/QsenI+DP6dwUMbfr5YZZpVp7iLRTDZIRN/2XdY5VN8vn9u
Lh5odhpD7LNlKzYEX+CXC2vdjfkUIwhaCr9hlCjYp1IqxUhtNYibFwXAfsTb5Y45M6Oe+p7ttMSH
G5SBdzrDVs9aHuTIjYP0Dd3qpk4jVsBXQnCt/GM4JSSm9O/E+0RUEX00p7JY3Wp/NYe0eI74zG10
CMK23+F5KCRtZpOf6lcgRz/AzdWhedBCf5Ki4sl19hcvhTvaCAyRUWemC8+XJwV2tzC8iwSCGTXb
J7P4FcgYS443Ua9nT06rn2Hn305xyAcISEn30/rCR/3g4Uwp5u/DvSaT9k4lj2bDaFhl/s9dOrJ5
fM+X6ChbzaTft7mzXVmdffW8R6PRyWeaZUzP2qySzXpSgAMeLaCPNlMTTdrJRhrHZ+tG/Yuthw9a
82EPU/nKdDSzSN4kJaePSSbP9H3eyg8m3ZS2hN1FbEnygiK2aKBW9eUJiMIVaKiMkfkRy9bOMp7T
IS5xFIKtq9hGZJjbvyA/b+exFzTzx+b/cIpCFvodvwwjwFQCRoH4m8uce0/J6fvLBjEvHZunLBwA
R3nKxRRQTdpaFr/eNtMcbXspj2OhkYzPhsM3/cO3WL44PcJqKCcpxN3Muq4LS2qNLCkgFgUAPBtE
y5iubiiDP2YvaExkEaSHF5vY4duGTPWbvVzDE8U8bZzyMRx70nnjLFaw53i3rjU52S6B8YRbZReo
8kOANl9t66d8ddJwCQFtnz/QdNgpuT+bRg+H7BzWhYGwTxCBSsLMML8+pqIy5PpkuwOQTtGR+4Dw
TbCPFgB5vrGBjcH+eSvSTHguXGSpkygFAgeD+m5Op/S/ZvceJ5ncjEczY3PamGhT1fXy1kErbncU
OCTM69BzVlpo8jCpaB52GvHV8Z+dGxDp9LXvDrL2Al0UMjz+fwqNL8OrO2IfVzJfSGYvoN59khhg
+xPqTyvw5ECwoMnxV8UGjQNQTnPjDVHzxcGkmaTQi21gpKqCKR9Un4nFB1n5XWwDn2CYhXi+LTi0
IqVl+0Lk317YdK76Suirqs9djhPQt9SeFhA8n+LC8y+CTUMB/UZcHoludSos6zYdWa+cyf8koW1Y
PfnVjyYjvao/5YgtT4r/fGEJ6cQcVLXeJsqNzo4i3bkEQpOmtNzeMwmhzFzX6HjxyJVko0Jy74fY
bKf/WwdxL28wuH95Rxz77HquqzSEI2ig0qq0tMWNT8+GHjlTTiZaxFvisF7l1xCjl0ABSn8ug35S
5z8ArvbfzZp+4EyozKeol830v8ICNEXaiIar25145Rd3nuzIrqInuOzY2K0D9dw9HdwHO70oFFm+
/CZPKR2tCq63qAj/hLASzEPYthfacVJwijMYcdQjVFLnMuXqVcWVhQClhbsMhncHZx6n97X+4QLb
+kS5rODGB1ZnmFrg10WxFzKEl3MNvX9Tr+owoGDBUBDOzQuKbXiJ5fCBxi7zU0SrhvNWOSwgr0cu
h9pmAIOSMsuRswvSKgfTkEtT0iXqKBb6vRqu1jNvOAs+2wrcZipAEzlQDOuFmA0Awoz0ZgpC0W2B
TK1lwXz6nJ3mXAnXbIBzoVjrv4ah+2vMIdvTRWlYCxIP1ukdAkHLvh+OBOrKiaMcFt+aFvXv/zIE
aIlxYRGG3gtg3zqjv0ymxCppURhcMgiVTiyANaAimPczA3k6kEj3+SoGhG2JzUDtHMBLu5+8ThBS
ZMMzjmk+XHWLidtqkfBRLoRQhfRb9qkz3uIpsvFayWDmSlGLOyVlTrgLLSII/4GDaz5kuXFC+gYy
+bXqqLMv5ALaITEngqwGpgOa8er450vBY0U6kZiWQWLuZLBzLdQDL++N0U3a5W+d+4yGrYGX1SzB
Aj1C2G+kNAGbILO92JuEy9YO7VAlfcc8Q78VMPAVWLLjWgexLEUMigcdqBzM5LnGs+AU/bJQFgnH
wBIKra1xCp4Uz5xs051O72oDmHvaDO4PKnOvgowEtedtVh+bd2QqS4OojvjFB8a0PxtRC4a6Y65K
5FT4hLb/NGNYWS5sxliIF0YTX4REb9w06V/a+bW5PU6/D5HQtkkq50L+/VodA2CotATchsUZEMWR
yvaLJV9Rw1vSLLmGDV6bUeK0f67hYA7f8z6BwmrZWoXU/Ijj9I3Spb7i0AVLuTamnFUECoqs6IWz
Q/UJspZJ9r6u64KT2Kw66+xx1+KFzk5XlZDlPBaDeBZ6SzONcpyNjx94b9wJH7O7qM0EPwDB8VM+
qJvQ74UWC2aDw573nl41ktpqpJFZY6I9jw/hTW6sUhFju5siKww87UA0BtynKS4Rp5b2FY7mbZF2
SEl62kd9vdbu8s5bgDYUndPBBlAjVrEx8L0EwRJaCaieGYqR3+xxcnDpIY+sB3hY6tXVvhITbaOe
KiRvyAbpDejnHrLJuxLypSppaA9QURJkRr+mlRsMaLfB8Hi/ZGAGBoGxj/vo5sqYh4C8y71bFdap
a47UdfDkRkvF7CyIX3hhbv7wbzLjmXSkPve0FTFz/R9x9a+6Wy8HzRgbLxjQvIwMZALIo4zc5qDN
m0zakr7m+XI/gqSzLIWMVa85HbZt4rP+JOPL/b44dSK7SUf5KQEpTpAdkMS1TdpIDL2qAgIPJIOn
9ngsemarxEyK5F5eBD4h8u1/+fyhiQcLYPgVzqIM4Ke/NoIarJeGIspurgNAgYwR6ohmpF/k5tBH
FdVpxZ8B37Foxra1egKYkSMEtWeDYpYi5cFcW9tevCUiqXRaD2/dCWKDZ4JiesCLHC3zZla0sla2
xfoPpuqZgPH5NWsZSDMsC+DkYM6+0UrFfHCY6SAxiT5SuJrtsnJ3D2PAzB4kA+bL9FoVv6TEeHlT
BT0Ms/ACDKocpYnGWRjpJh8wXx+dnfoftQWWC/NRBKuqTRgHfbPw9yI8AVd4nclYM0hx7Wuk8c86
mP2eG3xTDR67ZGiDIQQd/XWMyBHYg8OhplpnriEhBELgvxc4R0esaEXLMPIUiKC0YWEDo78Bwdq2
LqdImIv+f6gd5TtgrheYangWZUGSSYYEsNK+dMDs2WK/PLEergzwR+rpxrwvxqnS1Jfmbp3Woy6e
9sxD1wAwzcF5QPcR9IvEO1OXwHnFNRxJ1OV3vaPFOxR9byI06gwuvZ34D71fPtLLUP70dtRc7ACW
2W1SAqeYZYZhiaTHltPMIHc+nEUeMTUcUWtk4cZ8ngBgQRpsYhimEghpxQqQxSBNSuPx3UpMEZi5
0v8zB6NbueJ2Ubj5wc+K9NB2wDTnmGOZ5BbP8RnGryuJmIKbQdbD3BOWEuBmIXLI9Ui4o3cPbC7I
tp+FQnT+QA5t7BH5nlP2gmS3RkoZLa+YBdKYrkbsbNJyy/oFBHd+ZW+lhO1ipG8hH5O+Hgm87rsl
2S7XgQgjXExLSU4/OyjTp7LseIsnLT9Rh3s1BVAtuyph2j7rjqwGwPKcXZ1nC1VHFa992ZGz2YRL
9vtiQX20+leJeGQbpaMHirpgG6XYDLfOuEauqCKi0cn6TEc9vu2biu0ZggxODSiAyLA6nExYhtKs
n4anztkkvPemIpGjNRuqAB43ef9EnDbDEWKgtwdyuQux3MDwjy4f3ZvZxCh4c1dfuGn3OJUO/Rpg
c0PRaQnD/Zn+qJMg6C47iJoMdJnwc1yUeSBN5rLiPoVHzNdEcJzfDBiVwOM+v1N8FQI8RSF3KPPj
jrX+q0UPlxvaXiEK89cqOSv2YbQQNfLBmOjxfVmzeHAiNrdeVxB63833edT7JivSNj97M5CFK2CE
WYKwSJpgR4NoZIkADWSnY1owJyWcZq70f+JXAttYetaFdoQViHp/UF7pd3hP5YwLMFnTe0rxmtf9
X2RnLZffE3Ya6wqp6xvo3t7ap0tNSsM9fyGcn2yKjkp60QNxrHMYxx/32WMxsaWrCaQl+Eu7P4ML
QFAZpN7rmt+2NSPbW9HRkYMP5q64Ed2EK6Wjn5rKhuPV+RA+/s2+f+Bn1AHc+fUa3NLo1Xr5XFXp
bTK1aAmYT6q06YMLqiVdCsRGN6CXBfsALsaVocHtGb8Di5HEmWUOANHwh3CCxj47gpNqfze1TKzk
8ZGKiWLVIIMXg2Idxx5KinNGPTAkfTFN9KZCkASSor1IMOr6b+qjcO3B0FXCRoXf9LxxtLjQI6p8
sD5sALYFpQemiJyFOsSppRw23z8RPJsuEUK55fYpvUl2ybxNJ+UWm5cubTzMSzrSw/gE2kh0Osre
zIJjs4GGrF2F09kipop0MCTZu/Y0irmLOz7J/tq9t59pS3A0UCGsXdxsFiVCmRuciOGuSlmhIUlE
SOEXnS7oTaLJUjHbC1gpfnhrehi0wAkR5viqa25U7oW7M9m/4qaQp/y0ijetLKb5uip51Zg8iHKE
FAMlYD7FZCHjzAf5iVk7mqiBVYAN8o3M0RDgmSLXnQ/dNuVwHxXwn2PZWx7Ou+D0tJfi3NbNMB2G
/3CWTNR1g3v5UvEd6+SefGstIO7lnwo09ZNL7oizQk/7MzDCmTGZPS/TWtr+H8PgR4BBkU1cmbcE
qqg0kYANA0SBZbdF3LmYz2JWxXQOXyK7wYWjFDZRdoftJziLfHim9GeXopz2VPoEQ88J6IHUfQXu
VWhOd+ekAAvnJOmYXattQtw7w784j9Qa0A42ZDnYhVIY/NH8jfYmverZKdRcxSYD0rEJJDzmy11z
TwiX8UuTmVmN4GeuiytxZyXYHPU2WqYkZlQNm36PT7Vub0Ci7MiBos+pr44eMmg73c6CCJ+M1iZs
6oT/6b0q9nKhtW1YyXMNQN14y9nl9UbzCT6KpMNxcXw5+jq3bnI873QoEO9NJZYBuC6u50ctiJge
6f/mo5IjoGDrC4ixUfObfUi0gRPK1FJbrrvLb39ouudqEYyoObY0Q4Qsgmq7N6qFGLsL13o4GC2c
V3zcEp/Q72EhFhwf2U7J2I+QOotH+8D5bnS+hRvis7Sw5Cl9W6xNcvX8SnYVyL77lrS1RJ9K6SOB
Auj6R/QeFJuklp1gT4db3slhchNkqPSxU1xuMTUlClAt2/FIL53dZlUPuu6wr+MBU74SYu/NeKTT
xl15ZoaCNaeV2IwsU8X3xX351Ep3DHf8Y3/wtjTXdd/zbHWM2RqsAKUXyWatu76Jx+z/lZn9SkhM
sD88AO4eGD4ECgv1Ywtum50AZ5/PR+HuoPJ/d4Ky2yWV45tJiN54HZ8H8pzlsGifyq+eHXPIa6Sz
VyeAStkBvKNlKwX+igBV8YLqk1aZTELkTic+InfzN3+AB9zQh7PbU0zenuz5DUCyu88QcfJ0Ig+N
84BCAsUijyEiZmZBdw+WnOwlDK/AHCfb9Ji6YlCvUJG3sxBXkPAc1dy2VjJrz0eUnWOAoqn5g10f
WwtlVljnU42nzg8DAL020TasOgxbKiTVx501hIQgPW1M3cAnPSdbN6h1tH9HBufC+n7yI4s4K89e
fF+uvI1Eh4b57Q8aaafITPBmmOxUmKR5JW/OGlJpJpA9gGDIjgtlYjG9zejo3+36g0z1jobqEUG9
QfpL0fR/AgxHFdBXHRuwrfEGrZDR7bwCagx6OgQx6RjnScEkU4Y2bxjEx6ZBLy99DVV4LIuiOCSq
C1aDLIt6HSut7TvV1ocQgDn6cooPJDar4sAjnOwLa5phi6OsVmv40mInDlQl+IRhGztuG8XzlFhO
qqqz28+ZcAa4BXksXLEgbzsA4Hsdh17qAzyEl9dV6g7NqdGxmokEdiycxQiyFJXEbBSyv+54nKti
+ejxlzvNdb9SKDC+vT2uG82XQSeMLefVpm0b2IcyW3UpDPKCgl6xF0CoZLzTXQhmL9fBadw9lvFm
l2WqHn0EL6oWE4TUZ77MLvOCJl0tadxIVvwCF9v7ZQFt805UAOWZ2rQLmazCU4dlTX4BX/SliT4E
6ae5PBCj0FOC1FTchuLxDdv8WFg1wRz/O1TyA9pdddcSMvjai4RwSIppexS1iEQvJBfLwQ4YnxSw
GcGmnpUdue642Wj0zxsLs7nY+QBmfmyBZWL5+wqUO/vTNTMBFB5/xBMmOMvKvfMRz3pMZBj2KF0S
eOvuyK5uyu3YF/EBgBHd3pou0EuYNeuFh+YYa3O3qwkV2Zb83v2Vj6XnNTBvxTsqvV4w6nylnnPw
cXVsbIvWTwIXmlKaj360UhsvlElWBuXsFD+vI/X0EkX4ZpphLkAC+O2A7Pt9SWFGDfNFoFIaHDpA
QvPImTu7LtYAg3y8D7bt8ueI863m8o4Z8YA8p52tisYhYYa/xpNyqh3/GUfAgot1tcJDPx4ThV7W
b9Wu2q4ZGAJImXPWe69zm5RvGSwZMmWlkjW/cEJC0dVLj51E6J6EF/YtwGaZTvigUv6yYZShSEaK
oDweCCUAwZsUEr9etfFaFHETEpvLgS7ZVCuBCdBB1fzwANIcBLNHhf3vJA6EhEntjGWhsjyOo9Cg
ky1E9zzAdMOb4gsEbLxA+F75wNdUHMBZI0BbZkb+11gtwJ6i6k7KytTMfFzLgMZs2HE/svpGoew6
71+suInnlvlPydlLjoe2ANJWMd46fuOiIBbKNzM2SSvp8GOgg1jRd187W81V6pXQTnZEz3ImCuIj
J7UnWwDWYeLeBxbpe1tXeBtRIYg1YFfStjXnV3PqDHQkP8eArOqjMyNvsLepXycd9zcSMLjWQG9L
/zi34B/fNHJwKY9isLSdmpFMhmw9RbDfcO3/+KCOuWYf1Cwxd8DBjcyp5c4wEwseUfjrHUXR5QhB
TDURgceFLNu7cKUdWjFWqy04fPQqKNgcJRjm7up7ruGJ/qnn3S4fA5BwYKpABet4gz0hdOB5xBbI
Lmy7XOLWh55C4G8SrmDWGb0w5PgXzY+t3zfUnHIst2M3l7cCdkBsedfuN2fyQqDzBfGJhHKsruxB
TnLmdSa/bkEJcT90echGqp5b7ePVcHoQVjT6DGjLfDE04+k1zUAfYQsXATw1pmBPWJ8kycjNgOiU
sLPJdE6O41IqbYNpDhyp0+qBujuyS85Zl8idf2lNLa7z+aJo9EiSmPYvZ1nH06CkPaPAshMdKt1g
qy8xBpJQZjHlCrG1Yq41sLwUlrrY9ArmdNQ82T5D8xa9huHNNk6F7z/tuqt1Jp9McS8C9uwwoxT4
PU+3FsfxZPYOQDeh6o6RoleByjtbBBoqXNWY+yzPze91LgBLr2cYs05FpPhlLkf6k7y21vFdVlHx
zRugoSDeAfU2OMGNi/vQFxrbiELrsKKEnsLpdBKft5HHialkgU7xYmWw/JpRVh+gq6lXRJT3Oqv8
p380PxlLm2NRDCUmD75nrRMdqsQSrMQYYtCVheDwqgIkjmLrrX50i+wwYqMKFNChRGl0dXidQhb1
wXBw9H0D15PAb4GSoodi67BSh8YfzhJmcYp6YA8pVpCUxVVYKWrgU1gjMYNgBxbVgfFkseqKIxja
/D9SjZ1/cWy71CGklyTOuuw4ICDsfurWBEIFgZgSYDsZszSObz20JhamzqJXWTprWbeDPum+1BdX
7+zBCKv2P5naCQpsKm9G3PAzhHE1AoNhGDkmWRlk3eck6/2RkzTMR4kHzYw0uKK1bjTPPe2k8+g/
8rsvSAptL4OPZ04nQ3zh8PpMi4dR0zX+0TL9Ru0XHHbAfqsKs3EdLaXdAIAKDweC6d03OrVZzAY+
b5t0wHBFsHwigKoP35tQgVj5PbKIJUPMjCUZKQHBe4JcmXpMXqbPBDohx/tClOfvkXPkzxn3lxev
SKnse5+2nk39ublHKO1ZXn3lyV/dkVeSgD5IsCep7PvAwvpMIqVOQfehZOHKn4UbZi7do2UO3Hmu
wDJgF0C9G9s09u2HOudE1CGHna5Vnh58eE7rV6hF2rFWTkbzDF+livCRA/2wJDuc5vjLFL7YhFET
rg/QbwrnJVkEXDwUZ0ocQI7UZgdKJj2erIhRAgiE+7XyZ8zv3g70ZJW4K5zwRr0NtzEk/vKkcybH
/RQHp2tOvckJNuhpep14ajspdT/ygvYkv51joGcbn2oNy0bowPCC5E469oU6yNVSUbGFrnwYwGyq
CMlqcdd32C6awyZHshacmL9B4XxkChjcwzhHUfofLwe0L5G0QFNVnx4EiLLblsKFXcs0Ln0MyMZR
CDIQwK9F58D5JHCTibl/waRyMLpJNj5EpzMBiKJ2RKCTabge8851gFZ7LXpq8/vkJ/utAnrPenEe
+CHIN+GKid1Eh4YEgzVnZg38eOx88G3yCGL2H++2fpW0Qdv2VUMyApJ6q8gv4rpoXpVR/dNpIdVG
KKID9NavZII9U4j/8ldVHEB5M0stxyqnSzPAtYkOmZ2YfSGJEDuTcWRIdVexz/ZJW6hYvecXSUiY
kOJVXv20+L1Ywp/86MkPfoMQR8IkNRNuyLbGO5ZJymMyrN8zt8DpeITgr4Lpk7LViYgzfsictAR9
fb6b0y7IS4iuQ4rXaM1FloJfuB757KqDBm7GAktnQuPSM12fdB9OqnjUofwmmnCHFy5pX8jOV4cC
iPYc9+vv+mj6qxN+Sy6f7yzRPuGca/BXpzwRZHghdTXzOlcyTPqCrRu/gSHdZ9vpdduRKmxtsuIi
FAai5MW73zC9CwgcsKGCzh19J/19k6KoGSGDrjHZTARu9iuU0P9+3UuksQcdqGl4i5FQoJzNNCaU
CYxWTat2iObg3m84aqJGwVbjjpjAqUV3lZXmYDx685/Zp1ycrdxdbkHrVZIhAJQny4pS0DWPzSPQ
xLIc1qZQLLqXoNnWowLswbImNCLbdBbmcfrKAxH6nn/v9g3FvsyzVmZM/I6wDXQdJ7AvGUZR1QJx
YA1joRLNh56pf1Xp5eB6z+9JNBhGsis/Y8ZNBpM02MA3SFeCExlg5ebN+Ce8JEeAj/Cd2M3YsQTF
th5KVh3KdS/xfTXWGDD9HFrMTGZvn6OFvc3z3VSgoG17DBl8C81WGIijPeFlYAGD9dOixQUEQwN8
3WxxliuVtjBoPUqUtRf9GDvbj2rzwZyCaasVtYyX6HQ4uPhy2oeq/ca0R3lXAwFDFwzJnMfn4mPM
+2artPk8/h7yragbcW143J7S/f2laNCwNCIlmhQqrhiqdE6JQn62oy2JIlpLO+VJv6MScONqS0vd
OPFPrC/AGYEEkO7B2yYUDjLYNZp8w/TIMxobmHP7RpWmzIPW/WHC7agAdYA9VC9CgyxrT6/5UHeE
T1fA9eFNMJ283x+QBIsgmpK0DyPWguWN4eQQBE7j8W1lNglEVEN2qqGte/1rF6fLXPOqzEpR8y7i
i8NA6siWBMsiJUBcMgFfa4c4T5MeksqUS1MIxUaF7b0/yY30qS9HxmlyXOHmxAWYALi0j29GPtIV
dXXvEDVKhlanSGI/qDqo441chmC/uH2oaxn5S5+v7rMzmXgJJGhN1D3VrxvwqSZ+70UJY3gKFvHH
xEJUgbghow/U7ijOVzuUAM3RV4GMHWXjUBCBoFR7ULwjng6eOlaZDHo6tro2IDOktPwnZn7qfQx/
DT/7TMIHDb9LireX+MSzQ7dOlRmV1IgKHM1vQgJOtGn3YpjgJwOCtznLP1wBPiDSiDeQPVM3z/YU
mwLz6k4adrR53FfvjGnf97Gujgg9O7qUm+EJEQAsDDAk5bA/rZJVhcSW+AFr4vj5OuDN/k9OCZhB
hQAX2eV20CAPXT287n77SQIbGamDF2laz+BU4mtNhDC8ffIfc8D4N0fr4jmkU+4nsZzo2bLruGI9
E6ct5YgVwfK673b982goEqkOl1N/rAlADuMu3s6h/Vh8L2z3j8tjg4iUlzN04SJVou+fXFRnHrif
eSZW4frKAun+W/xi0eML8YR+sRuaHrpNHq+d3vysJXaFt0SaxHfNnfSBFmLXcIgVnVFU0bTA/y+t
8VtqQgwDnyLgsoHzSYXLP41K84fM3JkA9w8VOm3PU9zpb6fcPJMdyw514iVcNnVVSUZdeuDJeyYh
kvi+neK5zrxihThrgU0cTTkXic3ohYhRsbgmnntsWECmaf4pmaW27HiRe8Wt67jGOtl9RuMxF/kE
agSniw9+lBkgzXvZUUU90Ck4zf2Kn/A6WTyrUf9q7td/mnEo7LH4llwL9blsfZLJ/7OJWmCidlIP
rJfzr4QFiKj5oIhn3BFBEu63rlN7Kh2e4j+dRIUDiyzbqIgPNPjhTtVPKCzwwOgzKCnIYE4H7OvC
clYMC20bRG0BKya8bkfV1CLqyCWl9Jt8GEeRx/oEjVFZGyDviE+K3b4rK84OoxXPagBfqp4DW4nw
nyTNN1mTQfHciUMNoQQANSTiBUMMW98XY3358LR39kdfAG9/E12NAZnqBvMf+75XvB9c6pZoUzzh
t2oBM5zFYYPOvSEGmGawrpxnp7yN2MnxCxz3zZelhS1LUJr22HyrJKTUskKq8BrD8E7OzI5Ik6qJ
POB+O1wXfgqdOUFnT4tHs7abslgEmrGmX12PUaK1+HokU7m4dNiswUHn4uyYTsmIWRh6iajH76yW
89wwO1mwmWPSs4srG8+s9mtUOK4fKICzMqbx9IPo0+s2OTZp2po0U+1bORRqdLgzEF2JzzGdmUgc
/gEJd2R9Ph7EmXPgkNt9PyON+dE9ZPiJ1ChPnJUaKk7OTTswGtq4FG71eDLWuUYHhpGkdSuDr8NL
ZZXzMxEx93pOhtymr3yK20hfcc7h5paXMv9M7oAscCPU/Fp8Jc3HZkLeAJIsQ6FfaqlgjI2Gjmlj
ZWuyKdxGKvoNc2yacCM1eOx1akAKXKvwgS0TEEjjZzdfxo3XJWmfF/zUUTmx4sEeJIBqU0TerTJY
y8CWKfNMePeYbJohlwe73uP6Opu28fzyrb98ThUKt0JmAJK02/JsDaTo/9jIOGmN0dCKo6SeykBZ
7uWRjC6ChlP0tqqJTvfwQbY9AhfSCmvnzlxg15tf6j5VG/y+m4/zPv0xP75pfChli3abABwBWEKJ
mCeywerQSP1gjf4umNbWMt2mth9RsZj2FS5tK/lL4JtxHAzDggp0G7YUk9y7TDPhcayW9+QzVF0H
ZspwOX3HpxcnEWHnuK62G/wobQizvT7I+WYttqbXLOVMVI+8/zc/abvJJ/+CjGsNtCfn0W+naVY7
TehZD5cqD/3stnPI422R5ErE40VCtVdGuul+P4Z3hh6CouV1Y37PaLCG6npMwzGkCvSXxjdyxFi8
7c0jTTprXMwdhUcIY/v7lYE6d3zG5FXzTe67XylswPOQI1XhCOKegLWyWv/Ij98bHAcRmq1F+47B
NzXyl/Qs7rM1GOOM1L3Qy3gBz1jEfvKdWHdiyx/ZtIDz0PAQy0fychIjyOute/DAdy4WvwiXi01b
PhPWJe83SFbBICtCH5lPVoFNqFucJemHXIdV1wTRDqy5OLPY5++7GOBaRwiD750Vbk/Im39qSlfv
QetL1KTZCaDzSn2icGW+nj9mbaJl88yBKrRXThCKzinGsx/ABEqo6Yi4nER1M9JAULgUTLmI+PjE
GweHtJ5pG+utO90bck1kzv6plGg7Cli06EtXjS7FWM80+8unfcupWpdUZl0gxUUXiS506vm6sWAY
1k0FKE3NSFRKiSNuTlQ+qq1xwolJ128OEu6swel4RA5W+zOlLMGa8v4eXghfOMZ8sjB3gDCRBXyv
/7drYsWYXOeDYRml4gUZZB67aZnSoZDQLWwIPGHpTUvFGhsXFzpf0ZL/iE/t1MC4sSN5ZEgBtzkF
DLgDPdzzeBrwi9tmpMgHQwt2MtYGpSEy/xFUqZivbDa4TzQcMsNF4XkP7DcwfdduVV1WI5+Iobps
ZLVAGqcbYtrD9k7cJEUcm86vC7cfa3rDxyovTSMKpdENpZlx34zxhI8ykDUSCm7F7XL0PzJmTlE8
QLshVSNVkcVR8l7DEWBxQgn6V/6IxoNk7on3Z/2eI/irqoQUAZI5kA+VopB2gjjjkurwiIUoIsBv
Ui7jlEXSMPstzKemJb6A/hT41sMp3S147VBCDfjr/j2UknEfLkH7k+waw4ByhCoGZ/tC0Esy/fDB
LcTCBpFNl418amzGwKreoXUgAeZjvba/p1mfksNAAmURapPSI1LqDUvOA98MWsQW6p5MDy5WkQcZ
FdTJSjj0Dj224giXt3Nr6AZ9GrkuWVz7EMhnIAZYD8ZmbyqFvMl0GWsZ9jTz0DIXtLp21SK+uuil
QbgwotUieqUdLude9EyPa5uMhFYiIGetCh6eLhlm+doMeqpLFq2drTYxrAVnqJDtPELCiOG9BVLc
RULHUHRnOGcHpo7RqJBMofUKbLs5it97ARAbyAxiiK2g19L6okQZNDMS9Zufx3kXcR7PN/DVU/Cv
/UQXUXytFNf/ecO3BkURIJFrMfAWcyeXeOdWLg4uFuEiaWFJk9F1W6HbTuvGvuGE/dxN8AhxDb3F
JgnS1paDTL6OpiQBIVdaNboIar+kJSBRd/mhiERFqNQUpKnC/2bup4Ifg2eW2JuyZwQhq60KNZLb
G8wQp3BzcsQnn6OCZRdpGrAscncly31Bp5Hm2UxOpIZdmEFF2pM3Q5jJ+iR8ZJijGuT3dzBiOJua
y2o2TNY8VJZPIiNbsbtb4PGqAjBkbajpJz09WMqE41WVLTRFFuMrTqQorq429v5h2pqpnUXJ230z
WhkhOVCCEtMdBCVdS/L1CUAU9h9ZdgEkt9LCVlln3Q6TY6oAwhkq9juBLqtUEdGSnVsyhq2APIYv
Z4sF+MNiUNyHPqGpHQhf1EY+WaKoRTnCM2w+Q1Kud1uFtB5gUYFluAQHNII2wr4kUKzqAS5eRvZU
HtmmRuDxFGnV6zcj1ouGjdAwBdDsu335NGCninojpy39S4LWtzUgXYPF/c25Dhmx1j7dM09S+XjX
m6kXUfpltIdaM9OfveQNNThAEeW6rPK3ecI6G5wsgKbyoAp4Q/Z0gK4HKHcHMRZ533bBLEHCwpYr
ruTRMFii6OM3tjj95Ny/x8TMYODU2hZwXcTsPillFfmIhbliqtWF/xEyQGTrOXcRdp0P2AWkylDf
NILsxSgHe0j8TsqY8dTaSMo2P0jFbvwVcmpHCKk2tUzN204raP/hdVzmIIwGPCmQRDiaagdPMSPA
mUOQsOTebXRddyrhltt9zxPxI4zcIX/5w2yQDr+ScNdaVGo61qsxnxa+nt/byx/RRNVvOVWqngrz
uTvP1OSt3cVgqP3rZcRM7rQni624nwND0msu7peyhXP0j0+XVbZ8bCY/APYQ6/C0y37pqXZtsisf
6lIX8bnleX5mNZReR17qxIg3MsJoQd1Vhi5ozPjfr4BZHGUCSOPNNULLtj1+/VmVhRit8wuEuac+
0bZsSCIK/yEdL+bS2Gvkad5yjB1hzvhpoRRo/OpBYNmBMoXUwK2j+QXefkEp7dsGIjkzYtmNTvy9
xlCJJM/PWkp7AxLFyE9fHVibjI2t8ayv2pRl0AoKzEz2I4e0cI3n9bghwGucuqe/Rhs0RkaMiHwN
AUWsKEImiky8oeSjuh6JqkCo1gYrPnGqQVdOiUjb0MOczoWjiatHdDPRw83WYLVvBahZSxjvgr9E
WVqRba2xwYf/SZ0X6XzdQVT8rXDf0w4b99lirkqpiQ2vDoJ5MwqrFOvMwn+oPELjUYTPNEOs0BcX
wMq9EVsI6jvvWw73pOSWthScEq9Vv8pYalVgXoIPUXOC6uYMEv1GXdg5epo1yCdoPLRG0/7ixGqj
O35e4KE4/oX9nGgWu1pUbNRf9HdBJpoqDZZrEHOfzS2qIbQ2kgWhAIKKK3OBvSmRi04Gjl3aUMqA
0ld1CuKA//6gj/LZ7NjXT/CaObi+9MvhmWKcL7skoK5BQOtcjJTPRLZ4GBk64oPJLxrdqkaweoPC
ihjiI5kPe/qevEeqx/D2XybeLg87wkiP9jfab2SZIPD1cwm/3fkgGCMQBKUclqHpOWorkka64Qjq
pPngA8rfquSosTY4ydfVItocWL5W3n8Sut4xobj/4VvL04MdLk84uGa7OwrXoB4u8eOfGppPrsnv
hrX209GMkSETAnBucrDkQYHMFphbjQa2grYH7O/M9cmjvejD6ExMttSbzB8OIUUFDM72PSTIzspa
QsHcQmdC91HXVd0PEga/ZAK41sRRRyYrHLp5nD6F2CCF6sp4XHHE//3ZdUzz4mN3W4BmKiKp2/u2
axPKBoN3UxIPBCNFno+wRYirZMPo6+RN+DZbTNbZE3UEJj6ovVTNLE68eBAjOFwIf3yCfKKe90lX
R890QJKiNvNtuzqzoBfIF4ZOBxj+MlnjyqZFO/MedSkXpzffD6H8FLZOBbJGFQwbzJBhpZd0WBon
FpRRyCIi2mQ/hl4loQTmBTSSILcj1+5iE/b7iiJ+XdA/dXnhJJlDX/5yWVeBhJJ/CJf/6vWGZNQi
Ml2TN+YqQAPW8GN85SeuNuzsMiectJnOJqznVT9a14jS1IXi95UWGM+C1coC3evcMJY0sG6cPlZ8
kTmaUxQCBRtfICIyNyG8N+z6mVJaFogoBbXpozjGAyMnm25vPfElDaX1p55D1Gl7ybB+0eGYcYaR
ZGnHg+9rqSR0CYJ89kVMUz0KDJjN7hDDGNJZupVQtv0gpZJDvFUmBliySmqtN5P6YnUYuutd9oKh
Acr0wr4bQsD58gosXDzpHodhg0Q9M5Iva/QwODvvfUIw3zlis5JOYwIbM1vI0A32kuNJpARml0A+
6+pSmvjYECtx9VHpCkCl5chu56ztrbFOHKuVAjit9GoYQa/512JsN3uswdaTKCbtCZTuPZ7hIoP3
Drawh2y+9WJFHi8uXzKsVuwVCK2Tdz8PFMXTPPSRfw6tdW3neJeJZuetNlgM7oktKoSonjepxTA4
lLefQ+4jWyR5hv9aynFKtHI+lJc4yMakI7iK5NCf86a6sVY7ReTKvg5aZhcCyruuLeG8562W/PdU
GHgmzhSq5kkKWcu3MOK3qxm2tMNY2PgszqdER2emtM9yded+/lJI//OOs1TLeN4/lxCFnATqSpcK
i+XfIyZDFtoerNWmd3CTfuRq46KiERASpe0HMU9eJkKVUlpHqmFDay0Z4a9HMT3Vp3cnGD//n2RQ
VgZL2QruG/wDmgy4PtYNOp1QxY9iP7Hb74Y5x6rx2r6raO5dWMAggpveOaoJWlBzSlOTF86JYVJ+
D9ANxGYBFN7yK4dPWmOgKrBY6vdDm8VNJRl5vwyCf5vHu3WKv0suEZPWdvDpQN9KVUAl7ZDh7cR6
Hp1qkYMv8iq5dHa5LZJZ9K3j9DV/JOisAtgDJPlWAx/WQFierwbymJGuOePL3wYlOgbW10J6TP0+
PyUFB3LeOn4zktukTUndx6rEOvlBINY9Uin+gWPd8mRJEu945OwL1MQXjAhfYqkAk6u2ibi1dJv6
7c8glesx9BVitGloWD/JOO2GRe8d5W6kLi13EdSRQP4knCX/IACQNZvCa+IjbpV8qGAgdNRQzrAV
/d9r3GImkD3dtlypR4XiSVeFCeTe38RyzR8s+xfFOMC5OU5LiDiLW6UE1CYg/jFXDjx0oFxE3Y+K
IiIHPOQHVU0tjf3LbuZMrteoh4w7N5ukRK89bHNCxpctSYGnmsL73JDv3KTUUMbELzIwb6Q9/5QX
JrcxT93sZrS48j/E3/6Y9nFIT90WN4MVLQgTcTXAumlU5Jo4yYe9cEy8uUquCo2Mc+GKPPaF+3T+
XgqacPB98hcDvpmLZb4BDnKPUM/JFnUiP/hbwLrGJe8xsKNG0PRU+znFGZ2g+9t+2iDiblXvU9I0
zSwPS6CdfilptDPjo1YLpqR1KVuK2pc/PihSmGCFtgQEqhtbtGgczh2yIXztxnh0VT+gvyDW7rr5
Rm2qbrokoJAQh6IRQfQwqKcQhIZy3/pVII/SoOUAhVbHsCxvrJCoa8wAW5PyQcfT26IDlJSOKfuy
KhQ1hAXj54QVq21c8B3NdjzCGn42a8CIDB0T3/lUzuZklXHgPlRZ/As3Ax3Hg2PvYd7po7+2Q/WJ
wu7tk5L0c4o6qmzSti+MWMR4cckl8y2mfIbrf2yRIp60UzhDMBGfU88DJR+k5dqVKjtHypL5ECPW
gUaUNRgaFppO5dud7yQ7V5loPphv9+gz1qckHxjS4X2f+Eu+oUFIyUGLUasbM6ZWSQu2mZ8IG5qs
EJbN6XJuLLfDu0IPS3Eh6chKIwT0OBV840iQLIjJAuweM4L9D9b6f2c4BtdyQVmAQ0zgdGmeBvDr
9J2z3ZcrZZRsYjOVdneSNHPkOfjLHm+SFvJzVeM5yqmARV6ztSdU4Zvwhp2svQ36LQBXXrZ1AL9X
D9dkJa4MQzFZHTdq/EjxQsIt2O9a4ZQUFVq9kj0GRgTX9X9yvq82SYJSeslWxVqouu5Cse229a5N
oZqzXX6pgxTHIFCmf7aZ+sqwUVfiaxIvAvYwdZBrxW+eGhikgjvTAH6pXD5aQwFbcaTJI2CaBePB
g1DUgeWK4rRj/5eaBnuV+7ay72KpgTcNvZfttaNkK08LYaof7bJGah1nvDzQoTuDcuEeroS6/Rvw
FireSr8wliP+4o2OZpxX5vKO/LbmowJ/J8DZfPQ++WmKwLEz98tlcKPlOcCGxkk2H1mnywzUp275
b6X5ZLY5CvrhBAmgRBDIy6c3BE3fIrSzJfK/zXyz28S3psWvTFlgR/8eit/sNwuOut0AXljsg2UI
6/XOGZC9RTIWIUB5TMfxtvcdqUuBMMCtgs19fBAyAmJGjVKbhWEi21x5n3b/kprIheoLo/YSMnl8
QVIQRUiQgv288kLmrAHsZ8aLqak4CWbvldqIdjgC80VpJmngSMMlJWteths51G+yi5ZAi0KJKzC9
3sVUaAKsarNrYgl5ADoVMjXCHTPLcmzSH6NjxlIpsRt9onfMDdgEAOC/Mcrgj/OMGoXCWuq6gjOX
7Jif2XOeYf+sTLzvW66A7KlK+hRnQSUCAPhuQ8KYnDcwSxT0ENcJz4JUgpwVN8XqTwEedHjgcepv
oO1MoKsmwtwLB8z4+4bU+DUSKWiwuOzTNRVFvSR8oFzG+1ZyGtOtDmLzPDtG0c/bAb/Ryp9lme85
2qr5A6J+xgFlHrxsx3lZk/kR4bXLWAYeIQzvTBHm1o5N7A7ibPZSeNSHe9rXYM8XAvdZIbOYPG8L
/X6JB7vz8madrlw7jbOqnPq7PpqdXxuEXKermeNTf5d+ylDt32//n4AMgi/tAzMGbjkVU5OM4yf6
tUSmnr0Px4A+fnrVeimqMOscLtewLQcxOumKdXomPWbIFqv82/f0KxpTcn0HwBD7B0aFJGBwLUkG
0u8+Wb07BG8dXhScpPWua5cPgspZMeONJc+9D5BPoCRQSGNvHBGkDfiXcdusvI32WAnayCT9dV3o
c5bPgH9xYnQf6uWsXCfR52W+P98baGV+qKqAIyOWDgZLaE+LX7cq8f9yHxcNiXdlnLuYZxhD5F1l
KPio98//bQeGAaxPbJTbWVvTeCj7MR28uqouuBe7dAZKOadLfSSPP/ZGTF6TxEvFpsuS/VsozI+s
8y+XZqy9JAA7m+jF7dfaZpcul9JmXoNrkqrM6yDXJGoRaBeZSWJuYyKywMFDRTPpOLYIOZPhv7Mv
UkIqeWpnSEAr/fDO+sLWUC4P0WhHBBJrvwEdR9GFXmpYi/0GxIvO/F7b16sRYinuG6JS5FJi8IMx
52ml76T93i7893xx+9lyGXlaDoo2rAxFyewLKbmlw4sAlaUYz9mo7GlFmVCBye0QYHa/POJXWt4U
YlQ4YlM51Oo2T4BTZMHGHgrBa+Iyw4aRdgVAyYJAM2YNRpWo+Jktcq6YjU8LHuiX+6IAgS5N4doK
erF+qbYMxTnysk37+S7L0i+0KYwVh2i1Pe90VVRXelCE3+qoYumTVaHv4od+EkmeIlqVKb9AlCtA
IGYNUBP9NayOKuAq5qjg8ZnDtBzK7AKBUu6VkgnXPjqMFHaYNoN1hWh4iHByg9fIZcokvRMBawZj
vamVo3PJu+skUmyZU0GUoqchSZnviXgXiRouOHXCCQcJU4LLP68BYjpo/fEZt0Fgcq9MfkOSGfhN
VSOs2ds9tRT9krnDoOKP0jOTRggwrakxsSzQxs8tsu7YIFzP0f23HIXv5mvgNSkGsxD65YUQJyHM
ORO+02L8KJgbHkAuGVL0xYj1aSP9KUosWF274fQTOfBqqseiUlWCceqzN6Tx1/UfP2Vsgn2mgav1
3vk5U906qtPOUKf+1+EAphz8Lrq6tvGrn4j65g0JrIAMAiHul2PbfiBewolCJM47l7Yt61ElGvZx
bkNL11mx1jMC7PdcyQ0LylbQdUmOPUTFsBzpG6zms2as//++NldjHlGFF5iFibVSxD81XHda/GoB
E5U7k5rNkGvWxVShuC3y/MK+vhzHCI5fhV0+6OLInzJxhMJEgO7Qxpvj6AZs9zxFkl1hPE3bFI1X
6Ilq+Wc07A+K/lEfO35ZILzeA4EmO4jnhbIUutQ3ZpBqkayBGv78es0VI6rY20/RosyNAwxaAlUY
kamvS5PqTqaYhSQsUbXDeU17DXUqM8V8BFqrte15SAQe3uhWVO7UBJM8ivbdiF3AFcvFnsVAPr24
FqINhz7/NsJOv40jeXanmBn3Xyej6GoyeEgbQkOn/uMuwNBhzDJcOGGVB5ofDO2TdM5yhxtHAXRo
Iz5WjDSvSMXOOdXf4fsbku3bfLqkWo3AoXRg/K2+1paLorXsVTSksOetHABCh+8oNZL4dx0nUa18
0QWret0nhzpOmQpA645+A1SKkfujwpF+q1oOM9jtNMZXtw+ei8ztNZyk6Qk5orQEd7Q+0qfUtBMJ
sB5TRetmp7L7heBZC8YLnN+Inn6HslWBwZcm3EC9KrGR3sco1X7M7X7kDDpjpwWn+K38ymkvVAKn
6C0TdWSmiisuv08WtbFDBNnTVWU6sTHPbGkG/wrLBd4ep8Fh9LPUFWz2kDXOGN8RZagaFhvWsMN+
YZ4nkKMXNlyIsNKzhN+Vac56rzvIMn9bsJSkW3nqj7P5hq4R7MKxd+KBWP4Xr5xQxqiLX5szbaeV
bqfecd6DC7/zzK6wuVMmKZg81XGY4phG+Wjhyxk/VbFiTCjjibBI77epDfO3gQrNAz6nDCuiRQeE
KME2D3t+xFY67YxX6LwntzlgtT/mTTuTwrStFN4v4wl5vdSIb07Elkba0i68t4kPs8ye7F0Mvb+L
5QEWEEZCRABjot4TBy6jNqXtoBMrDT04im24CJ4jzSf+/DdcSYRXxNw2Huoz4thElgGQOVwBuDj7
kNvaULgmsFcSoci0qMWd4Mn30HH0VsZlrfCQ1xb7VbsJaPE/CaLAIjWUETXAyKBXIL4YqbT/kZaF
fg8VYGNjCMFj9+zRPglv/sxR4VZm4NEhAhlio+/xAwxWbHc4yGHk8+T2BlSmfZUZvmZalYq1ylS7
A2BOdhytE7jIZqx6qgssrP4LvdiEUEeyaH0/+X1rchiRWnucB2oM+s1DzMgHbwHhdetUVTxaqgm9
MKQCs9XxBfy5LO6FKJFvcmqoMBNfa+yInXE+J2mgWQ5bBX+XqJ0Da166gi2ZT2l1tCyiAmuDW12L
21nLLjwil5lPnx8glHU2wgXsGSwm29DwW/H9XOPIeN6IY/2f+KpoF4qu/qHrezFkxsHVKPW1kZPr
CGGBOtwW/Mh/UP8PUh5kgfgoZNt753SV8rC3BwEnVst9lqTMXbag3xIBA0/FCKgWflSIrCSgF2qN
b4vhzoiXdHe3B1ErS7WJG/xf5e1cAJhX4lNFA7Q66RZx1sa0y2g+2bGPOhzLMuPqqp+HYjS3+G8x
hZ4lW7RXZmuy0K6LDbAXVmMzM+e8+8w2IDTm8E1/TQKiSqC3PQpIrlbooxMyLs1tCt3OuziRYosj
lxd6t4pr327I8zHypN7xuYcOC144BrXhC6z9kC+ZAeIIaV2hqBpCb895gw2kJ/xEwbKbCzEmwigc
KY6dmEEIfIVxrDehhERm+o1+F9QIs9k4GztJ/mUERr5cCOGE0UsY7aq1V75thwlKTZZXQzZB+/q4
Pt3wkeVeMhxMg/EiczyjDNLnUsbfuCe+85JBYhdKaHUBhTop7Jqojba6gNmlu5a7FQhuAB5fAjRW
u3gk76mVWE1rDHhmyQ3fmSUzG0JEwdwUC9NTcTnIPlOvVhFThMOv3vNgJY8nd9ql+iPiI6utirF7
u0QJktf81lJYj24qqv0j+7yQ4F8lld8nEtapaq/f1RBO5TwMLKktpCgVGyjBhfzzsm1XwgPKRcxI
d0duaIcDL7vmeww4bETt6qtpS4B9p6MyeYNL4C0fnzfhmS00UFrFjw+f6G17mnVA+4aKeB+wEzCm
x5F7dgKwbJHq4bjeD4JXXsoDEnVjeB2BWN1SpfV/xhsM4brZrPyqgiO7aFz/o1gWUFw4r4fbvzy5
3xvVSzCRdpKpXZG3xvCt8xmQn8I5oqNJDRAH+5VUjQGMa/isJ+rBfAOca0D/rQmyEUQSFk9NOTsw
OEN5yzI+ikHgCM8eaxkgVDuXOm7gbJZD+jVoi2QbRu3imB9tiJBjCgucin9oK9OWgaDB4wpAOYzk
jVPnhrjNTpYh0olRtJls2S5Q0DEjjQyOvj0b2rfmc85b9nxS70JSxUMEARxKPWeXjoFrVrMlC+Ze
v49wO94/Lh/RL4Vm3arwwqGsnN+PzMaGT//vdS1Pg998cjs0Xd6cqwHpYGwEOvhMfZqxgqfWRUDo
LwBCJqFGlfzOJ+N3mq7fcCJwem34+EJql7F8Oz7YvCUWxXxaJbP3HFFRXwIstvCJK2dUf+wHd9H8
+q63mRMPdIRsJitnNPARyImIxMa2r+I3JQJdTXxPcxLI3vJr8lVKlJ0gg7z4mevnGnj7mcrVat7F
M4c+A0ntRJ6yRvykOAPR47XkY588paxxq0oP1ws1LU2Ew9M6oAFP+qRSL39eRymeKr9MAbNYYx8Y
fxPy6GBb6Vl294Bw11u0cUHtCr2D6QgrxBF2WB5xNMXJ7YSRS20mz28FCFTtNR0bGBWVUMmS5YWQ
U/oXIMrfk7HT9JqOrPJuHEa6T1ABEtDILdSNxVOomcF1O+mHQzDakz8PuVXs87jEvFEWllto+vrW
GZix6iB54lGlqHPsE/WF/KzRWnSaE0eFN4rkQobXpZh5YgFNEKsDlMbQT/MePRyZIOes0gN60b4Y
amP4ujP6A5lioDx1VK+mPjmZmTl0bKhIz/QroBju9S0lyta+aG2z4jKTEJsnJVLHKxXpOqxl//7C
4B2npjx2W5Le0IWas43biovYUxhpDTKROI6BRAUtyrgke1yhEdaro9+Ebsq62dNb0R92U4brv0XT
g8BjAbdxpNtoAe0C+GpqTDHfHFJW25WVyK/82sUPktvK0k6I4bo8Wb5j9P6P6/aW6xXnYJRjK2L5
oQxjk/U92aKCL8oGHh/k8wkDjUexOe5d1D9dJdOKCtHxb3XF4/2/vkP29aepWyoG0L6l2Tt5Czzt
cOFdVWl7WIK02gIYiQo4ATQz41CO+MWscKQAzWGHwrp6kEavT3ILGb85GC1eehulWEFeAPV5hYXz
AIz/yrXgi3r4Ov5oGKHjCPpjMNyBt3yxgSX7Eu9LJi/+Ew4WxZ9D4qA3jupnVxwDgJ/PH7UTgHjm
DKB8Hs78F+Bgyr0RGvj3ynV64dCWCp3bxBM4h2QSbPuUEeJ0MmANU7H/YbC10foNF3pjiVclsYDK
es8X3JuGJo9SBFVZiedYaOljuOo+43CVmMSQCyyk7wgJ+EIWlSBZSwI35CEr872VRzbLAMv271Fc
weiVN6m6gbZnz1JyBZifTntImM+gHnReXXU4pHRtpjCo7ZkEuMfy+XOeCHnzEdEoT5WWLhp1N0zY
M41+Vn/QHEUmqnpz/YqMWuLkAH8E0JHT1LM1E1efzMiVdGxi8OD5xugzMzk6iwvEzJlEfYVM6Aes
mrINiok8wBTNsJ/bPG4FQ5tuZ7GKU12Z0qzDR2Zwsss0mGuAI+jK6pdOvvKZw5+ISwp3LQD1Usnu
fJjscQHhfmAnoal0cCBWzwgNlBzRY2gSJXL5X2LTWXT5ejEOZv6LwdX34WYjIEErItirorFzwaWQ
6er3XGlYNGoVB1G8jZiiuRqhDF/DX6WYsRl1ZbSo15fZvSzwasGkx+3Q6+P0FPekcV7n7MmX0iP4
xN8XTQ/dRpKHkgH7SI3TlkKIOGqexOOYd74J3Yx6wuT0dg6+9pfEDKwNdyVj0wIoDSBgXLi3cdVO
bcgyyXbXVYrRXUNeaZMz4w4DyQNQXNaxTrJgR/4mmr7A2B5L/fZAri0nDtXXh9rzD2+1yVtENaB5
8szKdGQuhL98DMz2TUq9eBV4duI4fMb5nfHMz64b4MjcART4iVRLjw0SEOW6rmkaDAmrDh5DpsOR
R5t8ZJ5SGUv+zRzBy2zQXfPbv8zECTlNOY8HguLQy0yHf6wi6V/mCKrLA311WYoYmt5CQ6sDGr4T
xngP1uO3+QMXZ/11e6EpbX00FdpsCyWS+/PXM3zRf8iUNejQB71/4uNhcKz6eVzyfR3qHn2bXlc1
oJKsj34T/NFWz0gfOEDw4Xu8sIspIOoY4g60wLzptv9200GZv9C2oBqK7kif4d0nJRN2tLKm9YE5
igLDV6IlSUG5C5HfBrwjvwwgqUWA3U15PsjK0AeyLY9KumMqZwYufk0Q/LWeBksIFrccJv6B00jD
W1oDP61LBqKcsY8iTEh53ETRfoiNdTVT8ntqVUdBDPBWb16gbtRGskHybeCHU18skTK9ZDKUnfyS
gZpZ6kfhdFSkchntfHWgMKjaHxBhnOHTJn8zhRsgz8UvPJLeSpOd3orEWjFFy3Xn2lbGjjfdm9d7
pm6L0nDmmKFEYyJitFzfeZ4nQHwcHOg0aYdvSLEUhHEQMvDaPNlEjfSFebMqoHW5Uw244HtK4er+
HeptfiT13fGMIHrNZ/I4oDOGkNbZ7Cbs/gSoCj/xWjP3GPX6q3Lt0mKNxY1O7NBHzUEbnD7BFTqY
4G5wz9XGcU2R//U2hdXtKH1PuMbpTeak7AFrUj3+Z++A4RHBQVIpPF6cHWsRVbuk83MDnpq6U8UR
eqiZLIDYHzAyFJAzLTZhVLPPa7IkWKgP22yeYX1APUKzj6p3w/fY1KooGXfveDcCS/u9S/F4vLl7
pryjT5gJTFjxTc/3HlZSiedeZW9tBE6g6To1mz1fiMbW+VPqxgYheRtRA27VYa7proD/tDYzpsWP
pQ5Df4Dt74fm6V1J5nFvMxFuzCdDVwbRugdTDd5fiGKtQT3DnfZyR7OVNTKMNN4X11dOTBT3T3Ji
AGgtQMx81EGiYOy4ZroCVxymqzyEKfMzHSP+mQivB/x+bSBKqSKBfJLX+vAnyvf1zBjRc+AzMrLZ
AUZGykigTQdTJf8WTUOmeeUun8biPNZZGZaD/JR33DukpiASlSrkg0WUDbrisUD1524KZwxB4Ren
6yNuQRA+2Q7sxxX8LYfnEJbqa/1a8MnY57YlFWb65XV748Mv/tSIoUA68ngyUyodZ+rR9QQT5HVm
WekuQhtoknTR2KJtR589g50hjnJOIputmnFNWs3WXuAC5lYwQDIjIWqoFoLkeDp0JGks6q6+DY88
AAhUZMS+s0FLl8SITTbbWK7ruHnh8pgVUoKojxkJhlp1r7x37TZIT6182SdLXdx/8qSlFm2N6yH5
2w+KFxPla/X+DG8p5c0r3+fZAT79NP/scJ5LMX1pb3o9mjZW8V5CoQJLkgdZ52+CceWFqi9Xl8uH
QFKB833mSWczfJlWSlUvAWF/Q1zfMtg6VDMeRmR7J/7jZtPoEZnutuSeemvpjGcVVLT8glVTsrLf
7aZgNJbJ2cXOQwB9yc2WpeVZGE5XBsDvO44wRlOvtx8BC2l/kcGs6L77ePckjZ6gDhAjtqW8O7IN
VfWzCWJ1q29CQ0CF84aEAGjLkjw/tio4sFn817+c3XGFbk2ElJQ1nEow/ppxSd0iB9SKwVwkAdLV
dtew7aIjagw03BdBLD4d6OeozoC78fr3zFhRbNijw2c09tyxvQvJQq7LqXNBEuO6Mc4U/sN1s/rC
VOQCkZIaWRLN2kdQPLU2sDsHpWc3LkduNFm0vP6vo1X3NQP4pm1lcX62WTY/2jXBDOlX+LDqt8SN
09VWib9wGOChwktJseHoN51FUl5v83/xhfyIY3/KXrFUFHL9RijbW9XIMVG/LAGZdv81/1Xz9+SU
TFKtEoiQRHNLGGv4iRB22KrmnoGaCzET+rfP2Mro38iX/9WeYSXNIeEqhr6Q++ihSsXCBc2wxJxs
a2/Hadzrfn9Q1UFN5Ur+Buj6TQ5FQAEjuVzDvfi/iy2Ky2paJUFiswdeWIPfNoOPOJqbW7zyWOGC
6Du7GgP3lVxAmebLoxqjFfFzboydB468lBgithUfAryh5Oyymg358H3Xf7BOzFOfaVmWWjdj+Vug
kot/YSjz6sDm24Q4Mdq0vCK7LCA17HHWhclcBuTR2qOXnsbHTuXTHJm+g5T4U05bRbsotp4dgzmx
xyUFicr0MqtWyjjLonppuVi+e2gktCB5/8hAf9Qw1u8tGgnTVXuZlRoxvNaf7x7Mx7izBLIei/Ib
MZmE3U+eJjsF4vgbj4oL0pBbVCmNGphJfQNgqn/NN25RvPMZWtzZhnTLweBlnAs9ke7iLUbeC5VV
OEZZEpq91htxH5/gJRzZOnpyR1TCntAVB9yzhILBw+TviPfi8/Yc8QId+rqlQkGAZukA7L0eUq+x
HVAVCjYxteahl3aUW4z7r7PNXbewJVBve8cokPR28y3z3fOpbthIWQrhTXXHKFjXfKaMoqhDglgv
xwM/J14fbtp9WCz8Mqp5IkmRe34qg5/1Y7wFWwaBnhKXZOqvvgizkGjI7HCLst6WK4pWfEcjSaP9
JiImXcOsN5+K3losKY8A2kpDm9fAol5y4zH5QOqIoz9rgDKQzF4U/VxqXdWYUNxV8Bv7dvMYUvub
uVMSmDQaLfYr9qACg/6Hc8hCfpj1BEALgwmrc7YjmYL1cdIXNX8k0icW098z0ScSChIjQNIkEYUY
8sx0fwfhY+9DhUwe4uoCFIK+mAo9q98F8gXcMs9QdR06G735tULqVzl3y7sGC02Z7+GRv03/TDsR
FmqgqzU7z9IV9JHIO+gYPawV3E1yQidRbCBpW0eOKHDK7jqujIfhwh6Hs8es879tWSOvhhJKsBM+
HkwQn9T/o6U/kF1gGdbOoWZdeTL+ls0cZO5XeXUt5HmEUvHiNMXBg9Wg+Dcb64nEetYp9JAqjIYd
6cCapVtCSr1Dfuy71PjqBD7M2YunY+ZEgDMIeiDO9X2QwyCSj2i7CKIgYL1IgRV/+GN/ZptLMWww
QALsJdvMXS2cR6kHaIOkMxrw37ugyQwZqAlTYTmXv5Vcwdd2vCRnEchJGE4zZWbFnlZvkY5Kiv5b
c/VKxyoir+KSSzYAPjHQ6fkKZXy/gfSD68OCM8bJFJ3LcmUDfgZhjxwjwUYH3yJxDwS75fXrd61i
Pk+Ugg1ELiTaAffTzUUBTvygSGFe6gE2nBQoUnOJoNthzvk/IyNxXXYnmVlGB5xwnxCtLFcerZPb
tlVde35c4DxdMURQeChvNVU4cKO0May179/mXoYHDdpc0+N4lJXtsw3+l+SZt+mQe0ALkGuW5GoG
Ch6zYSCuD84XdVck05hQXh3zDq+Eyc8LJXylm34/jm81cmdmL1oVO93Q4uZPUOvPR5+QBYGsuYbe
lfj94lmp14QWxDceYPrRRjOkzsy83TfaBAxr02HxYfGUi3ZLpK4aibwyGMKj7BcEcm6+izZJlr1u
mpYcV1V2mQ2sBExTEcXdXNG/7O+CYpJfgJheyogQtjJOMZG/N4jpKVXwuE2WPsaKSGsqLijlxxTc
GGCDQX3ju/jXP912+4c56jhyQ600DiprLAllqieAtGezYd7GMdqtd6+E9FMPYmhNnoSx9hLPWtsx
uJYvn7VGbHkcTVX4j2sbPMpHhr7bNezfmwJfNyjsap/6v4C7o7E75NfVRN8B/TKp8MTSwGNvuaKG
N3K5+449Jtj1sU24Ui3r8NtEnM387b4es2Eqv4HBOJ6uxPb/VcvfcTGFwPli9HE68y84eOfJaAwj
b+sFLHNJveYCWdWEQdcgz0KnBYVn29p70eSNsrLOocEgLbvdV3iQlLYtoUdpUT1eR5WMKmrbI+3u
DsR6kT0tqWTG9lK/8OewDDPO0EFPieNGAQy32dOXfTyZ1QXt11Yf8neqbZ9F4965IuwejGYt6AWe
nulJXIbJmGIVq66ZEFu9o5edlp0ynlWH7vLuliPBsGMpPrdXyJxMY4SjldBBntxofF0k9/XOfoM9
RVwfDiFdQW7iqj5JWTs/GeBrBR48068E+OzKmDqmVk1xsiE5qr9nAKKe80EezEe6RDLtMggufDrM
ssq/Vb9eVR7Mrn+xFH9GZYdeC5Fu3RBd7Fyd8x+SZ3eQuuQ4JcqBNQDj4+QwJD1P2IlOiuSGNiCO
v7z1lIJdEwbwV+o30ZrIld/A43Lin2eHO83kcag4e+ASlZnX47h0yvByLsNVPf6i6BlGuAEERtAA
1Uz+BbjAHBdmfa0DYjYoKJRPFPftKtsonndEJVQQizlKYTZ+JOTKMJQw4oUczqlDzQ5Z77u9HxtH
IzvQ8yZ9ImwcvJ0IsNKwagBzwkMI593yRc9oSgorNYnP89RGw+fsHvqpweIBx+oZvkteFSbTUO1J
NCJ5tNNC8L3KIaQDP9VsUjy/Ilf7OkGMR/JKFT1sSnPxXuwTIzCoQFiYml0YvbzRwMtu8LyWRObz
WqUchJWitE/8cJoiVtdNlih/QffLTYZrcYdZ9cxBuIZ5SDxBgLwoktZk20nUeK8dM0vx76FKlFw8
mqIs0fadGTp2ook3T/VgUv2LHKRcIBnIhkCF1iUgKjRd61SS0meW+9J1O/+/+sI3Cd8TB2e5p3Sa
YnlW/1CTd/GesCLI4QppuK8bs6NjIlSxibEGu+0u7iMrexcoWi5KzqhwWPDbex/lX9iE3iUMgaWU
+QiHas0cm5jChOQ8ccAjxo76zK0R0lNzQEbWu0/JsBVqEBu770SlWKpHv2aYIc99IxS8AqMpLtJm
zePVEYfHfLEXO7Zxl0vV2jRwARy6giQvJzbnPQCQmRyzkzOCJGl8rNabrljr+ECyPhfcvrjOG+ZW
VICPbTtGVmKPRx/POuKUzpKyU2vxdBGkKU8cRoTRgZ8/hw0jLFz1d5hytR8K7fbNYgBH76Nzpv3T
OA6gi3M+LrtgET5ByhHBCbx+syCUfhr8GGzstUSqVNiTBTceXCKvmsRkVvjKGX2igJ11Ji5da5nj
OAyP1TCb+fVXqIpeC6gIYMysOGCdyGd24aMTwfGj2/PLCabc7fW+4pSvSo/EmbMqFI46DxD8V03b
JBFnBEiMfH1QNVo+HD37Y6Ey7h9CIVlgDESe9G9fiPLDXQb12T5876tlq8mo5CuuFAV+nBezNVxd
nPJeDP0f728Af6pFObtbqd6V+6uWeiCVwxwFoZB0NlO309OzXBhrhmG2+J53jgOxsrjpt8WAwAF2
eoUU/1NPvPrUesTq7u41AON5IvXTlSOSXYGHCYB+/yVYVjBDZwfiJ3Lx7b3UNWYWVEry5IYZUsyY
F6jWiqaWjRVPgGhl1TFP/dx34ZG0DsKX0wbi0tRQZ3IGjoYEX0jYaL8eKc6+BLYobXqtotMVPIo6
ua37f7m9OXOjg5s92Cx1gALBArxD0NYXLyqaAn9GnYlvxMZAaCEoG27qRU6x9wWIv2lhX6YQ4pta
V1w2qQZsMmenVjI2TpK9vlyzrvS5hmq6U4ikFVRltrnqfUcWt2V1KGlFgiWdSmRqhCF1MfVm5ZD7
cYhomm/fjqxEwhAB7oxAsMHQi5S58P1sje/ZYiKc/4hWSBYmntctop80iJFW1aeA1VM6M0GjPIak
XLFx3TxjIIzHB7q7ccjSnA3XBx6Bdwsb+FBTh8eTIVyW33jS9Do5mypKe3CrqqMyLEThSV3PZRHE
nfBbQuuEBStL94i1TP4I3HMm8Oc5I3lmeJOpRT/k+E0uFpXqWGJjNyzUnbLEUJrYvjoewKfjUj2Z
i/aflqLZgcpOdpsT1Nl8xROK1DZFzYaR4j68LQFomjlZHRFkEDxhf5WxEB3rD3dcUVbr9SUQrY45
4cPuz8tr0JJ7Kw4o8QdvUquc4jIamtm9wBebVGGytVIPUmzDQszGt7b2q1KdFJYapQW+UT2QM42+
qWI4C53epU54mFyQboWYxPqlls4IIHxbAGUnfanarz9B2KSNbpkwCp7hWnKPjLWW8MqPjZoBic2D
otH06+b3yzxO1vAHrHV7GAX9Q5DCf/qFbIdJE3cwi+HkhT613Gzu8cN0N0lLzIlQv7FDANBbVGBs
sBxBMVFRMo49juKWoIyXwhxn63LTmGYufjUq0cCJCLcKjsqzA5RmMpNElKNmIDupbbO9bjA37SQN
xP9v99zqvdAYWzTZPH122qMt22RpRwzthhtu8XTls5B6UTBQBjaP3QVUpwUD57Su9U8OZgr3+per
bt26tgLbuOwVu2APSKxavvUuGVs3Ym08rWUr5GBUYT5wi+acX9Wg+/NXXErfvo4Y0SvY5R1UfDb8
i6aNGDCWLnx9GIc5sGVrRwfe90VH5yD/A5vbkNaHZlGsG6RPnVAko8ZtQhqFn8vD60wRrx/sx/nQ
MsAUcz/DNeo/AJcAIFzQZygqBkXG69St7G0l2dJWPIf5f9hTprEra/iin77f3QO3bKxITesXuhvi
BSPDhBdM8JcNsOiTrYdyhFDsfbCD7kOtEwFqg2xE2iRxh8BVxjZNNXoN8NgfmADaI1Qnxt8Vu04K
qM73Artjm4VT0Mc3qZTFKhic1yx87yJUat0jd5obbLOoOuEDUR+ev6dPNJoKh5rHOKaKMmv9QDyy
MBreuki7B8jdrTnpo3Ug3eUJZi8Mjn2KYZtv86WBPWXtDm0rZ96ddmUrL0xVyAU+GpKw8sjnjyn/
Bs8zfeKsbO5ixplRM04mC90nY7ilK+EwPK201HZ8HIPnodOmyeI/kayz5P5yGuniC2Jc+EIoElAr
5MwU87goZuWCRHJhK3pBj96OsnTzfZbm9NXji8TXB/vGFqJW8Prk7Mt1gqxIb/iIrsvbuhD/FOGY
aW1T+oxD8/8+HNUBn9SJCH/dq5lGaZUVpsHS3+pAYCahMzRkfTu1z44sIrltpHuaDtxLMmhZVXl9
ycZ0fkqhTmroLiiV04oAzXtVu2TwMxf6yAmCUWzWlIrRdZ7dArnneEMuZ1PrfmKoYHv7w9vPDshN
7FewDs9OqYfqDA1ehx5owYi94QqMhyQL6+wkQMzGLj4Dd+9asD1yBAjkhlQQM7DGblt2EEDYnYSA
28YAgLbIf4FWzJIUoZwKphOVxoCC5HRlT+w2pd9EgFtlaBwVi0Dj10eiFla+rr+6IUDZhckGfCiv
TM4YNIWdSyBAzkIujLliSf9rA2eLZJnJZci+sEw35/fLputRFNd5kg+gEnblBZP8xZ9iuv/qAq6V
6OoOGXOhFc3GXFJBbsQYKwuhCibh39lU0bM5N4iocto7RjbOl53niR1JmCketIKB32yKGAFV7whQ
BuLoptzmiPEI1hwne0l6kwtY4F3/Gzhn6LuzpzGbejz1Qf1lN9IiwMaFbsoWueTgiCc+H3MwInFX
h7T8ZHSQadznH36UbB9nBZJWLy2fcGfEsB6QA1Nf5GmOfCYjNqOoOoS8dg9I0vTsWaY+zsLJOu33
ZNYFr8+9qoQULg4lHj40L8/Y6Wma1uXnfTD6a8EqNqoSmezGGPCC7nI/lf8Xy7229JJEr8zszhsx
QDn24HVcpcYpSwYJFsBrEU/+svCDVVEo+l5XIadBPepbgskYlVHAm985VODBlTTHjnhSVy6Tx2lj
orKFRO5KMUMrtsRzeOl7Ej++T3XiBaWn5zW+4feTexBs3q/JEG8ouPFxrcPbtqgMOZ6LJOkNTOAw
dWZeBbb81n1AT73n/g3BT8nOlnUxxiRk2KM382HIS1AY1ksKg8UXMy+WEWwA5JhNIVb8uNp6e/P8
6QHXOQszGitKLPAh6mLcP7M2EdKu9AGKc8Ih9UMOHl/f1PCX5Qr3mUEOzJunG4/60Ff3yOCgPx1p
q+KcfCNfb+IW77ZFbOoavIuV3aJs9HuLI6g9RbIjNRNlUCY/GwdzMPQlCVEH7ZqNuRcTIrPePeZk
Qs7tej+OQusC3jE42OGX1JJcSjeVtjdAdD9o+enWZqHksb2W67LgC3x8NMyRHzc7yP4u9oU4Rocs
PU11r43RBsny+pPwu5gEBy8jxvbx+k9ViddaUPZGXX8CK+rGte/k/nox8afd4m+orH4qmOKqCNny
ewCMRfqxmb0kAzz6ObkZav2FGoapQAcB+8s4CfGuCGOJVnvlhpvtSm+sY2rHzclZ8mCDBWwXBlsw
yAlNLMlIMr1nNSxSevdPGCv+g++73dDpmfulETAL7xht70h+G3y5dp3F171gs24byVWxfiMEmR7F
ivM6LRAWsj3FKsXK7v9hFG1udfe98zuArrCML/FSV8ScxRqHMnebBIxmtDNU4kBOGsf7X2uKOGbc
4LuacHaAL2lsaUppnlx+uwIjuIwdP2jmau+UAxbXnDWq3SJKIRfOvOM1kxA4Hy/SfEwP9Qxbp+w4
muPT8uEUeXj4FhQjAWWRs9vDryvUSFvcNeO0/Vx8MG3L1kSA5BNLcszRRbg/fvNn1QJ7qSSepzqk
jFOPKhXkEsAKUME8YsuhHjJSxxGZWb/idvqAFtOlCGDwy/qbDqtGfGWCP4J9CMbgmIlB//CBmAPL
brzXa9qsb9ObuhpYv37wWDsGxM1oI0f2uMuchGE9CnIirKNgIQYdZu7JZ3me921DCZIz+6msTmQY
xnE1np8bUXE14OiMQPYI/i9pngoHogJ8++432ZzULwOXoFRudiFP2vBcm78hHeXwVYJ0xOJN8Omu
U38kBK6HgySdwmdNI35ejhTHP0wzvnlqZx/ladbCfQMwgTR4OVn6uOxIHos3DtW4COD1n1MDAWQp
8qtlq4bXG6QHz1r/+zmckJIV86/nYhcQCUPyRLBhPr+347JqzEBTp3C2h1p1+tfEsnkOXVwZJXj2
nq0XOflVMDmqB+Pbw+DKKSmOoDqyG2F7gySe4fJE7komt7ri0ALl+OzqYPsUU2C9Lj01W/scpUbr
GGEI5PcbaI5VBzil/4MnWRnVk2V0Z+7j3a5zrNc+SZF6vrqiGwl5fBF3wHDsckAGXzGFM6OgLLNI
7w9QMIUrzyaVFJc50NrrHOPL/E8xMypTXu5fNuy9Pl/ssOtgIoBg8xeyzZ5Q5QSZsOJ+71MimXsJ
+Vy+P0u/bqd0S7+0OB0WZfiyGZ84bcs5fg0LlTmHUrY3aHBmdNNtOdm7kCj8AGI0X2N5x9Qc2v0K
pvmuSablavCV/PB3n/Z4CICCCETBjbp728YNiwNcE3ndlyQ2lQI5lAr+L3t93xzg7hVULh/iLYu5
7gKuY4zDb2M7pc6PTGtxUyniiiC8ZiOJKEocku3+WSv7JemJlIy+OSpzeJFrW3xb+Anf3OhC2SFX
uXN9NKyUYhksBrioEZNof3H0LuD+VGinw3jYaNHeadeEUDvJVs1caySsgXE/ThiA+9nTQEMVGs34
l+jmyCrwW2e4WT51YEq5d0rH5YRFB7vdLFim2VlNWanZswD1+eW1FBIVD/Dakgu7MHhhenHjXq6n
vRU1QDCR/65SN3CbNt+m9yYIgSzJfqzLlcbu3TiO22LfFm7ZMweR1Ki5wyj+zJ+6dLYx366CrSEM
GuwTkTu/48S8ZhRXDvTnSJq7F2a3hGBdq0+1s+GR8/4uIUb6Wow99ewNo82sKeXkFU+u40VawpTm
e3FDBy6Y/rlLlhrb3hm8VAWV/ffNmGYPrVBM2lanT2d4k7fYZ9ASCVymZvVeP8ngmf+EGUn62Ojn
192T+oS6B1dGet2RCF+pSaAom0ecwNV3jGmFsexI5MKw1eWbL7wLTwk9K3lJVWfxM2kwYdBGnYt4
rWnSzNw1LVNVPUVXzuLw4UXrQwX/LYyn17NW01blkl2IXCg5ipoO4S4aV/G/oBjYEyJxLb/qwUmf
5vxvUs69NQ8jfHdHUjcGYkSPswqd30dawKJnMg4ryk1vjlXVy4G2iTp4DMEOEHoUrGQX7/SZNBgo
1Uu+phPwhi59MdyliUFNtKXiZIL0jr31xCzyuOF8LZXpPIjsRL1Quqw4xWXFyVInuFlYdulJ9TJM
IgUJl1sxU09kceuzoDNkMNleVnmvs0aBtD3Vnj6a7fdRDuFQLv1SXZ4C4cI5Rk7Tdt9j/uFBcD0S
pW8o19uO+lEM9UY9q/VaqYSKCG1QQgK5/bIwIZvF/mj2Sr91GfgpjTG+dC6kUd3Xlr6ktEZ/vi8W
mdwc1zbEeMMSzrTNIFqH8YAilIdvKyVAyOr7UMDOUskaWO+yEsysdwSLIZZ6ZzspSZQbrLWafDIP
rcggtzq4lVMSw3963dnSS4RclRpdsX3gPb47GO13DBb7lPXr5QRt6Gkf2DKt6vqaOC4aIt/R4VJQ
O6ZOuSUo5hKunmw2bPyzy7VbDYIrmMUK7b1vSnO50Q6o3aYMu0CcHhkEqBFS4fVpPrhy/Rtl7/o/
oXhiFpFSu/UmA+PHS64dRFhT3kaGceihfnonKhUSwk6rvLGd3dhSsKXIFwulvzro0FzZMGATS9rj
f6O/YVuwTYM2HC2fgziG5VEiEbHbVRjRXI0wxIKi/4TFtxrbfuwaLkLKNRu0GVx/2jX5DRv2kdFN
wrK83+E34fJEwRDHDe9g1U4QubH29/1QrJQTZWvNTfAup1SXcXQRr6oNGuJNsQi12MfCoxmYxYkX
V4iEJ7gWAsRjypeSelvCuyv84I2OFAxODY+tOCtCvSeLODwOeMkbrq39CdlnfGORIF8HxJgOOHxO
etnP5nD6wPZ9+lgdEmd86oOJpcsX3+IJWuqqJ0s7ooiMrsUz6bfcWHmFss0iE+G1dviNDNEfSH+b
hDNi77MpHwMfEvOe3tgwcrT6dH8vI7ZWFj75cawnJ2jIijjO0Q8BcdGnp7+oTAu4STtFdsAxp+YA
2VPucK+bZQOTFKI04wLoOUNeRhvTWcTnh6GJKO0XLU/yhatQSOC+1ix9OxHpUYDVExQiWwJpBjT8
7lf3OQKs5t7x5dAj+kyl/KnV6XkRfghhCorcn3ZWskQhZDgAhluLLOGtZvQxqs4y552vfzZwrT11
sa6eBaiG4XWcm8STkBM+ZZWYScQNdUd3EVOkSQ95NtXYjVsbkQE/lukD6XSAr1Fpxn7qdtjKAGJ3
L7ifoGSQWEFARliMZx1Ry+kh0iMYvQcNKk+m4B9h/MD0kDCPbhN5gELuLvP5JW9D29rS8b3MHIZ2
MmZRSdbbNRVFLo1Vif8+ybaJMdb2RfQNSXHz3ENN5T7dCi15OsHzkluk1mOqMM0BRFzOJoTrq2hq
ZrTqcaXZ5aW/Rlv/2rNPFrlZLtSzxNFGDYbRaxuYaloMMWg7dvsZmKTsSAzUqncWJUov4vQDzai+
m5oW+5mSorU+Z1x2uElEcsQoGTF+iabCBSeF1OUEOXhbKwKV5z1M9JqTUPeFiE3nax3AgVexCsEF
80cqgirP3ZgHeRM/Hf2He7oRmp97Xs3867H/mTkLKYyX+ZCkmdvzRRVBL27njVqSF4tmLc1dvMy+
7pE8In1TFpvaaJ9idhFA0DaH9il7xSz7vJrX8ktLgFQgSLDgjmC4uquUlK7GjDjlb94rjN+YX1Ui
ZG9vkjjO/Icnr74niFpPa+7fxw80e8cnp5kTk3a/i/awzlT4TFEYc+tn18sqdAtFqgb+HEMB6Ib9
/dK0Ldco8yv+PPC7juF5nLyRAwOrcw6VuawlTbiIqWOZDC1bUDrYV48xyxGFq3x9U5PfLvzgD9hz
qXG5D4Na649iDtkPdQYBY+D4uRQHjyqDlsi4jceid8AZR+V7q/G0jjcYu9iJNO7iCyg7BRnV968s
EMkH0LVroEWAOgOeEDpJISYdBPN5K++745mPsTStlEXavmeGqrRAb24peqq7i6lG9AAgiLRN6Q4y
8n9lfC68rlDXzbef2OOxTdHfeYhDVzB2oVavkf6pY9sUAMaPg0ZOskg1u6cnTgFTb0gcMEpMVIR7
uWDO0lpUEOrZ12/0h4/GnbYn5V0WAIsi+MGh8lflsbUoCXKhhG4yz/KcpcCuHdPp4XhPIRO51rWH
8wf6lLlfWqjD2DRM4WIsHgVr8HTmx8FPRzofSqY7Ku0o/ZB2QaXdoRZJOWU7AjWCQVHkEJ7V2Y3S
GBlRlQbtTwsJcm1Mc/oTby+cvw0lLticTwsTB53Vpy+euVp9yBSqf+8DXemQx8AnIEBsZI2f3Vt8
SGEF/DkmC/B+ces11/p0q5xFv2O+kKsFcQGWYxVeI6SsiABBpKFKKqRmV0RiowMyvI7CoXU+j4JD
2RKp/QMYgH6owE4Yt/eMgo3NyOEb/3AW3qG1nME0O2CMOYHpXZ13DyDD/riAbiHD1fWnWzwBeNo3
D2unN0PtZBD6WLs7PBv9885AMrRWqXPLiLBuE3pxp1w4Pio80ox2BAVhrZD7xQL+mRtzftmcLZp8
N0T0vj9SgZdykKJkpJDltKb8DToIy6G1XneRzpz/j+UAhh+agJSMGpVlT/eumC9okbn4txIqcqbs
nPc2+OyLWYuNKsa8LBKkaSOyISKKsG0dEIPWi0DxtBp+BhrTgUoq6QqzottRoxjRtkCNEDSfeOfD
LAy3NxZ7xQaPRCeXQP5IGiggodjCXSeNX3G59ozRSPoG62jruU9aCkZN9vP8CkaV4fxvj8fCOq1i
xkiCKazkwt2ZSvTiCcMlt4xu2ya0Vzzuljqy04/b5grfink/60TecG4qOdti7qc1pfFHPluiV5zb
CzqsCs2WyhnwPqUJa9faaTqWxoOYOOkmsyKBVEkygi8Ig35VwjNFQGhYyK25QvXnPXFewXW/cVGQ
9WF63bRyMdFH/0DeQswszMCBGjDt0LAwxX4H62tBO43F36FgZamz64tHc/XODRqjnAMaZZZY1HA0
LLy8BVSSA4KBBPervybBEu1Lg0Ww5HK8WlDOhc6Bu2e2/S0grzMXgTdP/tyXb/uTVPmHYSNThSKS
ZqcxEaP8UThlBueKmgmjFvxkopaa59CU7pHV081SZftMW/sQAJU5nTz5iLXeCvvLnbE/In6cuyxY
henaltox0EPINX42+m8e7flNG4+AScG7fEh9eHFTwuVzvYEcr7N7/KstasfFnqvBi0JTLJY76t2p
fSijwCv/u/J/q5s8/+wBY16VSbxzEkDoaO+SQIMJHuTPFbHlFQKbgMkUvN3JE5Zkk7i2IHkDSMou
w4d1CnqQyZSTmCYNsU9SqDM4JkedN/0DhUTpTULWuOHzVkl6sq42Z0JYBdfeCK/Oflrt6RAudr3P
H3gY7b2cYsm7smKEvcjKA6ibfFOaDITgnhyq7VbyxXGT+O5WBI1FYEPBrAQ3U5cEPuagZhDXOKRb
PUdGUrNCTBnejkuRF9bEl9umIoFr5cM8jPUcCL3mvaHJEXYo7XyQKnaib1Evw5Q5zt7Yv7q22T9m
Crr4I1JcesICiGkmmUtOj0w90Sw49qG90rXLVg+03mHoiYSLE8dM86pcsCoQ6lKW7XKCz5tfmj/J
hOcfLSNqmnKknFpNS2ZSgEe9FBtKlMwhrAO5MKL6TMF3Grpz7N93uGykr1cAEensdRjdSxQ1fl+Y
9Ud7MNLzvL/KZZH2F/bS2+8wXDY7otuEOKwlQjvRUKcKEDYRomzKyfDt4xnr6BSUyolML95PyAk6
BP6aRJ8bNanHvmCdJl2aN4KMJlPTQuSnoxvfxJpR7O9/PTyJhtu4K9YzD8ajLRtm02nfwJ8tmwIj
HKU2DCj9+n0Irga8GpGkK4VIoc3+h5P0F3lA5E7a0a6BwBhdaiaOTb/NeagKJOuICigGLt3KfEbq
TbbI0xrFYV/OJVXy5IZxNs+R4RQYMe6ImRGiksjP4Mk4/39B23Q/3cbhGDp0f1lESDUFoyOF0rEU
NT1Cy8QTmyVmb/RCY4zirkINuEN3oplVDcfr82d7uizUcH0yhJcdpMuR+4gHS4ba9R5CakZOuCLT
jDWrI6wTvviOI8dUA5oTOoWnA/j2RF5p6KZWIfcxDnmVMxuOQ7IfjDqEKnAGCbcd/erXHc6yj+ER
27A39PKV29OdYhVqffV07LX6cB55uNZBd3DS+pi5g+cyV0Z6PsWHJ0hR2ioFfAap1JVmNTJlsyFV
Mt1a6wJE5Ax9OMOtHT1KVVr4dntY84k9B4wxIT9xN5D2ejaxZKZX6rgNZf4eGWyeHJtCGImod4BA
CnR0V5nDio+nCkubgqaZM0MMmHoBGuDJRy24KPE3cwofy50Hx5Xg6ecWPeJUQe0Wa1lDdc2HIZVu
7cIwzuMo8kI1ZIBHY1xxPUNu+CUR+vayz1IoctciBo1dlT90UXvxXAareQyunXFlgreef6BRBBbd
Edvauf+1qFBwU9dms9FIkfo+cZ52mIjLRY3N2d5qw8Zi7Dg4EXjDjwanQw0FvZ+gdySaL/uYZgT3
mJ70QxIZrOvqQnEkW8sAUHnMlHx/RWGkYcBOW0stpi+OGxzzj5Z+09p2hrLEhFXjWUPZEvDG1yJN
DHNXNU7UMvNEOeQj2DyZLc8N/eNQn4gm0kMcaVUmIlaErWTu4Kmj+6noWYfC0LBlqERej1Ho92rN
IMTyao+vtdoUv4QVYWe4ZBK3zCPc7iiHJlcwUq/0DxTtLVb8Fdtib1GjP/agDzKuDQaXXq28flC/
Z6mGDcDnzE3PxHbOH3t1Kc+VmxbbfcZVKJyM6LLxSZFiLNi+FTwbtyJSmDZ/JL9yza+dlSG3iOsI
HC3hVsENSLLPLD1PW36s1wQUDVHSYjP1F6NVUNT21+/RZFxPJ6/BrPV2y+BFHlscFV1zhKEbXCBN
imIVqE+kdVtfTxChzlJ0G7PclN3FsS4HiRwzzhATXMUd3CEzQlxaVFFHda1KVxKWiwLP2BbRzbZI
PVWOjgosRXYTP/qhtUNpj3wFq4Enl8qel62Me+dbNH245W/t57F731u9mgXxqtrydpMxgKk78+qP
rNpvR01gLtxtRJrvq1H8dU3hvV+xbv93hIRzMGNQc3xr/79qIVBJPxaQMiLRp0Wdxg1Uy4qm6brK
xgqDrKH+rokZ7CJa9K2sd3PD2HPEfFnxL2DNdnNq28XxvMP9OVxEJembeo5mqeVJon0fdjeJcms1
/a+zsoqQptTnft4kiU/BGpJ/stWpccOFHGEFH2A0FvPcPC0zfR7Q6SrArxVi6S9NjW/LTAxdy25+
Fz/xVoVq72Ud5JTrSerpy5nuisPsuxyWS2fv5HuSvRSvAr+7hE8cgLQqAeKLQb6H5nucODDKte7I
yfSFlf9BeYyODOmfQOQkZIbZN2n1gd9DO4IsXfX5BDsxYI0Z7WU1uqZx4bNAhXy6QW6drlTZe9Gc
6KlqKb6zrFXLQD/iduhcB/zmIp/ONbFb5mS4bNB3pMS0rPdcaihgVRcIMoirnj4h0uxLUTmF0E2S
L5iZf1XihcQ6jm0KNMDaNMfPMeJHTSJhbAAAu63t9LtIgUaQpNmIy9HubjV6KscpVk4S9UOPCpLP
oaUzCn9QAJpcaInN0sOPif+UKTTpjtxGQjkslm8MgdFkb0WY/QVW+OZayqcF836pAN0qRm0OLGWo
TyClAB9PhncG9YajjJwERtV+HH9hqGg3e57UNKPwLnqn6n6A4YBsV8c293O2+FTjHYB6m2txhy/b
Ep5disOyvrRgyPgM57JwIpZrssa/8vP21pqpCiRp7CJKf+xZT1TqLd2Pr7xRXQlRziCGTNL69Szo
bqDaktMzY6PNhVf+x4/cdrpjG107i7s86eC57tSkYRrwMwkAAwgwtUGDucyydn4kxbHLR4dx/TCh
2MSsxuqmfYE+/k1j1b/IzngAgLDVTx9jnwWClCpyjAJ1kG2tb+6WP/CJ2CUTMEY+jApxjAHYduyP
R28AJIkHEBAbbMMI77yNhyW9oLqhCq2lwYUHCVWV399FHwgCku1Eb2aW5B6vDGSXF3VqU/EkDsjW
j3L49T6UDFj33YqKfHovI12JJmtnQ6D6ElaeOVBmyegvHcbDiqNWJ1w4Ie9zYrvwhX3dk0HWQpyY
I5uEof9RMY89t023nmcYaQ9tVjihoS0IcLhGg0K0OttfWx9u2DEtcEdGSDnTD9tYDnN9VbgjFkA5
pXgTnpDIKoqs2vUlN/Am4YV4dskAq2CBCGZIBR/YzIJDrNeD5Gn9HDJ1pzavANlZQ68k66EwxQq/
BORSYrI/QjvFXD5DbvI0hpQuU62pzSXDvh89/Afj8wqRLrH7YAD+BuJp4MO2fU+Um7dcmefZBwpM
rzOcnhIOCCCCMEbwHTMP7gYkRlzynK99wXdvo09QtTZ+x9fr9hjifcmdkqISTALXYFrf/hdh+GOk
wGi96DuGLo400XSHHPpNVW7k3GPYdVg0MwRNnK3GWfRtL7L2ycxgoRKCn7/OpOgg/shXGFUem13K
NgM3K6c+xzHLgXvqKHvRU1UsYkv2IebEjTEgHnxmFHnaXOfQRG9T1UVjTbDDKeNznBXO319Qg2Wm
amWABAUOMux8DO1+5MmfsGiA94tGHLP24NRefaMtgRG2egBnxoA/k3dYNa2a1ZG54XvYO4FIHqPj
sQEvFeccI2FqDPhdA7A1AgwNhyT0eWrVTdcQJ1vyyr45SMAnNjVWXN7eVpD9Zc3rIqdIfCmXarM1
CPnLrxO/veane3NqgLkECHDHDMaxcFK0MRd7WRYG8Ppzsy7ADNbU+lmCPBVJ4YuS/EVnC9OOnq8S
GORTAxQPr7sgFnNFpfRkpWHmBCI9xlsCdIpFTntOx+SUj+Aow+VfyCoKW4uWFeqbQl7aPc/dBD0B
cFNinV7/cEOYsg+2TK/sPfSA29etSyzSDc0tC96hixDxmB3C5q2o+BnZmFt5QjQ4UirjUoXVd95V
iFM8bNaEi3xYWT/x3yiRmLRboocebURGmcDsLsd1TN+Qc78ls2cB0QyoNTtRTeHgoTAD0oAalR4T
S4a1xG5iY0xNVNoGIaCgbTgSaUIhtvAOgeZCJrKkWhVRGLqtPu/wf7DGRgYod6vzRc2rrQNjxOcH
4Hy3qUalfKesgL12XNjTTCv0OhDg9wwMMriNVBvKkmtG6kUgLnjpGuQP7Eht1VE/1eAFnGq/lk3g
HQrpL8QCpFbWaaGf0aI82Nvbay0EvixQxMt9ngwEAxTHpwNdlfTElkAyZpqnvpOYzzo2ELGlNomY
Ne+Ujt+L433ci5iymDjY9Lkijxtrx+E47MXYftrRef7TfDaX+6DFHEavNMbQcokzefkofDC3DR8K
J640PQ56gj3h57DEll7//X+Nnb/jKbwf5c0q6KUNAaBYdJ/cSx3XSnX6pq/V3W+wBIbXlx3N5IWt
XJSqyT4H93cr+lOaYMB04uBnC9dWCIqowOP6Jvxb3Xj38Y0nsY5MiqT9FAzSgbpBsdkWw6Ps8U+i
tI61GkCaV8JXC5Ko8iEkU/dBkAWRfBRu2xTkWpH6ZmbyGuU+q134VvYzlUrTVy16tP6AQfNs9SCf
VQQL7Tbfm60N5vjgL08XnEKzmv5urq7lV+MkZ1BTonrfmMCVrIjx1SIGhqcRS8eutqxp34jGYiYR
tVTArXlyiSSZFCfUbp9aFvh47DhOME3cMVocACqde8dnDRP26zHRwZ8CTemfEuL3xwaQFcl+1bQl
r+PIdZ+qkhZehpgP2KrGet8NHyYfQGqG3JqOH3UH7w5oFpUfCc844flL0CUxUFicyFv17SPJRUBq
uIkrxi+1rJwrtQgLim4V1fEdt//eXFwqWJWO2ikuud7d3fXAgxETPk6uJFU11AispA5A1BT9qSIZ
CfD3ULtvoyqY72hVuLPuJJYMiGbAVrQ6yCNuMS8DwfgKc5Y4HdE3BA5/LojDs6n4AAVJxuVzKqZs
pyPDdFioidMjM1v0Owa0JXsIptKhk5R3nlcJsU0OL6p65unPsZSNOVx96BeMTmDK1TPoY4qXcjq+
Wyz+DiZFdmDYLo05Nu0SFHJJqE0IcI+BuNYov59IX5PNVSqvmuPyIDfpjIqIcz9EIzb/X5+18rln
cckeIYYI2yDsU5MRyGaG6aZqQuFoq2XIhEB4PGBcGQtq1pSjkX+xI+FuqTlRbwMpmCcihsPouKM0
4IfZu8Ny070kH2Ci63sWZkwYe1hYVwxumWnn72wemZnaPZG2XN41buOs8X4l513UWmujoYtL88bA
2ZuOwv7XTo+PMy2/aLNQHucI/ex4WBP6iIBsaXzB/yS7F7wM6YzFHFE5w0vbxK1CiXyUv2G+/xOD
tbj+eSsrbzJLqA2XLvLlPKpVgxPe10tXqB7nsIAHGrAkdDkWYFy88/LyxfFQ50ELcgby9pQ2M81A
firVAopBnG1uRKO271oYcosOeEPpHVxbuZxwY8C/pa4WfSev7xnYjRsohxmTw/Rucw3CQXIkf/mT
FQ4cAtaRacIsmwRCdrci6WlbPaWG+OpqgOKWUN30CEBvHvR7oRL1XtGWEBC5MTw21Swy4Nyp/gWZ
aCHp8aoBSEEEq3/YEOyERHZ4FU+1N7bhnSR/ss6zFtXMvD62LazjhtRvTfP7M/YyHi2VenHi/FdL
LLyr7zH10ZhykXu9hu7xYdo+0JvONTb6OeWwbFZ1kFAq1cQ7S1Y4IH7XwD70ttGFIoiBdye406t9
9Pjq6jXTaQBIBBZTCoX5aZdySRQVnoMUR7do5eOycm8/8w6I5ifL0paTf68Rm/zoskuYtJ+UsGus
4bNQYWjf0cxD5RryzSSqYPhG03vpbTafJKV8wCmna0fo5YE0jEbZFyEqNHZR6JNd6+w0U9heCjQe
8XQELWivyZtOyrXXKnZQu4r7RSibBzU5Ai8XNhEFI4SshV77/OyaqIHkc2rWAOXyoxVQ0SZjuVhh
c+e+Kq8anVN6MrmE7Nv4Z3DV5780sFqDJeqCo6pBxCbWH7qioAJUDC2T+N/C+1F9cSjuIvH/81eP
gJlWl0DChj65drC3igfNjmkNKfe8UFAiF8YvS1KYrpfqToDIXsFGnX7RwyZ5Tqwzw2W2hbseVsC/
gxLuaVhM707bnAaxdyWizgfx4xqvF3++WBQj37qRN7Fe2+70X/fj7tUrZui8HXnqke6tCf6b5pBH
AuwLAYogUg5NMt5AqLw9dcTXd1qzPvGSZKyy5l1DSZbkhw4QaRugGyqmZydP9EJ0FV/tE1YrEUkJ
yipixnu0FGdUAqzgmaW/E46nR3FSwl+bhqrtFZM+kO9fNxutsO/x5CeA3qTyKTnsygRnhDhl6Xi6
EnDYhm9wn7sRHPNbtAytbVdekhuv3g5Hv1qGcpHyX64vypNvu/DhU5NmzND5RUHQuERWvCc7cZmN
BGL+Cp7e4oP1CGjWKoub7BoO5O24JsGUXQzp0Oa6CyEYYyMIrjdHI/5S8UhkYz0FpOTpMf8Re+8s
pS0yVJUxFEFe8h3EcAjJdGoxQjLkF6mtUeEr1AGaC43iCaS3SPlIRgpvZxR+w53XJtl8D2WJk5Hq
CGsJc+HG6YuxvtS/tJq/gJnqBcBijgBSzwH36AnJfLyIcjUnqY8P538AOwsqBv5AQkGDCNsmlSSW
Yx8z9oEza2Af68V0qQMRO7ZR6P1UcVConX3ZvXXnlnVzB6JIySRYOfKkceRpIfpyVYpHzQFfRMXt
6xkQqZdnkKVXmcbr9AHifBOMMLGBLFvxsMrlcFWoDyxWn54LvHXaLwjJvoLpekkvbr7sUsRnDCT6
1VYGbZjvMviIDFMB4G+A4kSk2wDR9szkmNVA5V5FVvhGgIbgto9K7DZ3A7umhJBTqjq8Kv9SmZww
jY1Mje9G9r7xlgKdsR47yRphIK0zfm12k7SbM9QZGqeRG8L8UXlcy1hYUYNpVa9/8WgUA9SlRec8
ouF2pphrGaBUvUQBGbubW27Km1vgheR7CP8sUKkFDBjC53jeRo3JqtNVDfHLKdRQXkYrZisjqZwL
zxk5e/iTgXrxPf+REzHwuMmUFusMraqAs2cgxWR75lyqlURorFFGkdyIQFJESDtd3QYn+moeAqiZ
Sbl9TCpTKjmliyQ7i2Kk5I0cshLCHlNTXPo0ZkZz1GX03/4xRgC3EDOcBc+hqFvGuo6YWYCh7I0n
ZmiyoslTRJUzpPCiAhPK+QJOzA+NkdQlqgY9BmetlxAO+uUcbzQInDllSp7U+YFWBm5n7LdpXO5t
zYy1rJP22lsDB/FWiJxNKNRqMj1zJvjEg++jdRoAZ9r9nG5igIIr6aj+uQu46PWzXezeZZQnGF8s
Sj1vrRs5oXH7j05nocyZHibM3e30pwdgOoPINqAk/7JhlLArJqmCibxB/y2s9UznW/4eJe3V4HAf
3f1d3exD2AM29qfZDecayMYHxeuGsVpV+Ev9OJF9/0QUlJffhqC8m/K4ziXhgtfd1dobpmL7pVs+
lLreRb+9RjPdTOFcbEowMHC+2ueo02bP7Zi2uDWk+h6FxL566e9brStvH9+HptvbYftQ5+yINe/D
Xb6XatmAxEYJe5xC7dFZWshIs85AH+QfsXe8tLKbp56OxF24JiYCOTh8ze2J/mOA9xRVhBeAn7Sf
E4uyFXHKNcmRG/duIAwMuB2tnyvNZCX0EIVqZdSCgCrwvmwGkJjkdreGdlsWePzsJrr0TYG4+Sou
H+VA+uJpj9SG5QjVwejQnkHxbv2Yt53+CHLTj2g0hJGebZK55+7Pp7m9BACy1zS/F9Tc3QT3Gjv6
TEeS4k246vaA3eSYToFgBcEKYqsjQeIWc1C2irIUf0Hz/cVbw908pwnbhVb26xGe3TTyGWtEW7i1
HnyxD0VErdBm3BJkWJUfsaydTPi0VN67FsBqi5emcg3ocOaquM0Xj/qXN9xHnvXlx9IxqRNAh4SI
n0h5/ZIBhfPk31DtiTZ6D41XL41/VK7YeGZCygyyMuDaSQlllOL9OuDb9V1DtoASJ5Ys4J4stvWS
wIagHUtO4uifTKApNIN/PpiN1pLtsPSK/3l4zW+E40X49LI3zdlZXrznbsUjan/XR435bH9BsgDY
z4joykFi0XbWV/zmLE8i9mnqXAW+7VLpv2DHv5WkAA36raybWVORpJD18Z0KTFaSt/Pyz2iyd51W
z33SOOszzMrXr5Bgn0DdSHYGzaK+EF89w4Pr7lNTR4B/lgpBSnECWeEKy/jYNTqCoXZzuRMHVgkg
xdMbf1NWxAd5ps42K5yIelffH/geMTsFivPPwCXnK0EtemDGJUo6NSDnM+DQPx/TQlyo0xP5tatD
wg80gH3zsOI2Dj6l3D0JDouS3ifgvUfQbG5NYsZO/Zk9/tc/5+JsW5/L2y7rpwU/qDbhPELj1fuQ
D3QQW/R7kca85JyDK2fEFwKFKTq0VH+1DZ5pJfs9dGuOzaJVS9CNa3f6inLvBO22Wjhbh8dTL9uN
Xu/h4izhJB4zVKAJ5nkejjKLuLH+fS9b9IwH60iz1eDNkViKBjkVJilxCOWDRZUGrV/6fbkwZ1Ri
XXWOtszyMcP9It31fKup192FgV/CAxo6ZUmtisCDFkT9wyg8xNCZ68j907teJzGmuxpxbV9lAWqd
IPfF9dvBBv3ZkWA+9Yxozohsuz6FpBMoWuMoXtDm2qfBYVtGdicap5ulcpMuZnc0P6K9joXpb3iS
Pl1PO2+9p3XZR8tbW+f539nJCcZKzo2VtJzbpyb3MGsboXERTCvPu/OJnhuRWUd/1Pzp+3PiTKjh
9lcjT0uK3io4KpBL18h7hekrJYTlU9Mr6NBt21jwLzIkwGSvsO6Mo1OF6t48nDnLF1Lui6p5d7le
OhLoL4ATnBkkj1e5M31MrCMCIbx6sMQ5E3WXpv/nXK1ZfCU9BeRxk6GRigoN06Zw7Qix8C7hZm+9
B8Z7ivtscCf1o2CVqwrmKRxcze5dC9q8qLMcL3mGKNif4qbJ+r5BJS+tZ0NkR1qeCr3Z4+XZkgJm
pf7MWRYDhR3Sx81x3B+Bg48+pi2m6bxKbodUUAKHPSjSb3zqj1BK2vY/lC5VL2LJcOKyKIPvitpu
qyG9YTKwNYOJStOFhng5o2tJt7WsQA/RAwkNlBpyure81vZxY2sFbFemdZAUXtsEpINbrYz8MtyR
FinIoRjSxfb48yXGvS7l/I4r9mobC4RlFHWawpwCeH2b/KbU+ooF7efFXZdTFJYklFXzVlpmpATN
jlSoEAgNcYQHjPOxn04W2pf1SmpMDrV98L3KJwfpc3+YakDopnQCdga7b+FJ/Rpan/9fpvFg5lqp
VWAzAP89h6BF30URl+MCTEz0kcgOkyXlsVAl39hM9+SjDsxFt24MAEnclETF4LnXQmcOuz9o3ky3
jbCgL8vpo58njKgLhbwZ2g+UQzrETz8xbm+8dG0T+LAMMZSNtFr6dotKIOylZkGTMsVy/WznCOXv
cx2jR5gkGeeBXZcznOCA0/WmN+6xDIo9nXK1w3oCjH1qbok58/sijTzhF+/fr7MKo/nwdWAhcJU7
8HLpd2mVeFcBQTwdj/azVNYYKpbu5Ca0XBL2AGYSAmgpfDOYAC6Pd0daetizNA3FZWWEHL66Q09+
R2UpCMaNYOf4+hz1lJl5UdOFFFPPGzJsMg9JfmDrCRglZ6/g0hIgFOrqr2Gx4znivMku8UMjV4Yp
jBz2RDUx+p4EE0GZJ+dwTW3CeXQmFAF0WNMr5IBI+vDEQ/LNuStp48S/LOTPj8VaxFJR2IhU0MZi
VZh9VPN62FYER32jM10F5ueJWUQDjARHAfRikuQKXDIKq036uqYjrhz5TRuIGl80zqm7pDidZB+n
91BuFcy7Ei31Y+iREMP4/PDGi9O4vbeHwwoR2zK3tKkm5RFpnmqnGQ4ndKDkwC/pTVHiaINKYMuL
y90jFsVX8JvbO39JPPFgDXMFBNlLVMFljZUiy00/zTL3W/ZjKMmxjXL2PiM0roOyoka58FQIJGuu
aqhGeta3vahqwSwwt1zdFPqPqG90twz4q0WjD4avh7XxInwbjdcIbVIaUVKQ5+F3Rl3tr8fzMIgF
TMzGVqSD4X63cvAXt0+7RrsR8xoWvuSi3GShLEEFLr3qigPXnLMn3c6jZhrZbLn9zgVPdPpTMMVB
qFtz+8T41ziBFR3g8DJNqsCzB8L6moSsEBeMJ5VgJsGJgo5Z2qO7T1719ZZPdFw4msicPEIHlu0y
m1EnYCitf9+SfT/yKELyMwzYFxGdr+BIBElud41jniSaoa8Q2b938vPisaOtCVQg7uO7Z5m6A8EU
KjNIeW35f/DPVHCXbg/h1vJbdycSZ7ntJ+7+9FqEwCk/QrI9pqWg9sef0dFHrFm31RA6cxwkFd5F
Tv+u52MNJhVEAuvmTNySV+4YooQX/8C6v0kaw7+ErNOknBXkr+RnmD6tLla0/j71Y1t8Iwiy/yZF
oImt1vLkAN3BTgmMbbninmb+1vF0ot0NdaQZss6A/tgY7l+zz3TlUCuqgBlPOLzBXs555O0nLaX2
Bgkz5J1asKNpraFcywWRdH4E7mKNYeZUibULDhZd/HIzDrf7zJOGpWRUYpHYS52jmw5chstA0Xhu
7FM7oAMoq05jO7H9fcdaEq22HCdE7ubDX3o+RSG/xhvp+cfnTEsBHP+tlQYjidZzG8Xa78YNX+Yu
h0BiD9GYsV6/GVpL0UYBPThctYk91T1W8fivf3RLxMotLJfptuBlDnOmKhnznwWvWks53RaWTTjV
ObEZziOIpPsoOyscSH1+gQbGXBy1HMX3OcwwzWu23/Zt/9O+5yhbbX26gtSlihyKo2wwFQqywAnA
ecKkHt1PzJzDviL/+zFfB3034K5h6dSW+PBkI01NtCfQSVMrRv2BhICi/8KHF5G7RgUGezvAv5Kj
ybtSltXoMr8EHnGcnjSFRT8PqanrdnoNnNnV2X+qH1PBqXG8LTsAcvG2NkN61OxDc+Qe6Kt1q0QX
R1cPvQlYyf3iC3XXFTDn2Gcf7XsNGGl0fNuINXYmXH3VqytnAV0Nw7XTC7T9ZHL8s/uNgvV3D152
5wKkY9bPUcrk2Nci0/RHQxE4GmTkF63Kf+IRZNw4wQoMuisTXGiq0LhQeAGCbROtc/r+SSm0IWMw
VgaoBz7+sUb5KBIY7OYd/JE0EQ14HF8PFvX40KtWsvcW6LcwXdpLnXx5qCzF1qCkc6UyQLOkURBz
L6PHgCUhrJlqOLdjRIhBGuMm9zPt2g5DhjsEz+Isxh84Tz16Pfb0JjTPR0aXM/JqXIxNcUtne5B7
dqq0mdNEdhbM4KUMIBANc+u52giqDfbKVwtPO2QcrrclQhun5lXJxi0LXN7IK/BMr0cicFEkgUWT
VgPjDN2BTXhHBifjNdrw/7wM5vI3VKClya6dTjTpPlfJVzfnKsNFZyj65QpMrHGBfgvW+qJ2qljb
Swu4/+GZzx7ivsd7oE+cwstsnIhmux+Sqf+eN86GNVfr3AxEDqgiwAHxnjH9heoncFwQa8DJ9iU2
nUjdMR/UTHhYgsGkttwYq703ZjZZcJSNe2VVZeB1Y794/wJ/ip8Wb95Ux8S+ktgl4Nkzeago/g25
FARey6dl5v6fVakLJlb6Li512AkyjoGZMLxLbL//Ry/JeCtcNbkkvwhXbFHGZ8X3OeMObHIKuFUw
DLu2jsPNKc+rDObP9DUuk4qxVhVrv78maadvXzm8LWtI5xZN0DS2xWDpnKtQcOL+B4DLeTaHWqfo
I3/41JSmMnzugP00SKgF5cpm49+OOoiZdwYvgfz2k9F/ij7AbvDLmiBoiUGxGLr7s0x+JiqVfpd1
HEZj5wc4E56gHdoZE6Zy9PmOpBzo5aTCh/E8jb+WVcpNTDk/7WsiQk3mEJa9uV3MxgRBMnu/dZSi
5u3fSuGF5yElGzLTK2UjZKkNglkvQMM3KiF1pcOz3p1psIV3HpauMiF0oPLkSQ1xH9GNzhiI1H/S
SYkNlY6V5zjumDjS9squXibzJKE7ma2A/YYEU8EB+iAN6VNYLSWINOHHopZ+hv95zmkv1BWg1+VW
Kpl/+uQ0c9TnwYKDBcAtgSozykNmgKsehc3arxAJKCs8KEmExNbfcUJa9MjSKGCnvyWQBwIUxKqa
IaNakPS6t2HASXhZnx7CKkcViBb/KCj0RicVflWii38qgs+uCc+555Djl5zefjqOsWBSJPZi6cxa
a2ERZD7pL1zZSkdtcm7R7Zl0DKW6GaPIEa60jwge9q9jAFLV6xfS+f4RtwT3oY1Vvoy2A4IQwLW+
RZdFhG6jGxRfZGMNmtGzM/XP3vkasVyD3fnKbqWJ83uihLsx4E5BzL5JXqhydOhbRvh0dHKC3O1D
io0m764P5FG4lyZ4b90rD6Y0+HRvOky/Db7Y9oOy0ho2zz1KczLwFXPw303ZeMaZP0yW8irxH86P
TLNEZ5j3ba2qNMG5x1HvWUfkD1QQrfSn2/RyvOeKENH2/QN8akMNl3lHHAFDEcPfNVMfp+jdGeiM
/kx8B+SvXoR1uQb8fibKF65PQU7XzJm2voNFlNHPRW7CobbT2aMXCEkNzWtbEzN2+rQ+34Uy6hOX
pULupy2jylVmnEoNOIV/ADZRW9qwA3SBKe/UCUiLfjHcWfxlZi8q/PDfWpuipW04AcmBmvlBqWjA
dFhTuSKhoI6C9A5fplqevfBEZzP/IkGHKjKFs3gU7JyUesjbHrDvgl6PUYxoMgOaLKY43WvLaPJo
te2y45N92tl8ye1kq6W7vz6IZLgHmV5kKQv5MDIuBBj/aCJYPNfLXU7f8D55ICynefSR8Lw9aya8
1YcLVReo+SYmhJGIBAeiF4NRimCSz4VkkG1x6WeivozuElKrYn02aqUtEVvX0y3/sJtn6ktHf+5g
pinHGrYCSAXnjJ1tUBp1VxmzCE5WLiBv13+QmGc2lMzu8ctU6zculmWdtKiDGQnhtg3hFOHBbRAK
Jdog9hSL0zT2ab8LueSzSBt4fmeGJKKKJY48yxQRGh+Dgw3mXXpXtCvKwcbmXsilCkY4sbFI5TDk
Ia4jXJQC6Y4TTA+xHTW9waaOao+BQAFgODP3KR4qI3G3o5a25wAT+DUlwp1XMJb2mwb1Qx1h00Pd
mkQvy1QWgH/Sb4WeTWVfJ3nlv1otpElOLLOpvTq5cierUpdStCxd1E6C6bc/NYquPRT+bTo79HyY
E0LddE8Y8loOTrR6bAGtXSgGmIFJISwmt6nXtoZNtClvAIZroyXr18qxQT5pO/JjEfHKykicRQ1t
WjjAgpvLxyZB+2yZYVwzsdeiEquiBqNlXbKUsi+nRPY800ZYH369YGQ67OlUFyUjecihzur2ebl5
kvdfcaEMdIAnCxuc+/twJpT8pC56i+MvBGNVhqmwR292D7Gd4JVvB7bEdd94VqfkO6mXAfnDc1n9
ywMCTDfPz37n+LSJBE74dIQMGw3E4yoXBIDQp/BiEeK/wrGI+1Q62wlxce29JLzVFMFd+D8yrsFV
8TaKfXdzC1j77JTNz9kaxA2XL0qI/aGest0Umv0HtBlbp+NTuSQgUz+915rIlmlC37vJKzz1Y9by
9ju/XtQpJPGacwlRPYp6t316uraT2IKJfEiTNs19vOvTLvBormvqWXRTrmdtWDUc3yPkJAiaKlQu
tI7rgr7HROUWvTjU4/QXehkHxnzH9ZY9Q6ECoL1gV9Q/rbhRQ7TotTIvdq39sSDKU+SNlqSyswyn
Wsu2PxNKOJSpeAgh5EdrRrUXGaDuymBDIfd1veqdl+fBl1tqGAXCdgUROVcaUJd+29m2RW7Sqlpb
1PEumVU+TgJKpXC33Dcjn2phfEr0MjEIykkQmcHPs1b+YVlFKeUUZwwredu45gbr9AEUTc+qoxHg
/C0Cl30rTH+V4c8k5924R9eXxXqDAQ99/suWdwhuIxT/RykV/ClAHxp+VJ52lFsgZnlnElYXzJuR
dXoutC+UeAZLlROenZiIut08QDM4BGzxfHIBilkwNHjZIYRm3lpamhA1mza57Zgtzud0CpeTvMXM
bq/w1FWBbHQzSuiDO79Vimiy4t+YQZsrweK7RZgdmVXSy/XD0qY+adrr78aha+KvGt9j5ucITtJq
Tchxo/q/4hu4fqEvviJPRuKYVXFZwP7kgYoeQL79ttjcYmPSqdwX7ojaybKea7JkRebXZrBB1ieG
Bx94syYAHvJ6TFQJ+/xKSAmcCbzu/vlM9UhNAHc+OY4U36yGBRZjDUrT8L5apRUJv2BfqkW6hgkm
EAP0yxs+fCzk8znSI0Xp4H4ef74LirkUOdzfsmoTlGEmldGkA2y2q5utx1le8EW+LRjJr6ocB/U3
dTufs7ZnqiAIqSTOyAQE7aro1ZmUl19FoluPypTKwhHlP5E8eaycrohSxmk5/J2pTz4iWPxLGJu2
2OPAxyMhUiShsDULIzK+aGMWg8xs1fQZEUAMr0nR/ZKK4aJ6cSyagHfPr7eVG+4M7mtRk+JPJB/r
Z37AhZwNp+uC3Gjuw3TNLTAyOrImqiNfnTXGd/9qLWt0gqs0Lvy7at2BPjHVboCv5vLTI/4DaBQ+
Kg7bVUu/NpUBzFHZZSw7E/81D0Cyox1P8V9atywMYUrW3fnR5p9SvZ7fUyNBpLz7qGXjcdWEVb1F
zEc/YGZaJVykI6eaCa/0rvPTUftBge3z/JMRCsMvBgDx43lmS/1AoskU9xw2REyG4bioLnqD47wY
R/mKOGnQ7vGyE36EJa+IyhcJJCIkPKiPh2/bPvq3765CeTk0lPaIVbGqKuQGV0RlAqePaJBLfROw
WkMugklIzoMgu6U7YdlHr1bxTqHoQR7eydyB0uqGuuAReTv0btxsD41dYUauoh311UBEho+dWiix
08vfYPEq8QYi3Q3WCC77z1cQs2tnbvzQCKfkBZgUcx5OwnIiy5sAcswzeA8vdBzUS1W8BBe9A7LS
YH2vpz80NpPnU3JPyTdGJDPgxTg66uOrC18f9X0trY74MFj5X6ispjVI0QwYYFJy9z1FXsqKC4Do
Bvv6PMsID8vhmcXrT7UetsyaZmRutPZai4MEj4Je9tixnVGSn0QR84HGIfsYG8Ugr5UTwcA8taHx
sPFX9RAAU8uz5hBy2BjnOrupVO66fhzP5aTKlBI/eFXC7PWeSnUdcw9LQBb/7aD/sJmS2R7N3CW4
pORd2xQWkQ8GIDd9R/oSXc+roIEEAuMEL8wjfHnQCCzSYB93wM8Ibm+DrzifZ5b4JWDghHon3+C+
1uBf5vf7kb1zpLGghOL1h/+eulx+a89sHBxS1eud6Fe7EFz+9oEv1X9sOkOQnM7RugQW4i8S1Z6e
P8zEr3o6tQtUEjsKsNCGYOsrYvLxd7A9d6H1/vDwdRulGLOmQqkxQ9b7lRCmm2gxHcT8NZ9ixQH+
IejdhHDWO4I1n/x0s1w5DdjoF9fT/IPc2XH7DadVyHaVr/TfVzldnDT9UtOm//UpJdISzlFjhivi
NCN3ZH/AlxVZzdmxdELcaImzCMJ6XnMLnTqSMBFQatz2g8t9HXlxoG6oxIh44Soc+NUTmVx5tRTZ
Yd5eofr/cevA2Fvq4BUUiBxmStPUZSiu5BQLxRxCbz4zEpfJN/G732s1IH1vLIREbHLx0hewSMDT
JrK1yfJHkVJsRkh2NhS08qOfUO1d8sabPJV2Ti4DldUibFjMvEWS9mkwscRiW5XomQlBRHvciJad
luhbe17LYSMeMzCa/I4iMsNUjviKGxqyI4xhBrbAaEycunzc9jMjOordAbJ0XYKR5HWR9Y4HxAui
Ey/GKM9/qrVoNIlphAz8Cgn3lU2Z2K0KJZodHbCzkpkzBsnaO9IwwobAN0CqkIJqy1MoJs3nFqDY
ftCv+sw4iiGSmKnCXZaGxSWX7sCejiyWq6pI7v6P734bcQMuAepeN5iY3GH/qyswPC6jsIfAMveI
87/qR3Cz8j9TS/QryFEoFtXD8DgUAcWwf7exkIYuBD1do+in5bCqIebMUa+/M6wEP1zGsZ0yCfhH
z7dbRM9HlQNIIREpdCdB0tx6g7WL5KjSZ9fcWdkuvMvtNjMIIDd5kdeo89i/egxkBFl0aL8WCakK
ObX/PAXN0SSvOmpmecE3OZEC9eZh3L/RX59Ai3oBbTdRmsFc/1FGmuc6qHLqJGwFoZGHk2MtEx3A
4YMhyMEoUDTYumQQzfbyVXtILjxrQ1/B9c3cItGdkhiUxnjX8rgWxVASWZ1Aor1EGVUlInSGTS4q
ghrlWLDVfI80IxJmk6Bci6dRqgGgre5+ArJyPBiKRMr1+JoJcxzOPScO+Qa1OHm5h/YlX3oRJMig
qB65NU2p6GrgI3VkA1XelvHYL3wtHd4w8YiWDvv0TOb+DbqJ61DRsqb+7ZR37EMPIib+Y/zKDnkg
kYKw61VuMf/KzCEvimdAWuETfCfvT7A+f5KO285YpWtCka/tLaY7taipqz/GRosCWr79gGSm+dpu
Xhww0X/8AemCNfQeg8fOUa4rkpvSDJhjC2v2Uikc0zl7rMC++V3uIPtMSmi75wvR0Z19LJDc25UO
yf9aks0YX1UkUd/Wt8/jkEuF+pt7JWaWsRBYy8aL+ivLf8RhcSNXkC5LjMAlzybry/Vz164pkzZO
lSfrkxK68kdfQ7XkWW6ynaPcr9SPVer9pf9jI0dHnKt4HmVcG2p9PUze1qQlpAI83nAiDxGslRTO
UMZBBYVJojHolb6qhVbFlQNQX11aIOH7SRnya2vFn/A7J08Xc35UcOk9tQf4UJ/l6G01xfjRANU6
XnTosEWMNbKQ3TfbWAC36YKm9J1e+BVmpEbvahebcf5Yf3Vj0qCZpUylPcqYIwM4IPgmnuaaI0K+
KPURDyNju0GE3b5qZzaj3zJHqasNRbPsjchAzWtiO87zaWK7ROj+J1poUDO/x4T5XxbD8nhbWjZt
Arhgtak6T+vDjC31cOr6oIIj6U8mEUtHcwOJk4IaVYGrLtM59QWa6duGScCIWd7Wt5D+SY7R2UyE
9bUEKaRWVqMnOWsPkSbhjM7BlUi7nTpul/u6pl50h6atEGXpMYv7wL7tRtdOikp8b9Qdw2amAgxB
T85+coDgwWFkz5YGyr0zeQueAI0LqcWeXVkpbddkYk2EPmANQuucphv5rRlfMaDtrizf6hu3r+cb
0q+qgTb3RMkiH0xSVdugvEPmHwPjTH+xS8NC46zqZ66CL7WgrYuEoTjFWYfaSDlsR6HvzQCXB1IS
Ikm7wRYC6aByZMt1sjUz70phaEkVg2ZxmsOB9tFwrNzyRmhT5LJunAUg/Yx1Yn+595QvQ5yUBVsL
x18znDpTTNEVbVh3eSwztdpQ3l1NOI3clvJLKOkYkPMe2xXZuK6s2MSdY7yaZPp6WVIgLvLH0Hek
uR8wHNUr5/s9ZdXUjFEHL7q1J0YzPTk7H8R/LLTC8TIeJIMT9KG3nnVO4/dYkegecf6hnoWtbVd+
1bPC8sDKXeHcAMWiMLsdBUCQJdbcgvFOntOwMsiK4afu48d6ZdcQRwkDdyXQBzQ84sQ44ESoqDyW
ASmLQW6cbQo9j1NOwT5drdRS1NstZslctIDTC860puk4aeDzq5AGQFP9TQC22pvm5chwHm/xCktY
KkEArl01dYZS1rud5JOyIR/u4I38YFCU9y0aBxqC1Y7vZyASDv5+tUdTIiwNZWhJN2XvI0WOrkSZ
OlAFtdwZau+UnBZExlluI8dNmlmBK0INx6bD7O3zO17O9f2Cfn+xf1iQ0ZA8V1HkbDEMeW9FJ2Ip
cncKdlzUr32LEvc0DfwdFGEarVlWx5JJywgqPr7joE6CqHAfyuYrJ9iTlZKVf44/AChyKzR3lL2e
aAW0ykOS65uYPj9RiZOlEbDt85Vdt4+D3IYifGeigkiQRwkFuJ/99lY99VTBiiTVHa07Vc3Y6v7V
lGiZjlo1h+Z1xpxxW7D+BMdu2BAGifxXMIgFtjWIIwYeuZNOK0m+k5pQHT+e/ciOlX3IKjiHetX0
cyrgjR98Xu8MoZVqA7XIyYESdZC4LyYatrTyCR1hX+7DKGgsSpw4GB1txXqzu6fQsxCkcRER7SD1
02DkZO00n1xkMgzK1RBrmvah3OHbcU7mhiAzsqxYh6lNUHEL2OPj1B7SEqa8+zFBOenHkr5NwEPV
UdqmHPtnaAoxem71u8pU/B+5hin/qs0pacVgXLzlRPOpOtCkHr+MHieuo751bxHNVYRqGi8njNXQ
9AqEZrhkULfeRZwoqLeVGKB8k6AicURZdPY6TkfBcDyBuyplnHmzapPdP2WTugGfZIJnWbBeOuzX
vDk/AqIskSWqKp6/F82zDHd9Bd+7LIoflshxHJzyADdTjMmV6mx72+4eJTOjJ4p5Hb/tZKzgH0y+
UleFD/W+1ZY3ZjftS0jvLXqM8nAD5N9kU60qFzhsrLoqpY9UecrvpIRK0PU+NQXj+T3EgqN7jQcC
70LD2U/vGfeP6CjK7JWiao7ZZSPhDM/oEvwSfoPQH15CSkHGMSv01M/Tagpp0qCHw83k4b8osXXK
jQMDAknJFEQv249WF97McYCsVtP+zWUOl4Nd1oogwJY0kOaTelmvZKHPUgMmlmI494Vgp0URzhNM
lZjWGk3HeyeRne+ej63K8qgbsHIPK2SLAu0a7H0LIt+RFXQDfSyvCSK+6/hzCL+ab0Fe1NexT4f9
+UUaOP7T2oTo8cI0z11vumgMA3QXGLaZlJWoYQfbKWWdsfjb3227Q0+EHUC2wt57CiaECXRvbFT4
pZTQXFbysslnlFg9/WL9Zuvunhp94OtSXOpxuc7j2oOFERRcHz6DTUtcNkVQC6u9XuSYxuz0QK5U
jQpPJAOEQ1X98GYAYZaEFbu7TjLL/PWLfkUeDwtONFLjTct4Ey/jzKYrJvYNCelb8VeZUqKaqmv6
Aw4qzZ9d1FfYybg7RkClOR3EUv5wWYi0OcDfjLwBL0JdpnfmRtVRrJAeaTrUVHKsveruvLacKBzb
e52l9w1B0wX226E2P3gEdQ4Ld3hbinI6s1tY/7IfA5bSlQgWl7G0T9SNJY27P0jOScZo+JsjI4GP
JZBWO85vlPKYVLgOrbk4/btRUk6ccqbmMWtSxoUgEmNjrHGQJsT1aDrG02L6O/aUBVwwoyRuACLK
2bXlGo8mUOn5b9cb6/k6Sc1sxEBfAz9wAVJQF/4YiwQKqP+PCfT3plnRwHi4WbzC+46885OwaWmP
UXFNK3DtctRvY2kOAZ/7nBtSYgsJh8OmgsJngdXtn8LMZ5mRM9I4WvVZWa2AjjkKS5s/SFb5KVtw
1Np1gAzHUc9BCyIdVpJLLvytgrq1D7pHNCdSVhC0HV+Xpp8oAHCYLglBMwqw7bK1ihUkTYz3dH+W
q6c7ApbnTJBs0w8TP5NdT3vbh7ylv5AwTcp5+qAEUf4LubssXaAOUago+3abO8GjlHR0nQfNDbXr
2WW10M4bfraXwlsy9XSWVth3GuMGmL0XoJT2/2dZdjEdBYtM3UszD1LEdcaMlN4fqT9ftl+QO0E0
A0UPnx19iWY4okX90mJHXaFxwHXUJ8WHN/9kYEH1fSkP2jlsWGagO0eVAKrU8gDALPQPzDam1dSo
9zW77iihtOsahotpJc9BzWvzuOQUBDb9k7x8Ds0iGams95mL3vos8tyALz+KD6CMqGn6aL+NXcHX
bHUxD6aXp9I/BYYPiz7LOReLrVn+Bl2lh0Yjgu7V0Kz1JBeOQ1gXRJhbVrijpogq2rZwPmeIIWrK
0xdlht6FBHVsPdt5913VcgeezNZtgn+3DKTi89jg+7OMEHK52lQsrF/nCzGTg1uiYlG+yCTwEwbs
BOSMAirshp9049/UnWUPKTX/SbN+6+ReVfrCID6jkh14o8Xve7FU0o7XsPFR38RQ/10oMgqCSk9v
+y91S1ADzYFFZd2/KR8BfpxFsPhq8VICk+AQFqZBASm3lkR8tYsDbTFJ/RvP5ncBBlEgy+QChOMs
2sWquyWzivgv6Ch/u1ZyUjEL9p6BEIg4/y4rA8C5sOhRzy3IEZh1rPeJK1EQNQfj5hj4axhTo97I
uDPiHQjiUaqly4qIeD8uXPzDwoQpnv8M/I4e5bpQmvSk8FdQBwL3Mao4Aavq2HiWVRxq2YHT/fcG
8yeLC7+6mrhbTZAxzNgGOFQgIOLupq60QSME4zxH7jTn/kf9wKoEfF5fJSQj8spc11J8kBau92L4
eMm+Qmdk+FnNEytfGLErC8gxKMxZ9UJXcAnp9l3trqjD4x6CbKnJ6wNaXJj5/dcfff8L9d2Zyjgj
QsgMxkm+QLpf6qGlmPd1uxkwwizt3IeT9fZpWnWRX7oq1+RyGjh1mJY56qt6MmdswoYnNg9i43iV
/sppThcL0kz3ozDKLIDkniKi6BNsG2JeynD4CXGqQRXaei0aobN1jvB6D1FsGIePLYbxzYVTrzon
wFmKrEaGCm0u9/N1DuU3bAkZiXt7Wa+amEpIZmvSCAWT1ajaftw/6XhuT2toDGgtjDAau5jN5uoO
byZbnUyXtt1E/uZ4Je8xQERXlXd/OvafetWuluwvckjSi+ecB8Y+K8ODJCQkGB0T5toyojMEYJl/
thnBGUFn/EzEan9XW30zd7uh4Ini/1PCiJRNooXaO7zucTtj1adqnIZUY6xZ7IYRTMBWWPD5p6BX
Y9fuAM/LGwyeMkufhn6XTuDFdKdlAb3UyREHOWm8JuHAeGoN1PIAX+FdFG724ADqD8GJZWuHobob
Ci1/GRv9RFXoQj59kJ5h66QNZ4L7q50TDspN5TLcGUo5FXcNWLKLW5CzUG879hd4py9FIl/hNyHM
kZCQdY4It60XMyV09BtBlVTsDP01LRcBhreX2JhumeVTo1LQ6AmOOd/5F7OvZ56J7+JygI4SHGyY
CNVcJ5FQpPV+nmD3lcn6gGujJzDs73DADPSd3W707tcgbosCKaHCy7lozGMCgLyqJhzbc0SfPe7h
LVbAj170QMyuSxQgQ4g/06a416ANx09EU6HP53roa9S8XTb3ayogoFfT8Q/0KOomrQ6SNrMBbL5p
BvWIp4RjmLrxe6a7Gk+0Yjf6C7XrIfegMLQA/TMCj4M6F7Aal/8NDD73kzjqwKnUjgPsloZiJMMW
yEPI+wL5TZwnvZsv4K+ouUZS4CrqUXdh/HeuAWK8/QC6vh1ehlT2u/SYhVGyjJNDe2LenhS5gEgt
vKcVcgGUvkKllLllA9y4RNdUc9bPIeWweON70x1eheAe5Kb/tWaR9hAVrluw97RaqZcCgfKKbm9Q
hxBFpdIbox1aSSlcWtrMpv+fRDXKHI3DB02dp5O9oZOGGEXoPlloT+B+LgiAaI773y7gTMx1WSyO
8+AWqT+msBGLnOizwTSistdKFXoqLMr4x7oruEZCdcKhUf5f/aboQ4E3myaWvhyxln38I3M166+j
XoKegzyYklrRiIlNXlgVrV869/nkmgDSDN8C06lhJQJ0ORtBm5WuOpu1uEkZn3w42N0SLDqgzcfV
vN8cGYOttN0WCurKwKclmQBi3FO7XxaDxT68tDG9bz+8ZKU0ySlxvCNT9XwaHMgBEbkvydudgwfv
wWCBwHfs7pHhhui/V2T2S2i/Zed5YQ6vYhroz6ShFaEbQYPmFp/MgqIKJvNAUy+Quwg0WyaaBDfU
xPdm2ZN+qbCYUM24kYasVcD3xzOTcdeijEnBDD5oB/YogUr3P40GKsNhMKAxQrsDMYNvJ25JEJyc
FF2H47tzqUDsZPd4bukl5wjbjogRLrzkJBFgx33jKtcW2D4i8qCm4G5LmmujkSPkVvjqqXHv1FMh
SraWEAnJCqteJn6EJRxGwdrzNBDydmYenIuoJ434FV2hsJZ02cpbHxyHojkmKjoRhj0zFB46yIGb
FtDJHyfNYwPGgszJf6mg+m10WHjNVtm/OmChwF27EmytDBeE+u3V68lmjR6vAw1K7KYieWeUgNLa
44U/OjYI21TJetNqhD2rqbbBgH9V9EOadehtu6+lMRs8kvrKzeIPtcaK/eJA9k76DkwrwaPdURlp
rDRWkMTCBbCS3T3CkOJg38Ou0tu9nyZ9Fb9zFCANmy3XVL/4gxL5MAoyMPw5yajzeOmNqszLvBBv
ZQ29s/dmbrDcLDhsdl3YJJRwTnfpHOGrR4A+hzgOjPESSshPTRV5PCq0NBG9hRJrXfUz6GQ9zXRk
egbuzAVikg6+3XeJsHLnvXzvLp3Ua8zDaDFuAgkM4fu8d4EqZ7yB1ZGgVsgVktzebt2tcUB7vzM/
R/pHdKsa7O/gSe8+OUjdJ7bNaFgYP0csgvUeFVji+yGMZveQDP2eL3fydOIQa8jmzlcu3CxXE0Sy
d8ZZ1jJfS5xdaXx5MYYA8XJVH/06kdSsHGdllXOS2Rd6n+O2FRvze5yCrc+R/RR39F9dUcKxfqUG
qVuj3ZLobs6T+mcw72oCMaNaZ/ykyhnVRCJGtXS0F3yrk9dg8aNHivBadoRI4lvSOLEesVmV2/Se
5HVfZtmll1/U6MyNiju5RAaSJQMbU7RCQWC/XKYUxTeUXrJs8SU/i7y0vZWuAC8Xtvmc7F40oxui
+iL4U7vTJTdIxFZn3kkgrBk/tPDWL4KyHhnaxalXGl/LVsJOC6HCemZKQUM+e/Wy+55vWlO6+wpZ
1xyv20XObTzBCt21paAwuOUd4CgLObErlKGmBU4TLwolShCbmlzhh4kpZJHL0agZPKrEA94Po+hA
wyKWrcx0iDPDlaw9br0fkeVPYYDopjqwZf2uV3fzIHJbL+WdajPnDOZ/fPmcCcexGpfv30z7w1cY
rl/V7p241CTCAvy07ymPiOYk2GGbZ4giN997lZaIkqhozJA+hAXAjfku1bdGowqMkViBJiA/Fun+
BpXCg/QWgiuvH8papUiZLaS59EDzp63M9zMXlyfa0oUcalHMdAKrfxyYaTtR4z74xA8qCJm1S/iU
J4l/AA+8gXXwxvBFsjYKM+F7seTvxzL+8A9RZ+AKPU9PZsd48lGMviAAh/+y1l/rzIVvcBFhc9Oh
V3KijcA0wvdEu10hAsjRGBtcGp9pvJ772D20WwVb4zZylylGapb+fVD6jnEBtJ4dvpUqlo28SyQl
Y30Ebit0KkJlqv3E4qJ+/hCBIqKoiVzLcnAFbypPez1epuytIavVpCwCFmTUZFcgB8A8TFKETsjI
pIWuALkhr82IdemgscLmvGoRuBgU5hLqibaAAt6Q9WpqtXrVaQF3u5loLnsIz59xm6dy2Fh3OPw+
pow0Umh1TqLukeODND8R8A5mJ/5Ql8lpCUVKATkXJKqbpEZpEn/OqjsmtvFWgAX9Jfw8soo25abX
B1xFpTXjwAqV9jSllQx5j2xI45j+jJU3n75nLmuwc0rDm57MyCgVLYY1aLle0FR0FS8XJeJeRGwM
dmaBsaaODhQVjb3VpxZGLxXKSaoXeTmwqzeox7PbEX4kakVDopBhiQFYuICvLSyF72neI8ETOdQF
+U137Nzo1OF2l5ZgRM6aSZvzBFyldA2XBd4dvMmkVEWM+aZJDHVaOYSkWLKojImRb0kICGh7JWBv
ch04YeeUZQAaOIfIfoiOIDnpMz8rmnLqjLpEag6AFLLLcwL2efZPN9BmpNX1Z0Y1iBkqe3w8mQyH
ZeupvMENgLHt7Qx64mCxi/ufkMsHDW7fEZqf+A2N40I01xbr3jlTzaOJ6DtAqibmdJ5ShyEFjF0R
YPSQFzhAtX+nLIsbjRgc6AT8Tk/Zp2lez9Pwxnw8wSxgttvtAsd8ONKHNAWzbEqYBCkldh+MUpf2
GgNUcM9VLLwVo6+ExCjFR3rQxu+Ox5gu9Ndv8wqa0xaTwUBztl7bHLJydVBcdvYONYn32cx0f8Id
VQ4wiQeYNB3Wrhb9xEd1LofxZC32UKRAimKF+16du0wrZXHNBSf+q27n1KPfCCIL8qv9bbdNiIFl
UV6cCIOtma+AeMeHrNV2S2bj4eAtPSyy8IT5uksgKdmFSbQxrfSZh9x1MtvTcoBMU7/2FILtIMjX
fNvQ8k6o5op6OMrLmAJzRYw4P2C00zGQTdvF9IF4HP8YLSg5mwDy+dnS5NmgtAxY5bzPg+HPF+um
PPN+fJpFfnnok0dqgoGbYOYrhZ9e/vjL7VPMWcT/Wzmn5W7mv+d9FjdsNLMHbu7Jo0fOGSP8Ey22
wJlIMJH9WX+zzjwzTTJEORfkI0irNaxVkoINooni3Hwb58Gc+oK9UCQTM+7YTcUg65ydtJuYMZnU
n4oZCjTFmegBacnf7ZHwGkX+VKtF76CspPqwM4M/bdO48P4JjTk+TPdjRefIHcJ+vHy2U/VTXIR0
VvHxT+OcHMZMilfW6+05mSceawXhiAxxIm+/yu7VAYEBWHlTg4phZ/ciZjCeBoRPBS5nkLOdQba6
biW7zBUZsU2I9D3ue2KdiwT4hqxSN0YxrukRzM+r5wLfRaSZp5PAMQuDoAvQSktEvM3LwQu2oz4r
08xtB8hhpeUXwtidhmMrBKd7WcCFQFGSrxTAWgmjJetEPfex6dpZkp0Yo83pragLHT57EvyCUXfV
2zFktOds41OxKGgb3FrgVYtQIsoTbRxE1NEKSU48hKgGPrfRIQ8jlsCydwI89qMx4arZYr/wj0u2
YaEQxcSzWSM9BGDPYeCojfKbE7utkFSzWogJuqB90yBqp7j8+wgYk64NFKKLGuNxcCP6B6+8Ms4/
qZ5CeiLLsCb5Qba/X+rvFc1hHSYcIX+5FpMoWRlJuYDc/QLgqfOq5JSJJejwdJ9r3es8UuNmqWFJ
NyKtvYXyv1OSlvSp7jPYuE8EAAOcyXGbh6KCvwR98GP8R1ATVj9o3b62pxpfxXJ5ckea+CA4HXGE
RNZW4GlbsSeOXTq44qsm9ejTOT5CuS7wMl8ddh9mPkvoYBKBPLL38NexYyE3j2PJpHmnZ110kxZz
tXKF/f3jpzq5mQ/SpcaMHObjIoolwjBs77gp20rDsQIQEP2k9K9ostKCjoVH3+aGLfwPYN6d0vCx
D2JloGvB/4M+Yj5O2g3H7oGDwFhhkmCjIVxFi/F7bYn6dPAcl6XKc1hXrccQnSWPO5GUziXIfyCa
NQoMGzLpb7ygYLU3FbC+JQEjPNPFJscubJZsE1qsYPrOtsvVfzmMjxPGyJowVL7r0b9H8NJdZQ2u
yWyL2m+IvcgAtvTcPvtV+p9zmtFETVtHueT4WCQh2xfgX+niMPfAeqK4EQhjjAZw6YdwOuW4pByG
e9vsPgI1S0Ab1tqQciSNDXmg/6cjjK3M8zW5XwbE1av+6HapQlHLVY8UV9CFfW6Y7t+lVj+VxRCx
qkicvjgE45hAVVmgNbjCLCg/PHa4PDUw/CR0eDeyeQ6VcVtMnA5TwTjBwpXWFedjLyo2vJX65zt+
VuwaD2VFeil3Dzbr5wbSfy9Za/Zx14FO+EchIUeOvVAcjuQJdz0BXcuyTq5GXJldBJ4eVhuIVQt9
Bq01ThuwG/+TIpPjwAcKOdqQensRt3XDhGQydQxR0JQrARiek3hjYH5YZqDVGCGRljkchC6zxDB6
TWOjiI8hyz0VgvLFXXpWkwJBa0VH0bHAaLjpTbeFBfLzFPZJCD4MeqR9hAtPfTikgUtFQhjnBxOa
g88etg7oNkYDdk9hn3mhgvvN3xU1bN7D1/apHAku/h7wp5CYXspBtkDPteJjGxWt6T6b9Z54Oeem
JZ2M4DocepiqiScWVd7qqE19LEYmmmPgHgdUZpIfNDwhcDYXG7Ae0TvYpl9EBmX/kuL9S3jD2cdD
kxfX4SwkLWfFs8G/8KecmClWYWOSYyNORNkEGC2nmZHqgAxostrpLnVX6y4O++VlKLHBmDPpywKG
B/MWuqxyFjR4KSd6rG9wL7DCboTyJUp5UKZMLQNVE8GgFPMFwsB3YSRbYmHQZL5zOVP8zUE7HtS+
Nv2g8aS018VGrhcmMa4CdubP8fUWIJebg5L/BTNp9xxHR1DrdPLAM8E6RVR8tc4v8s64qeetrp8p
dDs8mTHt73umcSJUF2mOxfrWlv7kcG10FnImN0N09MR54FKh9GfD1P/NcrR2lFutIAaLjDq2GWKP
qDxrO31Pj4grNMn4L1EP1dOcHODlaJB8HtuaxG+SMFJgjLAcAo5KurkJ/9su2nqcj9LZIr4fH9gV
wGizO2tnMZrVDJbNayD8UV5bzPzh0S51zOQ9hHtsZ8znwy38pibXin0yW6sCSR7AvrbnL2Kt5DtK
ZU5W8KgaOpecO9Ibt/Kg2iXfXnet6OX14WuLbP5uJon5a+NmMNDjPTRg5lwoVfbvwNiAv/2aZMZv
byicVFFV9Sso4DUS2BzsvNfc8dh/dJho9GHVEnDMaVJn0YjUHPIpndCGk+/MVbotc10l6O5NzAII
RKsznPam/pFpK6f1ixtCChMjwJAj2+qs4NjvG0X2FJBj/WTnRoPhRxCtKFmbZujTHK6UzzBf/P1U
LLd5mKIfqsw3vaP7ZTAamE+q4Y17assjXCIFQh4J879l2x9+cETvpV1eiFdozXNQBscfHDfpF/NV
Sq/vK8G9zpgsLy7jVfQB+WguHLI4Dosb7zCStmK6+1GBDvs+BVfGclLZ2SHpLb0Ym4UU9nhilu0L
zJsiChZBJvS8Vaz5/zxVoJQrMGEqrSmNLAbwayKT+04YODuFXFvoEDI1vwVF4B16vrEnQ5ATP09r
jVChr91BUYV9goEMk+xHc1zBPBIOxif5oWSvJKV6eBgeuRlN0dwul7dqreMlpEr/F2+mfz2yehyA
8HuggiFax5mY5X9pc1Px1BAi68pPRWvVWNfXh7tZ5mEEyukHLnXY+8G1Hod1MmM37uUlUmGR6rry
DzvpxzO2z/iHLvnsfvZnJYq+pbqoVOTAY6QSTPk0z3eFac6rIRweso7r91Ypk7h4MqMQOHzPAfm9
r1XU3/DUbFbWj8HgUj6OyCrNM9Vg+tCHMzUwRigILkWT1DfFNMq1qA9AkJVbqMBjxdHmkFKF/fb9
e/dqgY4pHThbJuvLusYgcjSwjSgHhd+bUuuxZ3w/574PMeqQ55TQq/lCjC30ZjcaBShDQZgQOaj+
xiHfHCJnRmUthWNtSNyvop96ZOZa+Zq72Nn3aQQEOPXozGJvPxGwhWmwSh5Ctojfnw053YpbWj7d
cf8wuRowGseSriQY4p/p+FVwONcmIYKlgbbc/mpMrxPZpPo06+qfw4dvw/6fZJjgaqxSxD8pSiFD
xN+atIHckNgniAeDO1tRYgMa2ACa7uRUutNM2Zy5y8L4YgORShBNpbe1NNrChHeMskFV/X9WSFIG
ucLzKcNYEd3/1F9t+8X3NmKrkYU1GleBQW6u4f70GNBELy+641sf1nMF8OPQpwRFUyG91S93+U1+
AFKtv4iTUgzDC4k56lAOITRHuS6fRvl5v+D3Ghe1IivfrVhrRPxpeiz7l9QLL6vcsmC6nJfsNG/8
spm9VZsk9ir/gKPG5l/Wo5gWxQYQbDMQirJU0V2GGJcODO3erpYKlAb/p7BYemzefVj1lbsPgANE
GNax+BUeKomJNgODEP8BDIHgKbEwG3Vx0VVVf/gV6tLWbVLXemWGTrCwuhw4oTIZaPmntvy/HOri
bclAJZSNXNDSO4vHHYbcnys34bpkfw93eCGxmGiNTDoth1paeFtmFE72AtMZNcpPrad+VXPq45A1
Q+0x3MAYcMNAofNMyNa/Xh6wy3vSPHExKGB+oYsx+ZuMLCQxQHFDKTvTmYqRkVc8daWUWiWwBUJE
ab6SKiad+ITaPriiQMqBs3iDu0I5R/3Fjm3YBOhg5/gY+AKzBK7+zb7aPBSVyU/Kj1+Kl+Ve/Opj
SwyYFj331dN2YUkq8DY5WWjbAWuNesW/CraNbgUIAnKTpXgPC0RtN0ZoA/2CFcwMpqsIbm765dn3
U8iVPPzuNld/8hu/zbTUozepDkIMtNeXO8AIH9+SJkG+7iwiVR0ybb0QnRtA+E9cRgkTwdOzW666
bb4a3tw4fiqsTlnjXWwFiBpKza8ISZMB6xfCtovYCs9ovjyex3ZEQ8ixKnnURMy1kxX/oS2sHDXL
G75dG7lfJqvcMhVj/tpwUfQwy/BkMDet+ox82NLD4HWAVU88ZEvH5J8DLXTutwJMeJ3Efrv0C/fw
UawzyqDomiZwukxDWXLMLlJlQ/B5SpnoW7EOxrX+bcLvwtq2SQ6D+jkjq/n2zWHuNaSTPpzQATX7
s/8qD7GB2U6OH71c9+ZtwyJiDgZ5jqbAqNn8xjaHqXPgs9WSzPjATB8N/b9iXffRQeYb/4N+9e2L
IaC5HBm4oxkLKfE9EdNwbBuPLDwWUhc8tzuEL8OsVkcNm7Nshq3YLY8+o10kNKPueAF24CTCCHCV
ZRLXRqxq9FupCydAzvxhALlREtiiz0M01O+ZTSanQ853Er+pSZBQ4tUKxBzTGuDiSdW2T1je85cI
wdXYKd8GZCzpV4WD2+ZBtIdziOV4svcaLqDoMBS11GFdhEOtsz8mspxfoc8HtyUiYx/aF2jotWKr
GDbW6L53I2Z2IIFPwE9FWkLKUrWJwgEXp4aEXeRQJ9yZjeXTSopQ6F35mH8kQ4bN+KpVKyWL22JL
2UWTj/8WxFlLWE1FN876SLixE9ARoRvdOxzW95Syfciz+69IXQ/2FSsth66IkZGXsLiS6P2pOIKB
PXN6Uzql/iA8jJe7NhpRc8bykAp+WF8pUzJO3GjuJ79W+2NYft9cIPTU9vogiSYDMTnBNtwrqGXj
2LxrOr6NRJDGYZRnGq2bIi/mvXSeOVwZ1jLUxsTB4lp7qDKwYK47mhkb1zLRASXNfitRoGK/z4m5
7+6Xzzj+x48YzWyx1Pr8ClUm06UY38Lu15tLCuythNToy++cg8gK1KJMe0/bgGbat6nZwPUwrik2
/iwI9CKpI25R8ynmMWJWbMf6QvX0GUPypea9zeBB3cQ5sZWhp8kajSCHxypPMu2YxZf+7LVHYJ5J
rRCyr2aZtbD0Q91lKCp2oT2pWcdkO0HqdIxAjUn18zE/9W0WG67o1bsqklxLGZPEN/XFrWwHo4Ig
SzduXb+1OI8uzDMKh0dtivJyuLuBa5x+bWTmF4bVJ5UctP77bAHiBzPtEyZNDdVtAFiOqttOEYgw
TfzHvVbXA84lCg014xfRJsjKkPpy+rOvfxNVfVtZuq7GwVgXXWHgEx3ZszzRcid1T4q16i0rQZh4
o9Qx8ZVO1wkNeEUStqdCNL/bEI63O/sTdkYe9Hs2yxS+x4b9vhnojAjes6HZCXdaGP5YTYAFUtBL
JiQL1kY/wbBwXkNpuWdyDL4CSm/5dXEp0lAeOe0dLxN6gyT7JNDHO20zUWwyoD3tYZkeXw/YQiBi
bm5+2v0s+1ThpjfkPEAL1yf9Q3yawAdlALKoB3BUc533wcK0fmnzwGSxZcpUuBxBu6r4/N4M+KKo
IxowL/c+5HuD+5mQRTZK9LB1lgbBa1OuenpmbPkqxP3qPpQGo+vda8yYEmP2O+3mBlCDfy6mK4Ap
MwxXZKghE79gUBUok4E4arh6RJjxIJb2rQyAeF73t2hlWvAsK4VBthllwV0sou2nm4zstIhwdhar
Yedw7MllTOERwgOlpW36mV2zSZz4ZYeBwzeBfke5QUSKT1HMPbGue4oBlN/8+z/8G6ebevK9PTOP
Y3+lAfALJW3w51C6l8h6qzM/4z+OS6JF+nGM0jRww0yhgbBs+rYqXsOHysQMCEomLo9ePaDAqtcb
/u/dnLblyiDFo9rfZUM9kZdopUmSQLTaZLXm+v0lYroClfEJcIqUE04FuZzO/O5gEDG9T030Hc0M
C9N0ikkRzCSJ0tVif2ee67Uxiho6Xq5CjGoq6duxNykbcFFd4bFwmXbFo8SgRcKprYKKXv0hvLVQ
cjSF73RESaYtmsMJIUGyiGcuLQwkINfY9RXA5LznsPzGRFJquR8BhL9QjLO/mTnOg/EUN9FvEivW
qf2YORu75svywIl74pbjS0T2r3cwvOEfuZAWfXZYSJgcrFxGpK0MGhHhpsl9IN1YypCI0F0c9CsG
QaAp0H7x4pLr5i9Z2BbEiUvsH2ydwbByiGKK4P0w2uYe6Y8iPcptpS9of8q2oYJNm1iv7qertu1c
U4Il6KqH6SI/YdZ8haVY86YQZCYiXRm75QW82nFDjgk1L8YF/+aACs+ydI0zLXJ4sFwEU91i4f7S
9Jpgr3pfgW0802k6MiFDn+hYq7z6nNQhpgYSevYSSre1YNxxuMwwXwMwk78EboX5l56VRurXE4ai
l5sTeQRRqCFYF3mAq0J+oiq0BqNf6XD/wsfw1EILgvUf3S7yopxWeX5rLTjSWmtTTe3zl+DKXynN
6nYuYcipfnpI/KJkjFCeAHwsZgjhB5Wh6sYXPMYVB/PVmZNeYJ50ZQahl6Fdlsu3ZCTaUo/P5P7L
tWMC1xFX3/FLno9GYjnXT5cjY+B+DmW3BU+w3KbKMGpT1Y69MjWpqwg83caW/nct2zlTFOK7PyCy
4iGlvijexbOrDYuz/6/GgkegVexlSS6yNolelMSGbdEid+jPU3zezahP86nHVGD1h6nTepkD8+/n
/IlMBW3sHZ5Qa9FPxst83dIUsL+Sqg/4dzLRMvshalLdwTQGDhQoSCo11ZrfpsWTcMnwZfNcRsk/
1YegZGTnyCI7nIcSZ6RnM1BVF1U3MafZ8tGM++NVE1NLKNRwsagMQ2Hzgg82ne4F47VKF/Ay5Zyw
QH5JGBOnKKBt2aXuZAJET5aEo8fWTp87tc71dUaiJVIj8W6zOjH0PbTB2mHT2YhHun4AoMdISlD9
ndoFKNRQdIz3iajFUiEGBbklhtWRKkDS6SsNreysERsap0Wx8eDghluLUGVa5NZqdPL9Ct135tYN
uILKBgG9KYlNgDLXB7zZnGAqbYrvWxdQJr7ZNJQCtYZAE5hUlrIvKAgLoXQIcJnDVZvWclJy7K+H
gFvInakdexGYD1LrBKmI9UyCjLahdGsi4jPy0uM5HRRqPw2shzM3ds3eFSkNuA0rsu+mNo317ON9
8WSyptZ3c11RTxw4D5a6oJ0qdFrIpUp7d0cL2qoeGt3S9c0sT43WUP0+3p1PHOFoZuK9PwpgaqsT
xagzF4TV3BTwo48TtD5Ow74QB5Pol218oQtWydqVO465F8ovsrz+ctnUdhbZvpR9RFI89GsiVR1n
UlWIl6/GEFCJwErMYzUbuKWJUXkTMRYvjMKcg6vXYkhemSwWC0YwcLnou6kqBVvc2hMoz2lujgAO
hiXDpWRroBzX2gZPR6NIRJXbDpU9fejDsAraVXJlprVvE+6X33RfalZ3Oz40fT9fxemQeUHLxyus
7uz7QZTcsw/RnXCVyVnfY3BlK7Wu/e40UoD9P7RGsJQSO8Dk36s7XUxKn7AoreTVRmwjaclUi6lw
R9Q2FHM5N65opkAgrqPJ9LlSaGIYHvGM7qJJHifgq8QL2ZDfKT30UDI8yZZqYKgEihtnz+316cTu
KwCZihmO2siER6wJuA8q9FUVc6f6N2N4177YBHYtPkFBLtoU2ip2vgM0oPHPq+DbZR9WOZXxBn/M
e01x3rnDljkTqbmpffvE5cu77GbLGDAc6jSMeDoZ/SED3lKbTLQqIpIP8ALAnfo4U78XhTVLpYB8
uD2inM7bjvqeIG4J1zGA8V7dzXFPdCXvM52xSrCvHS1zeNLEF2inLobXT9xtvHPpzDCnYcJqgRzN
ACKl7B2oOvPkbsZHht9fUoMimhZpTniILvjkGugtT5jXQQXYjYVe5h4JY/qpUX07WKrkqDQY8Uew
90npjKgY36fCGSD+fxDaYMez5slqHKBJu9Mgculv5t5/Np3gyqEDbI50rwiiHrvE3wFdd+bbIRHP
tcuE0z++0i0ufvqU1MduD13wOu5WXq8+3UOF6CIFHbjOfp/paXuYD71ri4ONJo0l1FioweCUCLYI
sQS0kexti4lYO7hg26s+Rcce1o3QZcUzljEDifvdSDfIjaXOzLJlSOwiydMr5KHePul2oF6bk+Gu
kfMBlL3Xem9EQ4hFm8meEgQzlZ6uWET8gvp4hrpofuPyZqZfcTK7xvQd7PCm7U49mZFtPOOBRlyH
OqfB0uj8Y6km4SdJLR9wNrrsmzHwfwpldf8lvsdl0yeFNjAYeRCNZADaoMatz7i6e0vq4gFGyrNs
ak7eOvLwcZoBjj8gLX0MQB4wJ7FHYTs/n3cCDOdksy0WpeAzwetZal+GgMX8EJLtR5xA+Xvbt4AM
yQ3hOPXpwToXJr0PLa/g4BKA2wotQSEHsfCUO2r6SfmhbMEG36JQO8kITMzxXYLJnsnf9e5ZjVA+
b98fp2w7VV2GGYRsF2mbddsJMKhhoHDm/uPR405sM+rJyDPcyuwYNoLSFkPS6vkdqlkLlxY8qFMx
bSE9idB6w86jjvxa9r+zgWMMETUVj2XmatDG3qPWE/kOJf7r/HLtNn3hiOzVe68ecplktpLUYSud
kTcBVrIbdrrJUiO/5f7hrDirNzcPsbetd1VoouuDeqXCqcV96UpIEVNPqUSTUYsB3FmoEhiUlXOI
LcsfAOehqkiF0f8D+94IHbYa6EzI93HmF1wdR6H07V7+zdL59yHI+gCDhb7C0q3NmOtOTMX85H2P
gX+ACBTno+4QFWucfPF6gWkPml+J3/BLJqNrDWTMLr/QvCovNb2o5nwiTTUdVuMXG3niXP3S/ghh
mBZcE6ne8orWXZSi9oJGm7hhxzRGbaXoe344/8hi8HSVkVmzxpIcE29JepFvihfbF5/WJkcpTltE
eJLz/Wy2GrnkRdIh0Cwx6jaz6dZOvK6vRRyU347GVgVrHFvgBqOAoBO+vPb/duHerJH44CZi55sz
7Rs2mHNUBaY1cDxjriINJJXxdn2YyG4OsWYSrSMPxADjvD+RVYM9rcEY0hpF5r8Hln0lqzPcTH3d
BEDtQWNgJY9ZxYXN5ychGes1RVyTWM+6t9dnbPLMQVn0nDcVMNf6/PabIGU+EJdpaappXQW+jxVm
5v2NKi5yUzRnOAWFgKspRSI99eWv4YkvUmVX2Uun9TWgXPZ6B7xtK735Q/4tT4ZGB4EXBB2OkPYL
sq8xq9WZhWOsI75aN11VdL6sWF4r2wKwO5qL2Hu4aKeiFvp/yD5RvLh6Lo/udUJ0o0rWIKJgkQ5O
I8j36tBd2QD7Fq3WAtx7+t+0yqfC/EVBQ/1Hrgal2Qg7ll179C4GF7TZ7QBZpv0xE7bbobgrszeA
0BMBea5GE70ZbZNWw8bMivKmz6pYbWwEvyhl/Xb0977Lz9bwuFRZrL/u1BteYiu8QLgTLEd7w3ho
pthz4wYCG8GSkHAXPSY0aBeHLs6fQymzx5kDU+04WJu+zdJl6hIYLR3iSERT0OWwk+x9ENVw8XNj
xAc8o+XRacgqFldzXcIqs4VagZrkvCWUcuSH36ZcRworVW2cEFQ9HuB7J+5Caa9tVSCxt5lHP9ZB
tjk9wSHxqxUx/6cVwuVO3k4tpp2IwsEdryt8Qd4ixfgX33cWbZysVLEMRUmPAB2600C5hail/wVc
gCYwWlauuVK6Px+9ODNEa4MFmpoLTv8hVDZCnQdFvmE8hv2rfNPB4A7a7z+wwJpepEULqq03y6Hq
lI4k0nIB/IJIzt3jIlMk2A2LjzVbJdFl9bIOnFFcgG450NeLmHaEONHjJpK1LCMdZWx+8vGlMYrn
jfV96FfdE6go9Gp/pnTyCiwZot+unqdWwQ40uY9Pn2pwX1/mk0iX2LDtIMw2BNb2XDqSi5KRXGju
3Qv/1nFJhIpqg7j7gjScrNovvCxgjiiIfte+EmX3bnrDizytOeYzVBGQuAwXkp+sfg1XRJykLiZe
hWH1vuds1blP4iCe6m3z+Z8u3xtzjZc9nqgFM5zm+XB8iVcs7eCV0z5LJxwux/3gyihlASCUYzXF
ZYN9fDFOhaghH/tPF36s0utvhRnOZWNGcDK7tJDo0Oj73suOUPDMQM6QvVkjF1c48afeNoA9e9xw
Sw1xRLXq50XgBPi0tNYBzx5tKxfSlG2EljUXrHK0+5jO1IL+KuWgNYmzedZm19lVpZnOHGDK38gX
Y7G2Ue+k7LATUdL+eXygo3mksXJs37XYTqcD2rv4cj+LTWUz/EP3EFCwSQQeyF//s759y9UGSw2D
rIo6tS21NPuCn7tBFHKVfJjyQq/vtBWz46WSyMDqkiLJ8fiah7i9XuuegUBlAroNxGe2hMMdOh2J
3wQFeXfRPya3Qae6VW1FW+JYAlROvKVWzbyVG50AZYYD91U3At4Rj190dN6qNDz/lqBk77wKohJm
9JmgWkFdth/h0trq3PxZumJSWJ0tzjsZHHoOtzup8HYo5QyFw9fC1HlFDqrYr19ETTA92oLBsF8e
Zm2OSxKme9LzGT9OTGeGX0wRlmVh2x5d2ploFnQI+MlxIoPbUBYhPHCMtSNA8yc+Jo00FaMQ5/fD
wSLGGpi8q+zYqkKuXxe9x7Kcmu5Rrx0D0HGdR8/I0HJpks7ks5oma8RYxVw/JhzyR5ky4htZ4lgs
w4l5Xxv2FCbdQM7FQ+mV//PwGbMc9IyXTSYeCmQ4an/w7TwQYEjSEF7cNw3WUUX88Ut/kMh3VHgK
aaU835KZwZuW+omWLPEL27TARNjibaFtUWKp/DAtuuyTA8xSudnEmPPuwB3VPLwQucvI6O9GqRMy
fnIgdYID0XTw8mXmokVwZYvCQVZDH17RBfej2cHIHdSNGQ0OACdZIs9DE/gY8yKgjYy/gt4gWNnf
tkKYNAbGMyHsAdzPf3eR1/EwzfEyIdASO8crG8c7H+jE3gsMdZ69XzTJnByNb4y/3BKnJ68fXiw8
+52CgUp/Nr7KbLOhKudzZea0U4968uVYEEp+ZqeMh0G7n5Jg6kZ9lBWhUucZrwIO2d9gMEIF+Qp8
JW+f1V/bEt2Qre8bCxw115kroDXrVJw0emvsRB9eDY5+U52xbMwOlG4V7DCH0ZIv/n2rzkvNCWuV
FNRr8S6Hg7SWjmkljiMER19WfDmJ7Xa4BQpP/bnGejV3XT5P4wbzsd8FRUVAL7WVOHe6cMGsSCHe
CqXHHNa/usbxIpyb8ey4rpIb2bXHPc1WJr9ml9NNbx1ipEon6e3VAliHL4HueI14G3TqAtKRLR8x
d+hgULagV+0uRBesn38DqM9w+2JMOjzTp8scFUAQdQDfD012FTqy38EVNWKHYWGYQMyjBlhyDmBo
HP2oHseBn4ATgpW2AtLIySPrdfjV3Xrz/CV8zw4uFSfEgixFDxI6lRC0Y/hnv6mc8qTWvVHSuxbY
RTtoO86BqGjArWPJKwwNyALyQ0fBtSMSswddGdvcdtnyqWbkJPlvAXX6qzSk4ai/8josGtz2bzVD
4b/QCZIADHUfeHXqpOCZJmrQ4lwE4wIRxZgH9uPOPv3aYga7nEw+p96ujfdh1X7xy9eiVphOcc/I
Ft1oWPJQ23Vx4KVjOkMHt6jRslShZUR3E8WPILQPnjggFy8j5xFVeBUfo1hFAaKXG/qAcKeKfrqj
L79vCMVDPIsn7AKQDZZgDeU+QNguOtoy3cPo2+yukeZy72SOYjMHWSKFRTvTHk1SrUy6ju6rhQnO
UNAaA6D6H3AP78vxX0gYj0Ye0myffcrscvlEeD/qJdD/fb7HPdQMWhMOzLiDeQjoYZxw3aD9QnmO
KN7f9+JwU/fo764YRCYhSHD8IxXdP5c/MaOYjKR3i60XDQaRzouGWdD/Qt+3+LMHEVAQgC6vZKsk
gEyVIvuyYan0g2X9oREACNsj48rUmLjOWSSidk+tMiv8Qst/CuR0t8+KYdgiuApkIWK/M/iVhEic
gUazXJViL4p8sz3JKFmtBS46wsuPfsZlgDNc3ibU+PU9i0eoGWxVj9kebRuvhA2OVKWNxrvTMpP9
r5PMr4vdd0vwg+VkFAO2vx+ycvp+Cz85KJ7B6aBI4mWHWiKphWnjPYA8vRSHtMi5IXy6G2rDTS5R
SygQL8FVIBdA2LhHHZWDQ7CsN4OWAmdaF+fS9JaNUYF1b5A67gGsK7eJC/o4qFPmEFMmOqPslKG8
NARzbuRvbGeq04/EWI4B/wgs6Q3qqxqQpLEYceoG8Q2jNd+l052YDVaxXlbvdVV05HmlMUdwSsVp
vWZk8G/MykKLLEOI9l/TNkknN0GtgLG+NAY0oyVvyg4ETp4fbcxu+rmZF4TAghB37zMVI3nNiheh
1drmVE+oYLkqZ9eNVEMCmIT8plgtlK2R3JDQdgTdAavmNR8YD834WLwl0gOTYGhlKguRa16USc4r
yWPynELcAArXkqsTJ3v+y1hreRJhw/qJAW6P449+ZuaAVmECtfjvve/sjIKxPIky2z1yXzaxMLdf
qhLG7nZIytS1cUu3n+0s8NoFhXCKPAqQVBbK1I6M2UEjQJGNVjxl0h4j7K393KS+BHLHA+AROAlO
T/XngBpnQZ1HMGSZLuGopTN8VPx1vtGzxC1nMoy+mCY1oye4Is5pKL6SDCuJiQ3GtyE+bp8m6ocN
nZMr0f0SjC3Cz6PeOEaDOdut4YW9DPOVlqJa55RblszhsJA43BpiRUaCkDbtDGFkuBG0O1gAXkSu
gcVdcCJjxk3aVD7fBaSXCDY/weIamgsxJxEFwtzZcoTLxQ2rABn1/aDXTonkv8mehGNx22LH0xvR
twuXOKeJEy5x9RbUOMeQCpKkpeYaugu/o2RecCGp1VW6T0vTf+zEiGOuJMDcB0doK/pDggTDFtDy
+k+o8tNyktDBX/Yr+KWZVOM6wb/GIrhsJ8eYDLnd5PHPnKqq9XUOF8IMfa2KeMRXtGFGMF469tdl
umYHKq9GzgCBcxx4rcKDKNCaUONeF6RsGvu6njyEzrs4CWUseXNZwm1o7px9FyG4GiASEqdFrNFq
A5hFailz/KIwGlUuvgG6aZLzSCcEqqOd+f+yZS5uPRWk00BN4OOmTjDwGtyDS6NuGVC5K7V1mgX1
nXkVc+xrjbSOgDrlL/8/LRKT/q2rsiYvLSO7Z9+7B9tbH1PXi/NidQE3Z101u0UNZm5dhNIAGdGe
IotGHXfb2vkOkAb3JCYrY/c/nW8x7HSbU6TSOGNoqtV6qcXLwQYoTQ+Ds9E+LTLC7XX8sc6+fHUj
NjnnkpwVaC13/7defaI86KJi2yxURyx68L8xqD20N2r2C0zeAcfIzZxg+gQGedfPb55rbm3FnvnF
b6AJRPybx65Vm1MXeCY+Tz0Z6bVbbj3XHiEpeeKdlV5bjglOUjPEQpCTSCDPZp4eW/yJUPATCkC0
vCpFa/mP7af7fwYVXPpFdLYITRTsvmjnrXVYYut67Fe2iBX+/flTvKYYkIe4G+hhpWUU1iT2tk4g
V+i02iO0F12ewGYStihq0dFYgVbYp+PJGEIjkA0QVQeCsNUX2r37m37C1Apdhf8wQ1E8dtGQhtHA
rToDl0i2+lv3aW2tC0dizIEGQX1ATrYknR2b9Vilp9kCgWPGfX2VwnCR6LxBx9EYhAyTsfjZD/ZT
nRRHMBB2oloGOFTTdQ5GbLDOA6737TibKd8NJI7f8eFasQgY2p/wPVYOS/kvpzzMVB6C/IB3Pa8Z
6sH9GJcQ+u+CoE051AltOgcwHVyjC9gPYo9BqzDr558X2E9AvgNtYd5CCknxR0J0HyhdDk44XN58
7BS7FvZtF3Pqqnko5/uDz2YnMFuCq3P04HuURVLQhIwriStfJeJ9Idg881rYFfFHxY/FPGjdoLV1
fT9BP41GI421eX+r0yEzJjBFccEU8nVqTA12tVgz2ZnQNlsMVJzb7r5zqgpkBJ5sQ3gb3A93flw9
E3U2H8yVZDokGWkGWuayywyC3TtxEQU3Z/lH8a1OYr94ql1Y+XdAfIJvaluOig0r2wE1weTYK/K0
20X2ose4D4kt3676FY3Qo1fzu9OjvsWdO35dnJZ+6nR/5JEES44JD2fsC4nQbXE4ob1pkNDxNpVP
vrxTlj7zeIN19LcxdDn9y+Ir6ybw7CioT/wunIL1trdlxKiVcluj9Mm3kN+GA4gxoihemj5Oqkla
i3VEUGtuleZhXBSnNM/PBKR1SYQqf8cWZDVXMZWkjN86MiP9KCTaCy1PdFWHM4DeEhqolhGZBXet
4trI60kKkG5haBYYSlBUuvIfonrr7pF+9jPZir/GufLe1hPr85bXX8rVkDXaVLG/qpuskDDpHHsV
wfghqz6he47Trh1nVRB7FyWGLfA0GbGNaPTgrnrUnNp3SE1PS/ZRQwBv+GqsPYiOFiWYaGUwF0zE
uP5Uz1e6rNfiw1NyptPbBVcHMaW4uLB661ocU49pFL4aSX8G2GrxAs6ISXUjSBgymSYMbPP2qzc7
Y+7utnoYFnLbgoEw7ULljUQWkv6IEq91l1CpYVM7lZ9l8ZFwvyvlwj4wccdHObzp/yBZ/bOsLLmy
y82fQlrhgRTVOESDQDvsKgHVOaWwJpuQo9beUhPVUBbs/Vjpb2uC4JnMQ4n/FMwzZFH+MOmATxb6
k4uH3wNIqO4Ma9JktJfUEV8ppoZLn0XNkbSazZcTHbSSw2Qgiz6o6XYPGl/bBovZ+vndx0Rm6CV2
Uv/Uj6fcuig9HxyA80dwleBgNlpTzPdvrr4DIv7R+ZpaH3uYIq/dV+FawT06Kz+fbtgNZ44A3AD1
/Qj77CX4HJiGvdsVXZzuWS5EAjqrG7ILhx3pdqHp9drS6tFHmSH5mJa+02tU9gXjJoZUos13yAPN
4RfRVSKvGxyr6HEglqKaZA4/R5GPZuP6MyGdhlHPRzFiPnkJ4+QfubXfth0quvbeC2RfOiYJrWlF
JfjwEJNAVB/YQq8EOJv/vHJra+RhrEAH3wvy6SrFShqBfcQTjdDJ4uvsPP2NAzT+WwxRxUdgL7+/
qjaco19Kv/OipnLLxA3KHGCxiEu4x2qYvUzgKPMSQUdVX9I2rsg3w+jjawcjFSgOUWwcYbBKf/nm
ZWT5tmp2ml9ml3nKh9OBiqmTKg+o7uDCeTPYrw3Y3o6u02nTRFNCrBXmvbcyFKBYH8+dDzuc1v9K
i+r0AzN37+qk124HUxc/Ls7rV44dDG1kRPa6Vpb5Y9TE/dxfyPaJuhmPJWchl5/xNGeT9QjVD9L+
EKtguvnke0LpsSkQPaHwPwatZTLS4jasv163K2HyG5B4Yvm1nKB+PbcBk12AAanAAPsMhd4cDLRr
33OQ7riu6xDOUdfwIYRBlGKxT/FSiouVdVXTly+ft52wzs9wG6V5lwiiHle8a181V7qYJSiU252L
1GOq+t4PNIzgvpPYly18UhNpV9jRTVWEW1H3xRDXy7UA+7wVSYqGkxc4peUvvDZplFjKveMpOMVK
N3+HNnFtJCy1WnvUJfjI7eVLj0bM5fVLNMFc9UDLwm9PU9JBC9FhB1SauqBqhuqQHJ/Pg91P8Vzk
HdOVFCeUnfj11Hc2oLNx63e8yUT5I9EF6IToeVF/FKlbxvAEqRo3V2uYhXyirc3we/Bi0/TL03um
iYWSfe2RvS55q+GCg3RA1c5Dz8Ygrrb6bMMpdYk1kRZLjIuw6XLxfyMLVfIKYtXGzQN990U0+xfd
HaM/wlUU7ATqAb2OS5a94sMIbmJHknHapQ1sObtKib9YIJjzrSwnBh0kAp3qFDsiJ75BAlcUsvzg
yy/rRYfRzUbN6XR8fcrFycvZgiSHCtBQnrUakwBpsAE4r4fHWobEMNjhyE4zoRUTHNEAyAifagch
jF44aZu0MZbh2eExvXsSftPd1cB45FSBJg3e04UEw1YOJFw+4C82xJAGGUzHqQ53gs0fGUEoLHSv
SGl5tWEcVQKS60YvfcaYiqC//5sCvCT+1tLwtCgslB9j1uGiBr6LuzVRHT+XPLtzEUIfAmDTsb1u
4KvTuRZW2OXItUa4I5FrPqKJmAy0aghkvZxhLLt4XwByb0IvpYGcTf2KH6LOyUfIsfNiwCN4Hq6W
tGqYKoQYR86BRhsLDKCioB5AMhcjAMM67v6llEMr4kusQj1zYmEFCpRggEFmvq53JAyYN7BRFXUL
n4l/wcH/L7dZL4CTz1N3bgepOZDFhRh48TEVE7T/gnZPOBXf0Ni6MH+DpeJDn4bSFrCSm5BYbeJD
gcJP/hwDGQdoXZTA8s0jnYHQlMsoftK4FIciJFB/AP9mlaTq+LO3WhgTWVVwT+v+Z7D02OWtf8mF
J5knfxoY0Xjw+1K4ty/UqKnq9Jqm+XFHX2XIUOm89zmZQiZVigm3NAcCEqFnLgA+PLQRd0VNd1h3
hqHis0BpOqS3WUN8Xs0pGGYqiWTdIaUGr/pLAwelhaOLu7IDyno514v+zy6cXXK/dWe72J3OUays
6CWkI/F5Gy+UXaaH7ge1EkIZ3hSxjBraP2y8L6J/aO0JrBJlrWdf9gvnRakcYIoAbQZLLUVqXiJu
fQ9iH43nmDDR6rylWa5r+f8x2xZz+V2+kiy5MWAXKt9ZP42oz+YFMlsYD/kXv1cO+6ZQYINc0bDf
8mKdkIXtRpAjs/HpO5WPNOIp8SJG9YQerrLAsjF65CbzOmgyVjO3tJoQpqHmv613xwlvSNsdgzcV
OgK9QbO8LGPhDLz3MIm24aR82VM/Tl9xWpacgy0k1ag73OPcoQMoSXSUGkljyhzkOj+piRttdhWZ
rMpRNJlf5oHSszgz+2Fp70EowaHzFLglAkcYATZgXLfIwZS0lt+P025eSEIZC+HO3hdDrE5IfZ5p
SecLy4c4U22FW3PB3Vkf/ruZ0DqKdNWWw6/4SeQnTvfXJWuttBbp2gyY1M/1TClL/dTGPkDKgwqb
AHFROf68qyrEtQ8AJ2CzlMtNNyRZz9AYa49DRDW/ONWKGVxhpsWrIcORETILru77OcJog+jJwH3Z
oekOSLmu8QwmCpAcIOzRu+GFKWYu8PjzEY07HJd03wME/xmjdn7wj07Ma9NmKW7Xz+jXlE1b56cO
lKFIcsVBkGfFYjHKHO0JjfmLzJqxa95L76cHqLAvUyRafNhJ8PUBeRBuLC8fqnUf458JXsPIOE5y
Wpkho3kEza80WWxzb2jC2ey2YdKyNVJ3bMto75d4pXkITbCH7Vhx+dY0LGakeapvt82L1WKyX1SI
btKmRnY0gjBO03q0B0hwlOArCs5XKjg8NhnpQd0ZS24Jor0WSM/Cgx8GzeTEE5hWK2fnYvUdUJ4g
fndXRE83+zYuVEWbyahmlowppoaqBshSr29eC75eMpIH9vMldepv41LjJ86XDG+L4pbT7Zv13FPh
4ap+9Uqy4aq2qAJwX+TnvIIjxuixsW+G7EAPmeWRrwVlWcBro2uZYWsfMxPEYohEwVzWo3kvx6id
5riBfTw1JoCzEw4peW1z7RA0tqKbvpE0O+OTM9HbeMIVbpXBfl2DyPUc5uoB7aILunpkh3LHBY9H
t3DbOYrMdbCfw8R8wpDJvV8sgI+V6qGxcJEJwAhkFAR13RF4Or14pyKxo+v6b5AzZsRn68c29LHa
3NH+V9pVxL0+M2Kq9CTsW8F4JoXrefC4c8Ou6+HnWtdfnW2eiYLDrqnLjSOxsbnXTrSedGSEd/zm
wzLtxEirzXE3qYWtpYfQ4fsjNQAtUhAAyJNJ//QBZXSI20/R/FvxJJY6t9h+v4MPVwxp/sF9KxlK
QVVr8txllaMMkCPftJPELXpiO85++hq5Uv4AgWFUiACKBRm4wFGi9Zun4no+LVEeeskXcqkU3Nfp
zkANLIXZ6lpBh4Y47Kw3shZQ811N957zGYuqpn4P9Id3jtFjWAwelFdk7gWjMpD/0NDpDY02xCwu
+zet0Uw/3+HIDxhNV6e23WiPPVZh0qERrsFylS3vlR6kuhg+9OOVkbgyHecSrjTPppDnsAUK7Kkn
8kNDG0vXevgqlhqS3To6Z+bKm3pqVhApYGpqU7rhIkNXea76BTcnX7oQXFFoJ555Hs2H/piKInvN
UFMMB6SCN5owPDWw8P6ai3kQ6mLMQFeWctzBJy0oduAiNLklKoMkSgjra57wEGQngZsAOI5n7pTy
Qa2yHLXQA0Q8QYkvko2iWDtrpuDe4gKzwutspJfEO3K43hmnoo8s0iCK1MvmOBrbUe9VoS550yrC
OkuSzo0YEJt+FpnPIPAT04TrXJSKkhw6keQ/O7YGSyQRxFrBgEQI6hnMtri7slgJ58JV+iYTbNlD
At/k8pLGWkzM5BJm4gihEFqQK+A7xnPWTOvRGxn4ihvpFzXuYUCIBxfv+/Apa8h6rOZWH9aEcXpB
f1tqlaA5ztSVvrTQss4Wl0p54kz7yzfOQ1LmvYZm1uOffIOOCab7SPEN9Vll1fhZMlCih0pvDBeO
feIXwyeT6Rv1/DaBsaylk9i8GHh4eq7x7jQQcHlxfAVPoZe7lgzefyljGmD3DUz0qkLsjealsvQp
tVv33XpThhfUWXaMkYO34eaed4bgQjnHD0NE/Y9W/pxf0EhWnhP9F51qYG7hLfjrmTMlmzV1hcew
1q1lefZSnA75GlCYH1RuYpXVXUF/rjTcjWu+Mg0yeKKpTS4iY0XFF2f0pTU2HkDHd7em7oiXRDFq
bQyshY7cRIB4ZP4LszqbhERrieiDwC+8xjZs9HtOWSxRtlMt2KgDkp8joyO5Xw35+ym4zgi4soop
54Bdqzybe7FN+DQYhIy7I9p6ehVJLo70nmnrGCRS8ahlcahHSpJ7eM9oaCo68SGNJQPo2HEorZDZ
KyNAqod3Oqmx1BSbFSLuxdBspOOb9/B+sZ5gONfcBA/TcpPF43sJ9JTPKcSOZYGqyrpjP0NEqb0Y
3w2O7wVrYUPGMcMU8/VIztIdWC+AVao4L2EOx2Cd5OwITbSb/6z2z0PqvzcDYoJVlY6FKwyQ39xu
/434EmOXSOex+YjNQzYaCk2foRjJo7NmDYngBonVrD+BC3GyaBsA/2f8fZpEQWOd2sk1Nfb/z1LU
1txHYB+ldkRrU87phlndzaIeL/1XbLdmqqUySvmmt1Or++fVIGIcNmQmZ4aGK32iRzTa+vyWPppc
lL3Ep+PZXQe4xpmFzooVnxlFZ/lZoynGmw18SK8tqf2DmucnqvXMKpOpJGgW1UWBe+RXyDfIy7tK
70hex34rFbh/d7vOBbQiiOLsywRbMyfoipbazx1YaWAnG2pCwHPgghJBHzdloJ/AIolEpqOCk/Vi
vkZ2HLdZqIGTqAhTKZxRIt6ocNsOdVbJEP0TkeVogDywPTYDACg654uOmgc3nnT2TdnrF27Zr6KS
0UibOU8IrekJszcGvBgCVyU5RwK34gsHiPj3pZyA2b5acxkiOq+EbZ2HBf5yAfal7KyKRogeVYVV
8PaOl3iukhGdlxvCGnyEPpUGV+ELUg0vc5L/2Tk4oeJtk9L3hp+7MdpucOfcQjdJxbRZPFlpz/Sw
8+WK7Z27uJNdzoaAz8zCKgg9E8fuMk6pUUbPUMci9LFIX8ebvXbCim41zpSK6OjlLqZ/w3FwAO5R
iGHWsBIwq8sM5A7zgqZCw0k9ZhN8hkb19VYUfFlymRa3bgoeY+lNhyX09X8tn4OiekIdQbHW6OvQ
EKQPKXdYAhoMcR/+GLxPyjjipMvg8s0+nWE3fBqWrst1R55mrCs7YXHrqr/z64JZaOCco3h1de9f
0n4/jBMvA9iSJiewS9xgyCRWettzGdhtJyBsOfemDzKOLh9Uaio8Elfvugruo1u7il+kl+dQjM40
S6fRAqiPxG+5wnGySKxNvLdG5CzYQyQi5HhRmKPHS9Gi6QwNdkQmpME9dn5Ovy4zIn0yP58fRZ88
vqFBzBgewk7B4ktM7gb5OE63Vu8Dl/xbgO12kYpVoFGDQuKm/7ghmG9WH1GW8kfP1SytSUpi7PWG
3+6Qf287QUJGpwX4fUyptn+xOCa9adZasc5aRUzYtPTPpLi2mzjqBW2uMLsyRm19qW82ebicth8Z
0BNGyF0WbpUsXl+73qwecvu7v7vZF+uziPpCnnjA1KQiaDw9C3ytZBswDM/opR2+Vay0fiuPafvy
6wG6pbk6/R1rUC0nQTLO9cR5aheXg7/XQj+i5cfrDU8rou3na5XtCj0rZy6yrRYh+h4rf+HSTnjt
Zlea4S4+m8gXh3oWCoXPlAOB53bmI92q8uSxwgquBbPAY47wkgEm3pITLof0wraSUWFsZRjgAEp4
UsapvLNgb4naN8pFsfLFAYRSMHwsulkRPCQXkdS/cTYtYO2/yNzI+0Q0oZ/peLVta72OwDaqLKtD
pcQ1PRMQ1CFwDlkGo/Avk6GM4+IJeKR6tCBsRpjPIEdGGeClMc8z5HpXoH43H6u/13nvHUDNryOw
tbCkw//7KdCinxAP/m/PfkS1ijmcf+F+xK+DRRLkQNTvEccFJmu6cF1c5oVIUZ2UfERplOm1278m
j5nz6XSrEXk54v1vLeyF+pqUciNzUW6kixUUwbcFf+raiK3M7Z8gKCoM1GQoiogIHJX3HX19sN/G
Iq+GjfzBISrxacuBfex7UFZNMZABS5S8fY03jjOjiOAzcypxD0UBBaC9DEkpPBJ8CbtFpbdd0o5N
dJbcbUybRi50wIBS0QBkRv0RX1Y8GgMmpBwY3PaDKLon+f02mipgI+/VtKmMNzGzNHGB2UZcUzFO
7652O3iKuSR/t/DsWEpRevvjhpLJIGFnTvopaUPcyRpPDjcXwU0eZqcqzofx1J8okix8HNi/9Aia
OCLzHDLvlyOyDNtFQxy3iyjtkngRTonc3U9QrQOe9S/IIl/6hVb55q5hrk8MQouPonvgUDGbLS5l
EPsJpOIk22ckAScFjbOgvPKL1wVGVc7ucTtsKf04yeNcfD33jgD06PAYfkKdNvwJjivp41xVd009
WKPSqjnFAMQyAnDHezjb9SBUD3+CgPvNtkG7CRfKxyAOBWDxsYA/ow3QXPi3ragQFvDmjLBBAZv3
vQwKxcw9dbz7o6eA1uMztLI1oBkIg3kynBADITpUJ3C2sWAPiH0u3S4TZdKBnRAjHWTDHc66A9Jx
OxiRKQlguYZuTTWIM2X93Sxjm5Q/eMIkn1tPBl3mGHPifBo9oGNCIvG1zaPRdmwWuSXjr6vxShvT
lwqNASY72kCnaO1ojB0qQlY7wa25CJxqzZB37ITKwdSpzQoamrigBNq0MY76juGkAXmL99iEImot
vSGJAAWt/g2Gb3lGh9nBh8p5WzBi5P2XDz+W10YyMcHuDKeJ6LQw/GA89tthAS+BH8mIQNOcG7Nr
ooyhCKSEzhQnY1hYkZ9UcU5lQMgzkAs7GkPRc+aVTbW7KVK+dOnfD2K7RwOyKMiWnJ7NYLVB4v7N
w1esK2Rfvc0G7GywmzqLDvQGqiIP39A0v/9hmppBYFm221ysWjkuskIgk30bXifQbV7AoM47cgEd
opV+24YlVDE1bB6LIoGD2vNJU5uvJSvPLriU4WUay0P6EEL9FiWiCNzro1/9+Y6YN7El1aB+gesV
+GJpun23swOPHi2izYIb+qvuGAxkKp+2LV8CF6TxiG1NP9ydRo7P67RyYG+/VZQ+LfqhkekEnpnI
xuQs0xBfiAjOhXoA9seHSx/B8Cdo5vk+T3eP52ed4NxqWxxqdicSb3gGNXiNOzRpU09RU8em/aS/
4EBdAOjaIoTBVki923vPTzVgEXWvJJOiVf1NmikqtXJ+3stOuzqFnte5GYWH/OfAgFX9lKeKTg7D
wWo5c7OMoobqGnOYwf74uCK6gD3RWIE4nvl52QUya2VsMeUxmuL6mce1YzerbPEUTiGvLnjutJVO
Ezj3ZEpWXbxB8aLnuyQuIwsvIYOBH9wCAvtaa3MQ2J83+TV0hHOZxXpUuKcr11QYF81xvgb3hbOP
owkL/ayb6alC0kmZDuBg4O9vVC19y1UAJHwTN4C1wdxk0GOQ0hMfP99AktLHlyhzJJ/9Kh5rJz0m
8WU52budm9cTM10S5Qq+1BBBV11x+aIQRngQUu49vqNU+H1T510r54tjSUCmqihcHDkS8932ZmTq
TdkucDIuV5GTaY9S+PYJPuz8/xvoA8gyiWxzmBMp/BL5UVpeMgd0IGnbDiNOtvv4au/5gtaKqxo2
AGbOYarAC1uu1nmUXMvCpH5t20qhW3fpBMwmZCEtEO9cT6TILOkfjJJBg3zgE96mJZwRLQtbO0g8
hAy6xCD6Lz0/0mHP7IMJ6JkPPj1YPNdkVGV8ILOjTcKGC3KCpQ7MOWPB9Be2vUCO5SoALUXZTcHh
xlrDI6BZw9BVKn2frkAxpICAfAjLiHqZHwQ2luWIxiBTZEhZIs+DO7iaybu6AJ0icPYELiWCe+g0
22yhIRF7eABH86oSesVtpkgtZeM5rplNkiddY5ylYUaU4PdqjGjnWZ88d3VW775hvdI5tXeC3zsi
gcGBDoZKPjVyyZG4z06Kkv2ydIQHRqmDFyjoXD1DqG10q3mCh5OIGq9Z12UsCtE0YRWo3A7IEknu
KvmISpcPXx2bO3hyCN8rmdegCtUKVzzBDnE0Tf6GZVkqyLXHqHM6hPzDwRSBIUX3Sk75LLwrUuLd
3Rc0kRLQrexLvtHBSUtzJ0reSxw2SJQ2QDeDBZmRxaRIgLfP75AeAr/zfjWfeH1DrjiA7qzKHoIn
PhXBo9EZNGV81I+VxkPUm5+1tsL3dYqFAQGEGXooH71DhvhIlNtNG3XtFSlA78qSvR/o6TzdL4DR
9YlP28Jxu1fI8UXLy1w/3Q7c/ZLin3lPaFlvyGjQLa7+sMG7rV2t+M2GSdBbBzEm5iHyGvgXmSr2
8qyuqFjtC7sT/8zmE6vwj27mwNKRwgAq+EjJ/iGgXhbAB16qyqYdz+MKJrs40Y2RDBVuSkj7MIS9
o5HuHVquKJkyjM20Gwns2LUKE/mZykh1uNExPfg/tvL30NObUfUlFPnjn8VdROJAAFts6Fr8zzat
bVyGlGTLMi97CitxSp4j/+2t0IeliAvX+5mhFSVdjfbj7XZcMTgCWPv+Wyrb2rj2n+zb94salppu
83sY8DcNADODQzRZ4tZClyS2leIQSAWr3w3CshfKH2ffXU1g/IgmYVfzgKS4h5iMAEEzBtrlSXE2
7T+AOXr9DarqsWYH7Af3EcpdyYI5Zjo2zYuwtQPZji8UclNf6/TSjHhqo+LNVTml22/bqLTxeEkL
u+/nJ9zQAmk5GM+UbDVH/2o6XcO0jaUa6XBnwhO9zBM8bdV1YBsiZa8yReGlPx6Z0a2CwLLjTe5C
4qO8LNRB1wkgYlk1SWr5+z0ToDwqkSuhNcTpqTHMERVyNLPMaMW81BsXbtlBimvpA/tqFAM/cvNy
sFkhYpl3VW0TFc5K2SN7hT8I+5vRM+y0U260w0BxmduZG70qBJ0GZ7GbG21CbvcGTNEVgF+sGELI
wV5cCAi71n4JQ44jSx1XmQP3HhNNeb2qc1puUSgKLwDntIvjsRAZZxxI1O4EIncUKDxRm+SS+VyP
uob4tpCD3iJz6fXJ7FXffL2VdlRi2tiGJbGo5BKUIYTS+XgVZ7bjAY796NaWPlC7VBYDjSFXjOrW
GvyHn78btPtdpqRPX8z2y8yRwX1ZDYsGVCckKNDNloX3JL7hWGJPwP3/45FtXzHL0qprokLq52lH
RiRDG9hwNDoQwxDiiCV16iFEHRT7tnawRSCmiBizW7G2nidmFSaL/lBbfOqZtp+hYWJClzyMsdVD
KJ5X7JzH/KFp34+0OpWKiaMjMhdVuNSiMhUDPYiSAzSbadZOSqHYZ4DNiDtKfpDKQ/h2A2+Bf89Z
w24OCNp5mmyvR2zgMVQesqyzqInG28V9Hl0Odqdm4woy4zD1AZJ3kjUtYGPpRZn3arFfVCjpMGEz
tr8j9yEp/OvKeyrC8fV+cEg1XWF7SvYXiMMKN/fWpSFmElFwA9mQQZ/E4iE+q5X2sF+2jj6mQBXx
bsGqtSI5RnBxhwiIlI2hXQf2hr5JjVOdViJEyzgAEj8FIJ+cwiWY2wpYPsfXOJPN3t36ZyRPvQH6
stlxuSEMjQa2tvcamaKW7DBe8hfq9q877HSinmWW8IaW5QobUUaMC5jTvnM669PGpNjJrVJpMl5X
CEttGX90Qwyzf58mdu7X85NUqEXk9waRhUOcpUZtNz9p3j4PDX7MAaVVu2j1ZJtkrr8Faely4JgU
uIbbrqOVWRSNBnofe8Vnypn+t2r/C39Ju299bri6+hXQd1zhP3XT4xgLdHgThv7KMSvlpBYzvaWS
OQ/rszzG7SESB0r1EP9C8R0FKR4nllxfF8daxvP49YWV+Tz8b5l+z6Q0nKRsBb3x6Fh0K4kLUmn7
6aEc2tztWrEP5Y7xeb4gCWixqX0DukB4eQDI0RPjqTFqkOcYtdP/1+q954RGoNCTuunN1LGaJiyJ
UGJX1HGdaAi1iLdnoMl85NEvul58dCMNmCBEHqZTOmTX9k3GNjVM4mKcEjMW63BiE6XXgdV42G/+
lPLcShTKN1hI6lq8KG6s4H+CznZSoTZGedeM8Eeg0GHaQJePZSUvt6dlsbAJnZNpOKkloV1C7Fzo
qPXwhivQe2WTiP82vt4eBDs/AE9D9oLzF0Oc+nKy6jjy0tndAGcxPqvhpHHfCWGqoLgae2KQKY7m
QvBkuckQJ4LUE0L2zVYXkP1h86ySGjD0L4MZVW5rmpFg3tQxw3Eqew4WgY1860PT4S6kpVnlTyAw
j7GJdYWiuXqfFAOoptK3miZ3kPZg1VT3bLKYMLjgRcuYWlKOqLzK1CY77AF5CZvCLY2UCtZBVUCy
rcNmSpVd+jixIYqym74xjGVQ+7bTL0rbmUOBfKaWo4iSj1urmzJD//CWkPGpb7SCoWS0iAqFzm4R
LFxEa06eRzrvm3vhup4wq5hV/vNoaJjrEd57mS3GLhVe5alaPueFe9MuPPGVs7lIIv71O1zwqXOd
tpRwV8d1lslSdJf7Zi/xH9h6zG5viyS8IjNPLdM+DifxwAmO9YvPdcGSNTVMSTfMqFO7ZKY1FmeU
ILB0s5A29ZBR+ZCVTM+dkt9iVD6ynqujyotb5EVGPTwZOCHObgH7M4kdLGV4+Ah2qEJRg5Ebnt6v
YIJM/gXpgWwjVhH51+itONNOhGH3XV6QjMiuNV/QCi5x2rw8/4mxxZ5K2zMUpRS0PNmOe7TDkaqB
8DNQ71yg7y0voZsE4oxoBD0qUWvdO6rBOo3GWmLSb7pWPLKxHpREt27hJ2EgRJqUgNA3RznLM7+a
bNgJHaqsYmU2aNXeBlgY3WtWf8X06NSB6QnP16ukyc06DmosDzYgY21JNG0gaOymlafMhB9DOkHL
MY4K/jR8HRRIPEeBNQSVfr/wtEL3WohaVLZbXiLaarTI1TtFbaIEtF34s+6qkIOPBy4cGmfzTrQz
DI/GlD5K7nnJPunvrOaf1l47hewiijwr7x0/VxZJIEPVYkvYyV2GBESCCHLdS6jdytTaxvqDrPzw
eQE71cRRZmyWA9BXASdTpANxXIS/35PEIL7QYSl2AIeH+FM3nBTekZ7TTl0Nt5RYc1oBiexKqW5f
7KBzBleulqtXaHty43/ROQqCc0FzQd6Tmlxw51kGzkk2eGKCQIT1tlc7N55DzP95aFahpfkCnAXb
noEWA78dQD7FdjZkgMLdE3E+gECWuLGcuTtIm1LMlU89hpJwGBV+QHu8ZZ2EjyZ91N44WDB9H03b
o9cUd5i9P5LDFXsxlLoE2wxr6Fn5/cztSD3whaV9R37uxw2BANmPO4PrKnjlX4RTjWotzjNKc0v3
visl84QAYxHYcOcxap9px0fC8miGXLrFO7jIFSZ24VWXKlq2mNYpRkLORby2NjnNCfFecb5RanIg
gSQmgUgT5gh6q6Mf6uRRl3LPgrbf8au+KIEr+QEpy/wh1E+mrFDn6K9JfJ0L1tFWHFSfY3aH6loN
DOQWEuortOyoe5Gtn5PO57Dzhfza2TzoXqlGWFS/MW/8ovP4iZqm1jqF1lzfCUIwwiCb9aTmF8ip
mnSHoiwugOjWc0BgPqXwXZIfXKeDDoDgfY2BG4W8lZBaecJ2PFo76u7OitN4T723G0jQlsr8beh8
8MyKJMnApu8yDjlBknSY7ChG6QGa/Zn2xUUFyFuydyvIfq08eeQGrHTt6I8MrtoogFHmQvgiJsvF
ZFbSCM4r5JSZgbUI4KR9BVRJc+rnw1wznA6RfQcMOUGhCphGggBsIA/eX9jdho68L2VbQP3iHSDA
rFucGTYDeqMNBbWCoOlryLNr1WBx4nD/tPQPL94yKFM5QeNUQVaejA+Szd6XCOKNAdKSEaZipQeX
bI5HbIMuvN9W5Q2mm+wQNiJ+28FbgJC/5F55Wqu7kukUFNJC49Z+1gGGWbilQkX9CcJS5JeCZ3pA
wFtFGZ3RSO1Gx+Q1XmE9Q8La0Bt6kxNvGpCnzve7UDY/ZZnimwOHtQfUwmdph2HthIkJMZnZfw+4
uyFrE0OtJov+9+DwKbfxm1Tb5O29zwdXNyqBOUY1rScsicG9sW/c3v26RaqQYgsWfNE9EYoEMkC0
VRmqVpPSFy9atBzjb16e/osjkdYAkBBAP8gzuo14qE2M9RcNF+qYyP+3wF15fXinW2tFg978sgKf
RMNBjRTyD5QtCN6bF0BAbjxGgtjW6QN8NiESN/tat/d+20H1gA3WfTKm0twcHg84puqaAVPDYY2B
QANNUIcKEvRmDyQn7edWg8tx+pfq5mJFcyUoyrSGQaQa4STQq2824nzCnJE7Kvk30fRuQ0lqv472
VDhZSRVSseBHZiNV7LJmAF91rkjCkU+kex6UQpEYHV3Qtg5psEOvE/e+sSYz/iLAXf7z2te1XgFu
V7UudPQzIQLlPgdT99JuEL4Q4TjwybFBfpue8LSZR1tuwmUjFpuMJe/eKQTREi/Q8XMj/4j6a1qL
qBskjWiDSfUVFeW6+FMOaxWQth45pSkVnV4MriA/g5BPdlnbMm/alc2CHnqTc40f5O+XNFMXukBv
mOQQWDbLKkd/CdfcasNIscrx5+dbbUqM0RjFPoiEgykhu0rQZd41vRt15VDAwRBpibrUtwia6EOp
NxiTiUaCgrQVaI3AaZbk31EjjCoZDiU84T+m5xzFuUGgLr/W70Lnl7m4YVx/WLw3gNj1S09zjGvN
l/ziyPgz8kgx9hxvPJ6IK8O1bvFopFW27e5CBBtXWYY5pneprGr8ogTamFozTrVs58m/sHL7sFrF
gBCx9TQW8aT1zPfSrPiF3Hp6NO1fFrqRmQ98hCtfme73UhtlUBaSA0v2x35GFeibmU0NpM5/m4E7
wVjkM8bol4pcbIzhY3gaKj6OQ1dO9wVETz0r2otp6AECOcavQNfK1SUozbc1sQKMDbgzQauy/E0m
dsScST8zn6LfvX78bAdYSTjnSgpAh9xASk7WiQD6DZ0JapKvHCbN1KFQl7JYd+Zs2RL8FcJBHuRN
PrWl/mtJjWn6jwCGav1g6hbpAPJtQQf7okuZsuBP+Hf/m/tJ2MsWgtPTPt2xLjoWCfZu/f14exN8
dv7EEkKYBrGEi5gL1klpcZN3ZNEP/MjyCn2fQ/aQxFF3+xnEs8CHY18wsNZWf3zRDrH0zq1ZJvNW
SUC6GxwVwMtoDm9gWQyS5JULfdEIxj6bMuRWNRuLJqgCkpNGaNZlKiQTBfex18qReJ2iOlopA13r
9JLb+Y2Q5QW+p7oy+FgA98Cp+qbBMUVtBThTm/Q7j0CzBjpA7s3T7Tedx346xpV0qwwGi4Ww4Bzj
gJBETvET6tqlFMDFBgHt9N4L+QcW5S+4KikQ6XjSxuZvDGI3IfdMU161SXCOgP4Zhrn7i7NWfx0i
EdWpDcPxt72d2tAoQkhhsHAzRNUG9iIc7St2vRDHJzb5zJ3e13RWZXwazzI1q65JD7brSnY0tTy2
di/XyYfSsP2eynMktc9UtLhGyS4NUpfVd+mca+NeQP5Ay1Zms1QQ/wvri0fKVWZ3OTHaSB9zUQZc
NvwA9cewJUKmaPQ+nFUCLyeuY5PUyE5l0hXpJKXPoP9rEEevc/MhjPz2R8GvBUNsFmbk4e8E2mkj
nKX7aGgBm8VT2pVVM0yRv+gLNK1LbYSnkMqi+EfVdvs0Czdq5wkpqqJES2JJxC03OcuM+e3Obsze
xZW4Kxro2Vgw9DCpSHNyjUKVSnb/0GQRP5C6usUPs3UgsdYRjTfUZxmSD2WlBDH5eq2MHmwLYWou
q6EqyXhTLm1J/94KDAGWA1DCH7RaZ+Yg5Pzjv/NwyutZN5cra7yMFFQAe5Oldhs13fivyPu1o6YW
TDvQSOx9f7MJYSBuhwfPDuqaDybvhrN/ClQGL9pkJ2V3PeaFktO4/9fxNYm5suzKO4FjdC5HMxob
9rqX5diLlCylpnRX/AqAeqfftRfnhRObvR2m3I2zBYj+1U5Q0cyopzZFE0FPjfORfieKeAscZ4ls
0DmfUTwzJwfnO07s+IYWqR/VRt5u3qE8wcoeDl9bXYY0nUpeQnaeF2x9tuXzIlmgWNmqr0x3X4L3
5sZxiv+pt6fRd4kRMwCfnzKqQy3ER520PzCMTWZT+bda/YmouD7VREUFia8jybHyroWkx2dBVUEj
x/gmob2uo9SjySrrcK++oNT0v+qOHD2vuSNtSVuqMOF0CO5pBwc8e7lq0VMMEiammkbjrk5pSJG8
ixIKQPgjlD6YVEphQpl0lTAxlDU83b7mF/um73Ob4emLJi4MigYrWZ899zAJKe85yAkpkXj9njMz
T7xgOyOdNxzGXLhkn+eoJ/Rb0AIUpSpJ4Q7BIZBEmC1mZz8vumab8/WdfzWiJuxoebLPrtf5UcPu
pipScamwnUzdSeJHuGVJ6OVkHE74cihz20OrP8HUUEU8pWhnmylXS6xQr+TVxI2Eig2AmBB6k7rz
9bwJikFHkJuTmgQcwNpUC/0xWmFhrh0WXT2qMxSPncIYJR+0yqlv+aXF+93N5a1YR2FSfamMpYhe
kz0n5Rm5sv2goUXSOn1Bu95dSBybb9pfCG50muuPQDx6mhyoopxxbkj/PtePyOCE1NFFjT5SVQwv
d1xrguuKOmrWO++2n923HTN5YGgoNEPiehXFF2aBCBbWFzIlTefFfwr11MANJf8eS4uyi/RC/RVG
8jxKfheO3M1rDx+Dpw+XTcB+s6ty8AModZWCl7H9KiZOu57lI/5lwkb4pnGs2YKJ4OwkmB+c/D+S
KaRaOpo8Ch7pZHU+a7XmVGJh48h75eip/OTcfneHtwtCnTyg8iRBAc/dy3Ebh8jcmFR2OIdXD5jU
RGAkxdWAOd02uSJNOd9pMLQHnqAEo4fGdoQmvZtPapAAuzwmO6+eF4Csygz0nWzeb6U/2n3adms/
lzWS2UrdnPIjx2W2r1WylnBeoBXxvzD/2j+oobUctH62YCcLB5Qo3eHnW3HmMjbJyUYjL9GZViUl
77kcFnFctOM/WdfFc5AsqxQ92ftf5aun/EvREoDMG+PIrj+cFahkSoTlhEvQIKo4inDuj6ndDbSF
1GUxeWsAvoaIuSz5ngNf7pXz8qDrMb9dEDbnIhZf6e1nOUR2nIxWPnb8kQjHdVUBkMYZ4NhCK8bD
vXlFj7Aj7Z8qPQ/JCy32Bz3R1wRCqErTb/4mG7ZqBHz8uu2LcIesg0B3sSKj8MwLgnOkc7SNrBA3
dzAo7ZbOKZe9YA3LB1TmOPxddkHpw0ix0PMjpjJU1P/gOXqRhHDtaJukeCTcZy9+KpUa0A94tjVz
4QQtLOSxzuGJxLh47ibzKTC1CVKy7i1T3ZZwZdjtJ/EKENkzUC1rhMwNbRidJ1cCfy2KQ7prJhal
JI17whih0yZh4ixif8Abt1Fc9ymUc6fwj2FMtvNA6sToPvgpdxDexTEI3FlXiHD/JEKGvupIHQWE
GLuuvPWJ3MOvph6YTrTKX80z41xjv1UBrsoOkEjkI0/PCeC4eRD6DuTeHqgg2hjrr5LCnh2P2nSQ
seiN8fuDLpwnXEuIhIPTORskehahe5Q+wUDGWX2glGORnKzQjsHs+TANHqBabiEdg/eMODLxjmPr
YSUOgjsc6i42LUHCFQXiu2BNDaSvWmEYzLV0Zi6sUUW8nPJKa/Lf9C4/Ql/gkjoeUL6oAOzd9uwA
Oecobt4F1JnPdaz5MiPB0wml8r0RoL353M9zcN76oqv2Rmk32rOvaLNFwo+2b43yzxvRJ+bZNIm+
2JrkAPlj8VMhCeCTECj+p6i30uanDZanl7oHBxUiK49ub0LOpALNViTyC6wKNLfI04hSj1M3A8Bx
uZb+Hw5uAZ15vdz6OsEWqNwV98HInvIEPeYz/mVAsXITKtAdJyb3C3fNJ4Og5RtInS3KLPVL+J3u
c9OqB1kGVvGVGV+WSAKaN/qr2Jf1ZuhkqLHdEh1VKkCfl9i8Q6rdWxLnSnl+lsEu0S/yr9xNE/pT
5zlOJy/k8GCeRuYnSiJlIZ5b5px/6WxfOuVrfikUNJK/g3Q0ZL+hd9fuu9WrtSIVOzd+BSOxFHBI
/Pgh4KRvJpI5p00WkGSWosoEUdiTKl/8siJUHlJ7NgzRdlQbJ18hsCccHwJOiCkiBgqAiLvkSlIh
LcNlO62oy+9d19CRtCI+72xxx4VDbQhtRbZuerLNjeOqIXvfWgg27S9kkLAN2oJZFeq8nexUV28l
REqs28Dvcbhbauj/Kh1z5rFAU6iVE4B9rmmNFyu/jYYO2oc/g04ZAUVTOcP2uuG0m2hIZAGzNss2
r64zpfuX0nXwKMc8P/6YPs7QUGwozEbf+3bTXSc/yQ/VD0Xx5GSNvpOrOkWaBg1Hqje6r9YiJ7Pn
sw23wzfXK3sRQ6Ay/KjHay6JYhnkgMhFwecKKNDO9R0+7I/4+opGvH7cfVcwNBTwNKP2SI40NNkq
XvHPD03L/t1zXRLwXLHUjBN60Ogp+OSimFPW+jjiAvJvGwdWoXVqiUjg7K2nTx/R1FFxTeEqdzLV
UTYqhbqDmL4dbdzInxF3gkD6FwfkdE1SCI89qislabgy2Hr9BmTHZZwuuSh0M/SnRLgskS4udUbD
1KejyllzNQShPUycQBnfZu0hcDwNkc+xYSsLg5WGZwo1MVvTu5dhSodmvQhYTkrepqcvkwD5BgO4
JM0AER4mCx7XtaDlm8mVLbGtPNgEcx4VdX0/fLq6gEofTV3+4u5E6aGTGMWL/TKiLB0ry0wuVFuX
7sXCiXWN9gmYjrNGs80RNn0zo/Ej7NbOW/wgDLgteYW8w2J/0dJ2m9MfzVOk1HvpdEcUzaxz0VnJ
Hf2r0/2Vbm/6Oxbowm3C2zy4PB/74/w3k764CQ1JksyFDB2r0RkHPTZyA+IpzejLXkj1uEicIRX8
BhKMx25jRAKlCpwtPJCIhxEbuOnSBKlp0pCkMmBxqR/el8VvgVpo6WmLWTOl69ay1ca6vFoDHY03
N+JQ4vOLXmT65uuTyxq9Ypsym6MPpKsUyZlyRANYtXECbg4+OsayFditcmtDNmmyoruq0ixTqHM1
vu2lpCHSIKtktP+TkpMxf6mMVi+/rt69TivTdIE74BZuZSw99JT+qmcK42YNqSnSyi74mqaLjTGu
824a1hwFVnG/eUT78KHdqnHHNrfYUMjRng1l9tGH+lYq8UNJLsutaAk8sjk991nPVGzVhrZ6E6Bk
MJpxXj7sQWOhYowkc8BstmVAlqEe1XYRSiwHxVSch1EUgXa8Tct2L96g54Fbb4TOCboLHdGTmm9r
ysAVVj2e0+UDzs6xTKZ9jdg1RUdBQoCP5oH4HVxGmzpzE61EGur5oG6yeZovZGusS7eiU5+Jdrbs
HTBUgPyUgbzW20NFfp6g+otSx0KAkvHxOZP2B99iN3uKMf+rWMkOF00BV9nvsX6FeAth5b12zPN8
WsnweO9gzgFTPMNnPVTG4sfo5ZyuHOgZjIx3cE2vnTvhesh7KZgjKr8a8DhJmVjRhlK9AKRLhPAa
Xsa1JS9sQJtsqpkpP7mh56F+5R3aRHwdwHSn6jLgoEdEQPQ4x0h/a2Z+1seC9QYFGfjsWtwqqvqr
kONRcg/vJtcR2FHGsfUHf1cug8fnYYxY0AE/eunTCrfneBVsOhf5yBagBL30lcvdrMk8UpV6V8gw
F1YZn4RKDMPqu19rIF9+ky03Z1Wn3MGBIW2YwAQaVSjXTFrRUUQ57lHeHfBfec/an6p0kQPjiIVv
Y2slIoYtYc2kwHtaESZxyrV5tKE+PTW/qmEl34qMqhK6tqDEXYwYu0YSMdtB+6GTlp7BcDfU1Lob
jfZRKJHnRrnBmswFP/eXqEXLlBxkQ7ZZFwaTQ9ngpdBaS7Rz5wNZNQpGI/N0qYGm3B18FEJIPevE
aS19QN5Rcj0IBnvY5BFyMkkGl2IZsLKm6XMAzn7lhqhyBbYqYWGT9xaRTLs411FeOpbdbyfZGG39
jOFgT6wCyqnvYfWDmS0d2vlxwXtCS8VW0eyf6fhwXln5U4d2/kc0bqvF6+GR0GkXEn28vJFuAAjS
YhvQwjXZZNp25vmCnPhVEXUQ4/aEmt+REPxrgUSlPpxrs91dw4q4vv2cQxZuly/01sZDZvYcE3Ln
LQxmOWZ+yoTMq9XcEG5pXIdnjJsz7Oi+TuR2V7ruJGEfIU7/tQ5yGMs0hN1inlvt30iAPv8/K3A+
p1mB7oTqzc8ifdsPmQ8n3t2vZcQ3WOjI4L7RpEqEObL5mFd++rFzQ3O6jXDQvLM64vFaxGGxnex0
dfIUHcYMDJndc3hgMVuKSZ7Dz84M6GS6vhoRHl0OE4mDnokqYDS2sog6p5x4P+mxfRgS8a3qneTH
rf6yeLYDfQeLOgwDooGIMirrLUTuGEtO4agCxxnHRXfmMuVEi24ONMFXqOMEg8Omq8+Tj8zRfpZ1
cVX9ESb6/2+fDJXhrRgf8DyJqgL+LQJoak3FSIEczdvKOaXhwMfuHklvsDmhI8+UtQ9DuhjVOTHh
tc6Y+qOvbiwSqMN2BXKrHUSEMYNKMo/RjyELUSfA6ARbWdYpR7+jEJpXOjpSjBeXIMDRIkLxgKul
T9YhTPDzw5VKp++C6+6+ZiKYYHhSJDC3fbS6FswvwKFcCO8Ky+z5h/dqBUNk4xpuHA4dTQZd08V2
uYl8JWZ0CBvFDqTYvurnKSLUq758hgg1/6R95vKto/k0QjlLiu5Y96uB/KRi4wJhN9PH12xwuT09
mq7SNajN4dNhuaa+s9mvhsf5+nkg1dJ3lifsaaK894NWRIWfDJkpT1hau3PamVA9ZjWgwzYf1a7p
AYUqjpcNhV6OdZtCjHfc3gHFYanrWFEg5hdjQKxwl44xRd1GjQuvc+x380f8248qta/lf9b6knL8
0ust6jsDqY0jyxzbq6vJHx4D7GDfGdxK6w//kbJEY5EY2d12z+HeoGgesZj5NjQput3FS4oGCddB
fr2TUy99wJDPzJeQZyREZ0VNN4sdQ3E9SajGb3RncXllcgYzJJ8DsRtfHi1bfgsIty42ML7dFV9w
6peDqzTJb72U+7yeBe7jv5lHQvHGYjHXuZbz4kwAk9duvgNoHNVA4SEukPHvcVVy7dE70RHXm4A1
9f0fNQFXC+aQ1GjCxXlX4fGSdTfTy2d9qK8ZMCoK1xjJ3d8C8vVAXwRzv0P04JQViDxJqf354+iD
vHmmV+GX2O00tHXam24Bwyvr1kuthDaHLB9tDC/mc3APCgMRVV+U64tkogqYCW9GtYiTikRK70Sd
XWRdtcqAFApG2gq8mmcD1VxpgP1/npOoIV3F7aIHRtFgwpoVO/qdJciLaDafbIHRJe/wZ/p14sbI
d34k6LzxwgAZ7R1SzFdffjSfPvyC9FoVfUtCx5kKCboA2DAShOzdZ4xynzZzpxs9XMgZrzTrWmw4
bIoe7av2nZ5/RWyn16TXr2GfWs9JIqlCVieJzjFdxNJAfirgM5aa/pkehaA/noFAxGCANsfbAzUP
fD1tKTtuzc7HMu+auu8VqDWDRkRVBDEMC5/6j133fuWuJUap9jxTJpILaPy2ezegsilMEcDTfUrY
FjjvzdXpDBaeA48tTM6f68GJjPxCCF+ZygSNWeHxrrhWBM0MleTj1jEkS/6O5vYtgXXXRAUywFOx
vJoRjgSM34jXZPejYpi6osmZNEAWLv0DHaKnsFnCq3eUv4AQFNoBp9rjiPKa2kiaDJC2g05t+hm3
59s1nfMndd/m0O95CF2w4qNRXp5s+sHn+LhkI/t5VGmyTgxUDWVjS6SM479X2Y7EkzAwEK/q5tqL
yMdJdF+dI+zq4Yy+sxSjGwBvvHdaptMhPyvLzNRA+/YxSY8KTRQy8OUwl2PSPRk+khBsQrVC7dgw
3Em8QwPXgGXyR0XRRQwSQ2vt1OhjUmvixoWCiVDIZo525TbT2vb5XU9e/XNc4xl2ZDL2uEMgS+EJ
tyS2Iqr7hqIQ8MCxqHUvKgQU6fBlePlPYocrk1WZ0CLwZyiA4P6Hbhuo/hGo2ZbBCuOzPTlTXWbL
b4ZP9wXWhINzz0jK/5ZJCp01NGCg6Qa0zSfCoOn6PKI3NuLPXBah/KJtzqmu5HNDhG4zjQVSgPG1
c53zFvZlZ0EEVuRzizcO9EXPU5vkJVd+TerOEzXvOjvyXEvN0gzAfr7vP2JcjWPOOH+VnyL60pzf
pdKURz8hMArXphFtWdMUTdK6KnDFMv5kPZ2lwe3yRPp66v+mQNlZEI49B8uzuATZUJyBnlTMdHlc
iYm6pfqPblJp8zQMKt577RpqY/c6OWmsuQOvYw3ZkrdAfk4+Fsx3mi7xeGuz4QhmaiJnHOoAVGCv
sTZNaedGrR6B8LpaQYI2cyHHKhdWMBOLgD7vOpzeaT5rU+6PpZXH8WFy2VLB2ZERqnn935Zp1OG6
dfcW/zU8zh9xBOmMANpK3ah5b6YJiWhw3kr5G54ffrBGRC28jR8XooxV1QbA/OmsaEZBH1/e6bo/
7JUXhGp1I3nlVDgGbgXF7EpbEyPErqUmDk2rdsJo1MbierZgGvSFy0Xh0z7XOEqbwp+RsDhkK2vI
FlvCGk0+ziOJc2vnNhKWNaAJGii/aO93QVoIwoSxTYEHZd9zzSAdUJMOyabKAi52UASPwS5Z+NVf
dp08nSl4WJwgxUamHa+XFeeJy1kPHnViaRHzSM3MQw/x4kxT/R9eq9VWzXeA8Jkze15wOlTOVJ/N
JnARfBJ1oUwL2ARGgfPF9lLGGapN4LqbNrgC9tBxmllJag5FgpVSef9VdRIb/DXLIzwTOpAoNgUd
bNkByY7UWJfXOv3n+zHQ+FWOEOZehjhvZ46ehgMH1dXmLIvKLphvAPfa+Ka8qsgwfIJNU1lUym/B
n1Njp/YgDdfQRLPDo0C8p3EAjcG4d83eWbJNUnaVNcEX7pLuWlVwL2lrRSazqyhWNSDXysvjLLoZ
45Vny7gtIMjB1/1uVQYVzP8e61OD31IXYNK+gm3pmm9Xk0A0f0Rkw9R/sMtPkn1TFMCGXUFcLOUt
FD0qfUz6hBv6bM4xL7DL61cyMgRqZr8B3v93+RoJylPwvNbz64u2RcMruXFY1LbI1+rhGBuRUsIc
nmCim/AJ1CrOeN5LK9KFDSTABeNlrPqIsyaVrQ8ZXt66Anzb851g1GJgFuZq9MAeaHgR6fGVdSqG
jyZs4FHtQlBYiPTq4yi5Y+2215W6WliL4oP2XHq07A2FM7acHj2ORgP+xHaFu7ya//e2qPXvUdR+
gdZPH4dDNqLxFbtyQtYg5Ef1Ixa6DIES4YbMEtPStfzZpR8T/SjHcQqpCHBGdJ+nWa0chqwrSURu
5e7NVj/DjurZespPbsyPfBrbofjLZbj+vDJ+8k+1MW0NSeJSm1t0OOda3qx1rvqhYFotsMamYoXP
YLyM2PqmA5ljdbXRPw55Lt2037X7Bs0N3NF4hA+IC5yhJsVwdDexo2Fl0D+JNhNrjeYCF9KkkONS
78hNC6PYUAZiBrporEEuguPGZ2bLlMCN7agkM0qfGQScBRqrfwJ7sxB3ZduGN9P1QCgO9ydLEOaq
H6o6QGDLFLZMIFys4mu+ZtIm0HgJqfCDrDhRqKEM+GEINQ3aZbFosOzmWmFvzRWdroD/8iTNguNO
gdZ0lZ1oDNOoeffgMKP20ocYQpRaQHQeIGytprFMeafoFktMVjlpXYQSEIVy+mbcCuwC4eW2nf3z
PbxVKX6PMbMWKy+6KwrZjg07TYqiYJO165ccp9fNE+1+R7HpvlwkQZhKhGnrhBw+Znegia09fFCi
JAN0FENhZ11pPr0Hfk4RNLDJ4aghGW3Ot/5fvWbn0MxK/oqDNaFq3268Ea9v6FIgR0cowfh1P59Y
/uv9cqh1oKcDIvqMPT4T75Mhp97SExfE29NZ2FLGiYztVudn5uj6y5kzK6UTXTuSOkd6kWeYTw6d
LyKnnP6u1r0O3xETax2SsythP9zUOj97KQKky98JOTgCDdpK1MPPgjnW1Do/ps8YgtwO1oUdxvyG
x5pnG5Cmemjp2dswAE2m8GdO683YyhiGDF0AeJbDvITCrrGMC3xMC+lNP02TRwSn1gwpD078SRTT
tEEv0ZcHf283IboNb1GQbnGATIiTyV6Lya0PyYYPSFRMwEQwxfws9KX99Cca8qKLPpTEzPJxk7vF
H+5ouqZskUhCel1EZt+o1S+FDw4qhZ3e8tca/t7J4X2pjTF3KwenxPuDRtEGGeuhaU3Cqpoqdtp0
JBVaZxjTeiiE2qvqwj+9yKldSuTnPSvQhglawcs068nAJ3qgIhw3+2h4PQWItwkOo7mCDiQ0J1/n
hevwnSD7QCwJHO0wsyDqX9+nzYf6lR14SCrP1tGdf3I421Au5squ4GMEP3iaj9PxGa8yqp1PGjKd
SifoWeCtHJICf6CSWdQgDi2UPAGzi9mQOH+ff9hbo8p25PrIWzWKQVzUqtSn+L1aXYxmJJNdWz9W
yl5Nobfa7V6Ofi8O7INc2cTAS9HgSmw9+ZXXE7Re9VOH67vvwPFVgYWoQ18GAovQdYn9do6YnAux
SOtichU7co6CqTkuRpNz+2dWrbhkX9eoDH16rvL/9KMyx+evjzt5wDStqLeVsbOXem9habDWnL1Q
u0zMmNaI+qIMEVeBvftJGKXUkKnN4Te4YL83mqOpio7E+0y6aQz955p6Ep7mgdQLROqkmXmLuF28
sU6TPeGPIp8LnVj6rnbZvE0zacqcm7c5mstdKpn2ZdVISj/jtYeeRc+/VgGthYJs29rxz5prZakl
Ysu3yQwR2iIpFxbHy0t4uOI828YIBxXaDPuWcE8bUrDEqwGoW6ioitCu6gTndc388fMOrc/Mv3Z6
lHQ5ukkddtKcEjg0Xbf7WRYCelRRahmtQ9tHW18CSlLw8eFnGlcscQKajuBm0B7Xd24wlb4pZEaz
i9qC600HsITq8wGXRJCbE05lWn5D2TkxF6pOFed8Eaiuy2QOA+XP1HMeu/Ng426QK/UdRZ0jiZM7
ofp0aGho0yp4kNGq0ofTMoFzjpsHB34OyVh5WPJZbVBmppEJUFGnU/TaEOfpW0xpmXD1I3XQwK9z
lw/ITYqHotJs05QNlpSNyF5wOSDiJjhvCSnbLwydDXal9iZ7ue+Ha1NWfeSXZBrH0qsxDASGy4ZH
qOoXGrmElywCb8ZTMUWD0OHXzUgn3TrRVpat81ouBLSCKpqHV5aLtLZ8Ve4P+uj7XWMyQgkcGwpe
HLw+FuFJPjDvgGzsli2B0xhsirOcH8T7GoBRSbN8S+xpbRmrGtvrUmOf6GJZML2MlqNO4gkBDHVS
X1jgOG4iSaxh4lj0iP+SZNUYQ1hZmcq4h15mxrWVCcVZgvERc0xzZPDIzWPF0nGkB/O02T4iNQOo
epHGgXUdGBaAN357o9urR8E8Lz9yiZ9PDJHyZRukV41rPPBYfMkVn2Q5Gjp5bCv5/UXKCWcJr51l
4eycp53LSw5vfpeNQGrL2TdmsBF4iYvnigPHRAcvs/yni9+asVuCO/a1C/+OCstlZRxRTE6+NUVR
AVfxSEXAfBLT4mBONCD64hICM71COjoZ1qrcs8kBHAu/KWUljLTkY0y4H1UzqCqvlDMmRdjwg10V
RHYkHvVH9QL39DO2cWrrdKdxcUCaep8/xCXVlqXbYp/KvLXs5dS3d6atICzIRjR0fLWL5vBMUfRj
u6wcJ1X0IBVk93EkjpAMZXmvZe3FdshTsy3KEpXNMTraTDUjEUbG6dydyynV3Is1ObQGjclvNbL5
tIqm06+GSiFL8Zv9wZE99nB+JrXzuM6ogy9Vy8WP9gmGNfLAxM60qHCAiJmIfAe5iJvEwi/eBPsd
pk6k8ccDathiWlSNHBz5IqMZ4G5a+rfac2Avh6KRdtjKKjqZCz26atk/LyNutYed9sPcxO4lnmxV
JlWSaEROJQkZjvEtaVfg7t+v2Kc1oy4c5sdi6B/k4dS3BFqtTVhzQmEFVU14jhdlMJt3ZwyVZgom
TjWgGbRT9p9xqbEm6CPbbGkYCuQLAkU3Rbj/hJ7aK8JmAhvwbaKZc7RzmyppbX66VcuZ6HB05pZ4
Z43UsgNRB2k8wtAlmyhtUKag0sDrF+czFThpkz+NrKD0Hk7kN6P5JL+k8SCRfBGrg8G+fvSC9mrX
dptMmLopSi82vxgdE/3gkXiKPiWSwOY72nhAnYcmyaNr7onqAGEoVuKhyF83DyWlHJUEO0TdoLDh
o4iOBTV/zfOC7RSNKF4MX6KCMCHkCaqnVkfWMA/Ui6GpEtROC0YdbFkLujZSyzVBavYpmqTyEcyg
ZEiKVd+8nJvzJ2NFt+uReJujK+aqsbCBPWYPM8H1qF+fplD9neCfsgmntfIwLYjE9BePUGglPiWX
ZhoPId+Sd8q9UT4uCfdI83BXAIqBdFhzCLqn//5WRCM2wEA7JE+9j/iRkkDnu6rzHPnmL7f+Gzzp
pdvrI/Q4bNOuTckX8M6cpmfo+WMQWskN6eEZLeFLgShdcxnbr7StTF19so3b+q+c5xGdjviy4fcy
th7iT3Z9SsOWbUYSFcxsQs9cfFRzVAqCc59zqxurtd7qKQDDni3yihmOcAbmpSYDEr+JF69WBhps
9ML2zrio6FBBkaGUQMzQkCPrTBXyNMHAV0qDqt5yxB3Jp8vPTdyKutTUOSSX+t4NBiWuy1Et66q7
4BxuQR9MK4XFXM9bqD9uyysyn5QcnFJr+sJOgCu1yIFdoE1PXgw1pTPalauRoWFKs13gsqWDhsbA
2m3WAhnJVl1ZK6gv3OgnRyuZ0xHCLsdrlO78agSAhW7/211meSgWb88nErxOGROzGNpFzBmLWQ42
BqOu11o2c0h8dfcK4F0gZ3A87Row5/MsKciFejWMtelGh+qJMt18kkEcXVV6cLd4wp+UihFh8I3C
qKD6/AUJl8j2YyWaQxTREBrsltG0qIr8lWWppesbvkss5xQIoBqWPuN7phf009cjAnSzF3Rn5dWF
0rM3w8oQm+wGnLVHDFWyvm08rSMcMIV5SUKADXMaWkOPmpcOMoF5cdD+l5fF9qnw8W9aib7ZshR4
vq77j+zdH0G/05OPPCoKPXw+sEuNypP1dPWExVl43t+bHej972k8d9AH+itLripxCZfn73BSe4C1
f2L4A9mXXuO4OEgJwquKt/kr1gO3ojAi7SElpR1ZM8BaOUwflnma2wvcehRBIcVHPFjlRa74OYgg
jDV+XGuBYjjJoZhhf4D8sAYYR3yeW8KEiQ+zL0MVxmaL+Wij6CrJqP/hCy93ozcbyPTwKVOTS+wN
AdmGbLE+y5GGbC2UZhbH6nH3fqiTs09fkgricaVshgf5tumlt50jc6YLUfxn9lREs8T1FQGREQXu
f2xBnEfusRBTA+3qV7nh8mumwc552hhcI/l+0DYU5a/uenqkULoRkv+LiTCbasY24yVyd/DjxNcG
A6TQ76YsuUssv70j18AJTA5d109Ja6mDYl79WFXj42E0ttcY8HnYdX2ZB/pht6S3/4afSrsb3kXx
MuQ/OQ1SP/CKYadu2J8Jqtx+DPAcBzV+recqc62ZPLmBvCbzZXmNUbMNKsrA/e+EtGqJVSCa4/N3
/jFTyxPEbj8AD3WRuaqELJC6U1ibIujR/EScRSlr+ZUe+cxdXdsu+DO6hmn0wFMh0cPb4S1TN9o5
bcFKMWjuH89TxfNAYZ0tbQxrfysDNcfpDozTzZ8qfQ5gAOKbE+0dZwwxDWx2/mZFEUu1dP4QllfX
sbBbjpFPm63fAazlaw9nRiLZXuUxlkK0pdbZm7//Mk1Vw6v0SrmA88cWXBTOE+CAHPQlMEfw5HUs
dpeefIdJdCN8Uz7L9FoOEGtQJc9wmQHDU0cpCMBPMqxOGGVvqaSIhXAmFXYMF8RP3T5dtJgP+4Ya
y1Sb0Ex9FJ4xm8Roi6aWLRXA5pPkJAnOPWPPRBpZ/cLY446bzEqAPaEJD8aA1eZ7oa55qgMKlLLV
pn2ARiXC2u4xJKt6sXZ0MFxhjtSkSRfx0+CXuAbnlMToNYR5vyxdtCBlTMorxTdKU6DbRNsxT0bM
nagmzyQ3f8pxInGOPmnGWvC10NwtTC4Crxeov3OAUYuMOMw0tPzEHuVgkeFzIZATnicVBaAplVbr
Dix5qP3/YWB4oEdRjgRR8muhzRAq6L5yRweWRG5Tk3pMTpJ3vxEuhqXzvqbMp09ti5Pj7Jv3ODl5
NaoXzci39hzZb1aGQVn7ZKajF2IrLi4nmNzdd+QIZZR7WOEe5XKCTa/W9k7U0zfxCUpzWXCYtP2z
SFMXTSjwZhugI6TtVROZ65ad1MR9gReKMDLvo5mQVxcWyYbN3ms7dNpUgizwT3iGblRglIHsX6Ce
ZN7fO7QPkJksTsYhKCMSGOsM+OQJY/ZE8cF9DuQEb/TGu78/C72Wjs0V6WQqWns5VxtTiAQbAwNO
BRDW91FmhU/f7DVzd51SYmpWHXIUOEKW5xtttDmmPZoudOUIFWispJEv7yM8sP8sWMbVzRI/do7V
DCCiwtBfLNCOQASfBk/sM5XTRc03/tz1Pl8h91ML0SGOPrdQRxaGKEPtCn1fitEQZQWiU/62NsYO
LN6TcjGXFCXNgJyoPrzfZulCJyJpU8YyxQZwiHlmG6autcTlFE3L/Z417Y+FpwIV4mnvjOFn7z1M
ekCtHJsN3vyF1EUDyCj1Yo/xiscBJUE7G1AYJ26EBH8oNHoikyWhMWiSVqM90bUV+8L++oTK3Drn
XAGBX/+vXuMKBYTEkZkUbFp0uH5RlwE4XDWVIcGbBAlrFpMKF/nZhTprZ1txF5AxYBXdWacaN8Zq
lGKe4pgpkc4hNEJZ/QTSHOPrZZXT5lVtbP3KnW14PnjX5Ma1O0eAF4+K/wjIwm80d4JcoGOb/xTM
CNsKldWpU6mPYlqfvOHHmQ0lwNBnHJXlO+O+Sgv3Tlf7u/uz/DVP4DGKmghWksO+Ed3O0MYX0RRB
gOGRKBbRO+m1Bta6R7YjaL7mvF8oRdfqysCDSs5ZqsbIrjiN59d98nJeIkEItztKxIeQQeUuLrWt
ICqnQZs0KFgo/4Lj0fM71/BlvYTJv8OeJrW65wCVEQmkfgMSg5s2lEPLJhu8eG/zw3xeeTnWKAs+
vWrTemhiSu/bJpKDP7JuvNr2s8+VtqkErWqCvodwz+M+AjaEgk2NF5erfLKr4AD61Z1PvNinAJsJ
AnUMwuZzJB+LslQbFbrosF2Dzlllfj1av7r9rO22BZbzHtkU4UYqRp6fmCyn7+7yNCQIYxHP+mPG
+iyhAzF7/TKRZqE5D25AtLDBEYQ4XV8DnwtvR40R8UlKBPvQrzhpIV9MwO6U0w7sW7bzCJdEa85E
Spau5DE8p5x1QXqeD7ui35woYoViBW487VjkPrXiA3SIw2S0+/JhojPkb4NNckw2B2tKVbzbdGai
i4ECyDidAVJ6jTjihcjTZ4mi0mgtIv7OmLw3PnsWueOIPoIqdhyFgJ0YxBzw6r/H/nIFHPsTgdno
a626j6n1J/q5d9ES6hRTblzcgfQVSiGv6ZTLS036Cpxrf0odVap8CPsGdD4BiwiqmL4nVIlqXP/P
x1P+jMUOyz6DFXLsmQ+6+iIPCN5EZAKT4DiONKGM+rVjGGQNheJO/sFS/rH0hP+omULK3cy53LPS
2krPqpQTRx448XzEY/adHSheAyn3zWt//IiYZ5x6+oAs8gALkDa53pRbzPVT1PTh+zDU6FgFRQ8N
E/mwLvRhMXtBlLP262GuwVhu4+3Uxoc8cdzRl4NmXH6m5CnSHciC8NUT27Y465emeEqzKOH7NC0A
K8xw6NUEvjxzC90Kp0QNvnzxIkcti0dOuAg/8B92P6u51KXw/BtMTvP0JPDbXAOmd09M2NBn+CKL
LdqjujlAcX4r4H8HfiOFKUKqK/S+tvStzpCONhpE3JDUqUQXO82vj/k+xpWzJ9EDphfWCu6Da+GX
F0H/w8A486Eb+qACuXipvwcHnF+fFZalDhZh7i1j/HA0immKbb/+SVzZeixnFdoZ/2Xu5IlRujlZ
aftExbcuLZMtgTpQJ/nEFoUkYqSInsjk7UzIdeU8QXHkE6BHqsveK2e224TeBSGUJKDZw5mnT8cI
QBhfdi0WOW4QXMap9wml3LIjCJlskFh15CTOa1HWGQGEEcp9Xd3HtUyhoksTsXz3Bq1yc8V7xL+4
JnFxx7qY0vW8OvM+dsOs4Ch3VPyYg5hHKWJyiAof+F/i+/5NDTXbEk5VR9lbZmmj6Wf+DjlaNLju
PVbm3uxGLpdo16TZXLJw8eewhQC3ZllMAl5GeruceMEHqZ8kKnfxQ7PLhBhubNG3Or+X/dBhDOG8
GKYtOc/rlt2LHa8s7Kb4WDV+kHULjzEiznTMG9FdwunLoRRBbqJ3F+GJczHdtL2g51ae4vxdTW3m
FsHtN+pUun4FANr3vvhRhXtkEqQkj+pLoUUAyIIDfTuW+Mh4jjqdmlqn9N/g9MugNEi1jNXq6/IA
l/Iwz8CcQHL5fceKG1o7Eb0L7aRjrZcCaBvL4OH6WIy9oJWqDJ3Nf8cqqX5HtE/LOVb/N21BGeHH
wd2roFFhkPuXVseyhx+X6Pee4EUEdK6BUVBPvJifx4zecgKeq2GmEAtUY99kjtcQMTpFUI1teD/p
6IGg3DYv3TQIrJs9Zu0lW3D2VpcOklyz3s1xPjSqmnH8H1pwBdAW47xEbLGRCMurwRsPo7xdzWeE
DFexMDDDVbTUKoR5cplPisBX9jRQat9M9ugDTm2O0xaA8qs6dIJK+qivkm0BYZ6bSw9iuhDPGY7f
iUs/Jl0Hsc+sOdzK3t9Wq6H7Zgi92BZG1QExVSZWWqpy+q07kHL+nkw6vxrPygfLer32XQ/yflt5
cQ1QvuKQ4dG1tE/BXGRkDnCBqAf+bZPsySu659Yk++HlBJF3q83jYIztH0Td2Dd1MAmCujzaE/J5
EthhQEqks+vAtiEBU1Mr34x7nq1fnlevXRYXPbth2Z7hWAkH9gPyGibZxZIIlNKBRipyhs5B1yrV
hglgnhbw0lwJp6Hge25oEW/afKqnubFrLSq7UEha2Zoo8omH67U7vtGF9wmCQuloJtU4Q6gRuVW0
6RbO5gs/L9+ZdKaN/USswJG9bBlJwSoUhvBasNxETRUcnlw2Ihl8CLWy3nP30dQl1EOsxDjG4Qa4
Pmsz7lSAYTDtVjbuIohvNihFdy0dxlRHRk5WrSdGWPLgTEV8Zpk9n+ql4dE96gn5kZRj7XlDQecK
6D/c+5jX8rNxE4WjsNCsNfy1ZikyBiukKzwZFWj/kuTh3Kd2duWuX0RXW9uzj18bGMqtgR4KjhRG
Ez3j+fYUzRqTqQqih2+QvyRL6Y/fUDsBV7bwvRaeCeQiwSeMJ8gm8cVyx4ffnANJ+WhPtJLI6iBJ
E6GUa7DKwq7jhn7zEG1WCDN58KG1P2ivktYWwwg7UODP83K+iAmAlTU27vuaxy9KCwQfXsu8jqX7
es+S67Rdzm7bU0s3NWlEfx+2qgB4bXuv71sVxdNNxnkHOZn18lHxxAnHQ5cvElCfXQiPCJ0nVgxV
kuTgW4qV3UKHnWdyFT7omSE/4XqYFUDCjpUTCsNU+5kI3AQcsM/LC7pLhE9YC7CUn+HrouhoLk4s
tRKvClVtD1yiJb5JynjEIPsMNMFX4TbSGzXysLmQ5dhmaUkM/chsaMIe/cHjsffedwMTcJqaDO2k
4VxVHHnpTk0hZM2tbZ2la3KCGHQZilVKZzxIYQgyiOE2djgCqoRCjk/mdH+xAB1gAmahoWnfMfBM
Gm0lqhoI7OR6K0GznP9z8q0VvbFz9pfwAV/et/H4lomI/4ymbPEJX69ld2ISt8/Y0iL/Xd5L7+42
l1TMeN3mblJtH6qTwmoLP4CQCOBdo+cS31IHVlVAMTnfHZS2q1zXlFLfKJI0ikORTCoq3mjfDmzZ
Ff2njzfZcgpo00mMpjHHaXB1s2T2v7/m73UT1ENL2cbTIoKvfpMNFh+TQaApaIglmAwylEyx3X6e
to3gyyugTNR3R+CjWEXVhSYzofFCP1aP9VFzshUjXMcCoZM1JfrAQcZ7TFn+MQ05gue+397W6w2S
r+fMlnv9g/z1R5CP7heUt2/maph4n4rfvOyN7dVQowTVWZnQ70Y5BrpfPQftMUVipVQFcsrtDjmS
uav49XoK/s7fY53GkANw6yHnp/Znu8I9zg/eDR4MAZtc+JWya0KvpCecEj8bw4uUCFYQBwig8fxz
O8kXC41Y4b6Gw/UVgscPxxnpBhqJgPGMviX1u6K978uaQghsCakz7I6MaHfyFQGGse1B11BPpCKe
r+VHU9wr3wPrxe1XLayKHeCQuB2b/+pu0lMjJe4leEwEUXzaSgCSuLNPhlUN1Jl8V9++wSlNiG+J
R6BXHAZPg8u5IWTKHQX6090T+hulhxFum0TU/3qOhqsosFyAWKpYmNN2MB3UYccNHH3d/h3nPakK
pyz8RLBNqMHvWMDo0BLLiRDWReQW3BpX55QyzfInSq+zOvL/hvIHe2j22vEwqkmGD2+V6cJepDD2
GCiSAWIzpw2+0AaSMIeQqiz1+tF5skyNzsFP38dG8NfzO4K36axJo2xIBntiL8YRijUnm9zBFik7
YmspUsWeYC192NSOaESfJrUh1AWpKxlN4gcQrZFrKLRx3peoC66n0hoX82EG10ahj0YzOWn9npyF
ybC60HKx7CBOf/pnpsvPZHkZc1OrhO0EN/Ky6Tejrm3i23YNWZIRfLDO8n/kalvcvga1Fy0eoDH8
QX4ea7cg+diyUcWK1rzN0U9ny45mCLC3hrxDC8H/qAzv8HD6AfDXyt+CHc0rbsfuUM6GFye4qpdi
qyU/ahjpYCvCKuDpL++XG4bupcIYnID+WzpLMT9cqciRDCekqjZSidQ4WtUsqhmsWKSLxMWW4PU0
oBUGjBlPy10GeolMRRAS3kqt7E8VOIwum/dNq149S6dqDJEMqOPhRanSXETP2Cg4q1gZqyQxniXG
0A/IKYspKllyLUzwv8nWgodJvjNuacbEYVJre0CATg6VTpWUts211UHwBovbH53lO+CGyvow0e/f
bRNttV+YvPdsFmbbhRKtAD43yVD8lGZd4pz4a8tjF6EBVCZER2uY6XpHRGWKWXImCM6FsyV/ujmH
iig9ua14RDvymEnPhIvqg3WAqz5E282ni3LYChnVWpXJ5zCgg7EDXR7d6vJN5Co6g2iX00hFi7Z0
CaKsSsuO95cpeeHyhRBL3273/1Bwjfs/Pz9KnjlJQOIW8Nc8vPqilmAlzieEYTbs9UAHjl8Plv9J
/gEv+t/jpBJFw90NSgFLC8EIfyqMEPoYHR5vy9HINNfagJUucjOQYstBUjy+L6jhPTzJ58opwqbS
PF92oUEXfHGtaEisXR108goZj3FlVsfAKp1ngZoPxzuQEloMjJj3SxxTDWZB7eT2sI9S45FIN5et
6i4R/WZlDmnz2+RkYdOUMNmHEK36oXQWJaUe8U/hyivy442h1taDTUJcnkBzRkEELDV85N0+4Ilq
NQHpGmnRjV1niJTflffH2pCixRB1K+wPdXqP9H77aA29JncfjLjbOSy9lSqE85rNc74yY85XqOKn
fhveYVDBXBbzGrKj9MsezCv2G6mlrMdr7qDDGVyT9P66+muCrXk6odhlD5fAaYieSC+2bZ858xPv
MA+6JZA9Z/4X39K8LUx1ZzSekOYcDn1szJCWr6Do0dd5nxUP6GAoLy3HyEG3QVJjbpwswmcpPC0W
EvY7MHfhF5bQuPeB+pbPqw32a4oXfmtKJ2aGDKg6/O4mBV7p006jZ59+lXGm5/WWh72plFBcYY0o
YCGTTDpcpozpEcgZJJBEb+VxWys5Uz4pC/NXYNXLO9kwEz1HLdzBnx/pUK67vBFKoJvOiZmEiilt
5YWyiR5U41Vf+T+qAeTJ3d2eklncHjaJLaefECxHPyh/pGSI1BuQmfWVHO7eUUAYDwxSouPZpH5z
0REvxAvdS0uZYUvLOliMp7qe0tmnpV1fTwdDXvJCN0oVi8c9LS2ufN3FR47MwSMMtYraDTGb93/6
c9H3Qe2oqUMEltSQrhDtP42P7Nne96A2/oc5ZEvseiuj5DGAyOcuHX7U8wh4tKTEZ77sn2HKjgpJ
jYGBkTvnADYYN0L14oK7zaLv+0cnxzXAMMTAO0DJ8gePA1XDNnF8ugiL50RyFVBtGtOCU8s9jb7N
bw3/KUwnSaRIdXv73IPz8YPhudQ9kka65oJmlhrVG8AHf9rFtXi+1qHBfAubN3S9n1/+LN6yqEYD
iaxJJq8CPiBYoDIb5rkqsj0qKyA0tkLShqLZsU39pQxrkV++OrlQnAsyAWy1GKj3M1pohHk7s3Q1
ZmtHrop9U0Ty+gxYIEm5gb8Y5XT/yJjS3LJaenFlkjrevZS2ecUeaLo2ELMrnMDZ3SpaTV1S2bZG
8PkC6Vs4aHgAMM7KtFaXJTiS29IFi6cAT6ve1yLqMOQKxJ7Vypw1kKDYBrpnSDUiPSgoBDuqTU+7
hCQuBS5+fR5YBjSUx5Ir4hS0G5tzIAR28gOVrBzQWluM7vCuHUq2Pa8mnNcInTx+ZqL687BGcmwB
uPezWdvh3ilupCW/0d8NN40te14hLlo+5t8uOs5sgtqb1w9Fv1oLH0LHq7AWiAkzsAFYRnCXhHyn
1r50LHmUsrvVAPbb6lTzz7CV5lSraZ/PD57LAQIL6UD7JcKv9B8zYsdaIdok5d3B3HWtOXHKq31Z
vYP35vyc+HvmdrQ8KAHJq1M8ihuoTEhmsYkntA8agLaEpq2b9AAxpE2Lz3GpIXONkOe/3B90fYA+
0WYoD7MBuIHJxVI9ka0aspr8AbAJLKrN6aShVojxImo7vsx0CE2K3K8ba0feqrBvUqTDw/+lAEZe
vmCi9ZzWWC1x/OkKAmqdS/+DupE+b2ycBGBNb5x49YVSuHITnzcO4yeWT6uQCMB4XyvoImqKQg5c
kCKL5VZzjfBqpg1KSLTtGB2uCbdhEA6DaWb/63Yl4fJIE11niIdCwtZLs5EOoKvOY23lDfJKFITW
K3kABxmJInc9QrtJ8JSXZDD0jLgc2WwdBi/LAJgi89qtCz11yg4spDoXQN2gq+2GqluKPVl9kmM+
TSfu/E14ShVqAoRAPfyFBTHxN4rbP/+ak5iVikM5U4Ro9SldjT/7nUhaRNO4tpYNeed2XKMmcOca
oBcz75FRXL+TCWjHKZ277fsv57Wwd4HR0YDdGQaSmR1HGqttqgiXKil2KZnAGDCtSU/7Tcnf36se
u0h0AhKAHP1sIfadPo/ep6vi0iUCALg9W48ZARWUEetH5ZZhdI7A03w26YHn4oqjQgrwqZYeB//Q
Iy1mVQYSpJD2b8R+FYTkcKdgCV9K/A6BbhVQSYY7dMMatErykPJMlgAokb8LsNAIuXU6w1xWODNP
zpcDaDWyKmf+6XmwHaZJ8OGGu4+QZNn4unb9jpzp32I0tC5W6mwgLTitAHdnM5UexW4oZhj/vT7Y
BhJQLCDnqbLmZcR80p0cXr8uub9/8n5z/aarwPmJvAzXnUqPF9UCic9qwRsLIo2J2dUdyOmOOKfP
n1RruNlNRbqij1SHuqZ/YAFZyExCGXF9jdvra+I0DvOZX7Vsaf9DFQbOUOX/0gLe8GFQJ5O9938P
yxUZOPVoJVm8n62Zxkt1mp72RV4O80vVL7BH+W5jW7UFeqwstkxQ57qhXRnHOYfjc/b9sZdoZcvK
7d4lPlUA+qp6L+WfuhJ1viZPK1/heyqDRTe8lzti+B7kBI5LTYSg40EhF0sVzpsDnW4lOyRIU3BP
pVD5LSDUoU4sgejHcYdOCPwwZy4olYm1d6GHI0AvJAYFUiN6oAEVsgaX50zB3IMIV9TDGo5s6cU6
qvMs1ohkOZwgidExky1oQRNT2ldLNGVPJDE3NQ0uXoKHEdcORilREKT1sxEFD/XQvsvNraCGfVX9
o0a+d2ks4QePZvTn6099PTVQzAKv5xmgCE0F0eJnrdL6fKNyRoQ43o/sIrw8sho0suoKIYv1sCet
IgnPc8QdAm40UNRIsIvlTw3zQYfgmfUmOwXLvb2Pht7rianpIH03Do/TFMJy1UBzBkjABEvMMxmP
UvhWVkpy+3pCka2rTRoUynVR2KtWc970oLMf1uOMucTiWf7vWGi0JjiuwWhfW2Hn3V6AHFQl2eh8
Ngx0CXj5tkLoX2VX+E0ao7/q2//Xg/jnyw56ic13VXcS9Uz/ZzlFPpxGTjJ74BLNhYrLggFPOSZI
G3taniRXSyZF0xZr2PKJ7zzMk6y31hW8xWA/snNcPhf0c2vj0zlGdmis1bvoxYWRoz0Ro1HZqysX
EYPiNHrKXZGjB1QgcwVWMukQ8Dtc26HWHlLCgjVLWA/d1dOoDUJAZ6SIkmHNn1lJQIFOtWxm18Bx
UXZCtPjoN3e2JLNP5I0SZRLFXGPXhM8dtkVAmBJPljxi2XiYb/6/9odncuz0USGcUGtWH5ifRBkV
3X4o6xdKbJXWxJPh/5bRF+crGB+PFfeSpgOLMSOTkEuQPq1Ylu7ojIwtHjILc3kClw0CmSFChpN5
r2AzARvE7pGgAktlR2yPxRnrdy7nJKRXEAR5F4uOOEBcJngPyIprpUJAQO5hRMN9NF/3rdpIu4Vn
kq+DKreMC8yx/8DfG3zV1fBZcOhdA+YO2tcVZ3Gz8G7VmX8tjYnTdmiVCDTivHnUshM52CTXiuF3
GPOBO5IuT+Pee5PlYHzav+i1/0+OhqOKOAIjwvXN2Fxqtf77M/0le3IPk0AXoBnfT0jCNcl66j8k
+tS4P6rMJ5aGVHg5JpoaZE2Yp34cTrwE6v82rt3WD/+qb+Zajq4mF2yldyxAgoxdXcuF0MRZGtwG
YHma492dOfWhT97664AUL3LlKLTRx/6fpfjPnvo3dDdIsv3lAFlcHTeQAyRx+PMdwFbOQWMoFpEH
rttOrVd2G2o9o8fPNs+D+1nPq8ItK7stMLJdPWpqJceHNM4ojmOmTxFovymzTFCtj5fp+SXulCrd
Oz9yf7UtF347U6bLjdzvzlYK796eEJjEam1QjobXx+h4qPHjhzaJysbx3aZ3WzJqi42Xd6i/fmON
TwYJqKjNXo7U0GtvtI/ucdRI+/2Qg5u8lDB5CzIxbbkW+uyIrp9CSE4RDQRRKxXQN4lKGWKhf4eV
SailfBw2CVGYWPXDlG545ykJIHYYr9eAPEwJBYvMGnpn5TDy4xnr+poTTTw1sUm3kMvulqW7r4Aw
/a45iztdcF756+xByueW7u4xKrsqoxl6fR53vJk/WmCN9tIMCOxcq8ArPl1xGqsF9SurpnoQXDe0
KC87kxRy49MCVz+KQ2ihyp3TBj0sOvksqflh/2SsgPmPwWOOEZw2nnm5CIMyMahvTy9q9H2oSqpA
NDDehK8YGu+ag3Y/d9wX/y8bEadKdvBVDDYlqpNoLxdPdHUqB0o/VKaduB0Onltgx8HiW+hRd5qk
AXgSKTsdASSE5M9mg3433fOoTa66A8c6BaSsHZ6pHa76CbFeD86D0nVjJSiVMcs6ALI89vcoN+mQ
tcVQ6E2qD4cR3WQLlu3FcxKGAt9ZAA8NZcHxlH3k1zO/3LmoOzdFq91ixyMyLwDQ5YclKC7uF9Qq
jIkOyp/Aq319mYzPq/5QTHK/9WmHjoMMHTE29JB28D9hJ6qeAHDEjkP9cRK2ppw4wkPHsHVECy/y
ffB4oc65OoqKSRPwnLXmImNqCROyquizX6BvIdd/H2ByFOSNNGW/r7/U2Kf7VnLbAeL6rDBzQiyy
X7fwD2PtiuEb7MjbzuP4CbhMzSozttjC7qQnVtgrPBiVi5nRzWoehckDfsNv2f3JOl2qzoiHS9Po
H0KqZtMa/DXnZ1rHsNjqoppsS+vP8kh3NjU4f4Dd0oJtPQqXizguEBGKzBy89+Tl/4AQKsND/3uJ
KNaK3lLNmFZH1pVYuGpvnhtWGzktXTa7V9pdxaaUFx4abY1J4jMt/T9aD2kpzndQgAwU0OQ4DOf9
sBULTiRGpOuKFfpkB2SNQRjQXBoeB8RYfbnem7s2eSYX2oZpzGTQSHtWJihXJGy8rfKnEre5tjuG
f6bokjxLj6eWggGiYxNSabDgdxSBZOrOpJKe9pyS/u45Xs8cRp3fq0XCV5UsYpuxeZaRbxt988FI
27V74nS0uxjsUwQtgcjaUySjwOpAcLWaIWZMawiKswz+182aWT3jFu0hOpTLD54PLe6A1YCK5EBG
8ELpPpzePNXSxJlxp0G+qKD+YfBR7gQ5n3rWPB4MjcRYqD/b1O/DzjVfw221y5JLwjgk9QaUkgz0
bi4yuMZYId+YeXq4oTBmhXSHpJkVwl4J+oV4RohLlJI2LumnWKefhsqpFyRJA2q2vRM84+EL4MbQ
narZa7WTtpDCBOJe22p7Dcfaq7RyaQkdUmBlju5w+1TdWFaz6gPuAw4TQ3cbUxkLLctUo1wyb7c2
CewNr0zPyRRUpK6RlYFti6h1WebCwQcR+ciWfqOaHa8Hrz9IqeiKSLOUMXGKy6Tl3a3Xb6+DQ9+0
MkaMbjWiZFjAVro3eHc+vfdR2fAgTV8Zbh8WXouguJYT39mj4lhxk4puPftXLWIAJ7SN2XgGkwZo
oluPtFTL8KlkhqWpn3nUHtNuvDTKbWPcBfVqxFIwsbdGM+qHoU3HH6SeCgF2t/Rb6rDkG6OkU9I5
+t9asw/gHrX4GQ663bqPgWqvj3NZmRrBjyI+5pm/bJ7H57Kf1lDvEGCytmkYJxr/8jjBTJ/qJvop
MRjdMAa4u6dkWEnU9ROi9HWMJIz5dKe6XNzTz3ZGAKtu48A/8vQiKlxA2en8TxN2Y5w7JPrEthzo
LZdlRqm42uj6+ylzrDC0OvAVPt8/OT/vdJ03Br0PVGRdB02xWI2Bw8WJLUEaY0eBIlbi4PmmyBrL
YDSKlirssFzqOjgposl+KpVyimprEuIbmOm35IXwDDRZz0Bl/5OEOD7ldXtPxoeHRdgKuZv4WuKT
SWJzapWWfsOiI47lrhVOlHvvuxiyMJROHYcnXIgwRxjk9cNeU4Ihpf3hg0QpTDllDLDtbBiLgN/a
irSps5HMw098OsCPa4PJSrvyN0gw5u1dNcGzvFZV4pAe2JTOVzVatr6cXQTP4lQJ5nBzsTmjElTJ
Meps/5xwvTbYTfnhtZWoKu9ZtFb7TGVN5nSKFeVfy095jnKMsosReHcRV/TpPvwmNk9DiSsbROhv
SqLNCI+rB5BtwY5XMmYS9ehif+RGzeVyJlatmhgVaDD4KxY67ncHXefBe2GlsDmfuOpcFIaYWWMo
loX7zHKhDOhcmIqenqXTjXAqbS5Sv8LNaJUHs1bgBFkSPsex1FRInoSQuC88/gQlmxDd/N00eVKZ
C1CuLopogTpBOFRfVnSdLt3Xel1YKoM6bOpO5Zba2R5YCaD3DegLM7V4Rv+I64+qr3C+hSvIJN0V
4qyB+LTV7E+TLmYhzN4aKqa1cZ4mYumxHahHI6pMAD+tZAKv9VnIe0MBq5bpB9zb0BHM1JDeWgD7
0poL9gk51+griHaMKtVXcfakQjByoxVCvmU0byx/R7NIuGKDp0XNB1m6CN5qB8TvqdlnAJ06P9sR
Rg6vfw+Fhjt6mCCcmJp7VV2IE5+CZwXBLxYeZmNW5BZXJX7IHpY+LE3eYyxaVFL1CbSQKpbVP43j
J+CJt2vsYqBUky7RA7lQHH5jxolUKc7ihay8TTKwa0RC4/MRofAsjuk1wG54/X/aXS1caPX/3Bjz
nmTkLkje+JJu/F0JzDvX0viLdFpTuukdIF27JHyq8BiTaetX48Ec/dClQM1Kzyo4edcLg2tWrKlg
Q4m99KL+rFPbtjtDbS5h17GY7srSQwNJbUNJ+xrOHWAJUyBTdHDxSUS5wKa0OLNFG7d2cf4hgTTI
rG6Dmg8kLDf1/nYErbHVIdMOr77UZ2DO08B6+OzS+4V6eQbTUpQRRV9zg+DdxB10MDvPW5rzs4hx
lQW36mdoHvLqWEgi41UWpQRQ7t+umP7o10NUUw7iNpIl3PFvxEZBl2hvpD2ocQ0zSCiT01Qw/vNv
AOJDQX5vg3LqtfLozUgkawxEbUHgaY0remn5GBM0IDXwg7kKP4Q0TWSIn6M6y7sK5M/WggaOqy94
BT5UCoauwMIx+rSodUdd8JVYt4jRcxrYuEuffPaCSMdXRGwoMOOBQxEeqhplj4wAgvfphg7KdDuy
ZUibrDyb+zutNCl0QFc5W2aVJTRNXyl+tfGDdG5nOha9XvK7+z7lTrRpQ6r2x+xX9w5ZLPJCkQjw
mFUnLfPwoPloAEsreJhBU7RykYfCMqpGtnwN58g0aqEEitYqzLIYVaR8035Q07Y+1G9R9D0XqgY7
bRLgs8kekcRZw36JB1O2tJho0VZDRMVElwzFxyLFicPB5RfHO2RmlS8rO1gXVOQDqA0bZwwpYFYY
L+DwwEOVuIE2S6QWxFyWu2vILxMGGLsjUAp0uQn1Cjo3xZLKt+4uIJQ6iZuNsktxUeQe5pyBxN0n
kW8OF3nMxiT5x39uZNFLNIeGQPzxoLDLdgj78CNf3QSD+yGVlGP7rXj4cdJ89Osc36NAxNzu/wBq
eoM9yMBafTC/D2ynDzxJrumcwoiviKDrRTZp9pbWneqp8hppGXzsU9CTl8U/GrO5/Rl1D63uzXpY
CKDkKlNfb753rc0AyF0A2cxEf1UB4KbXPpeC/n9+pcIpXNFiQ4a/6b1Xn9+OrLTNhXP4nNyPJUjJ
u4bs6qx8tDgWiZTcNeS+BDBUdxjYlFtD2z/CtX3xj0js4U/9BDdoS9T3yTO+Jo5UkPn+cMe2v0ME
cAh200Wp/7+5wdfW6ZOiGbtL5/T6H88ZG67Uj1Ong7/xSy+eRF8fcsLslxINVmVayn2FnvZdaXu8
nZgIgTQgpReQNlzqpUrHnmplEAizGpqrHty7p9oO4jB/G+bZgF8QGEDTo1xgq0VnT8lt7fgm/N0h
itXFyc0UydsjI3FuSw+70Odt7fe8O1TZYcnRGH9lUrGSqdaUYMvHSWbPeTZ3sByWSxvmkt7Is2DF
lH5xwin+0CEETwzlLbyuc7vA+cerRrVOXwEFdzBGWe8yP795XZoeVL6ql3SGvx7b6Qj2tWZX0PvI
v3gAuJj5QHKMo27TineDMz7dR4wlD9vDgP8hIlWeCVuK6pXiZ7ZYr5/lcXwFDbdk9emITx/WQ8cA
Lyn34CarslmwCu8etvzWR2X8J3pAbnrwAWUM0x4PEwNOZzBDo/OqjdgbmT3bOmLxEs4DsD4m/TQd
JM6pIeHalIcEAt5IFm4JtwXlHq6zDq0nVrwIbQstzmY2l/sOpAoUGxEDA5c1hetVSFbVHOsbrXC7
z1H862qKX6E7tmU5WC+tR/tujz/qqisNCFoY36XRwZS86IzGasT3pi5Kvkez1Tzs9pfPt/fBCzla
SHXbRQixmDvtt1NsKtMsSe7vHoWnBIQivKJkXVY/PrmBxu/BRSyU1OA6ypN2cSE1HUf3B97njGbQ
myn7tKEEZsbAoQ6fpjbaVK8PAH5qpmrq5R5x2ePxr27bU5Qf8lYsmCEeLtlxoqdeat9DMCyYTWL8
L3j7GLxfi+391WebCZsJ/CpLMwPqwMmruC2BIqNf38FQUqMz9OnYs8midZxEAQQCys86syHSlWMT
KUK/MS3TTM5I1tB4+JCAMyjDkctO/sGtvYHfVUt32RgWOv6vl57bk9yLHutHxJm+3jF/zEI90YNJ
oyVk4BBVBa5RaxaQJerwEC0Bv3gR89HxUuJ56rkOxyC6rMx9wR/2pO3ijZEMfwit1y+ZpHt6zQE/
p1c2K7GcQEgrRlYk7kRG6EqfWfM67gOQvSyiJnLEDXl8HzgFw4WccnpBaIU0FcSDqYlKXweZ9hmY
do0FBolpmCTIOpomZ8OxZDYR9joIQN2Re4VPFnfMoMQs2P52j5vk7TTg8+d1vwoTvFpf/tFlmVbE
lKOMWapoEDBLM8g7WqYfMrGuJo3jlroZVZPMa2bzxS6fiqu8v3Bgvpi/5HBH/W26FcUFrqOTUTga
GFtSGikvYoZrDaSuSX7ozq3E3+ct7oiFM0BB1lYwpH/mAnwmFrJFs71vfsjMlkGaMFXgGao5OCsr
PFtAZB0l0Z79ifoa9sw3t/Zo9to2ZZA19XPGN8OeiRAWdCIKqHkepsF1A1mXd3vV4Nx8XIgWI3be
+e6/YjYVgKD0ol00c6iCSi3KS+ixFO3oY14FlvusLDILBuvHsZZsV9GONBjIcpqWNDZcUTLRGaue
q7lxCvUMlfvRyq+3vqxoYFv9AIWDWPNUVcWmIg5jQtrfFzRIiBMLhGPgRlXujslwTm8l099mGiHn
WjKNQlfRqkg1bEj9wAw8pNjLVozToMdlRHb+5UHybZJaJGFbn18deCyg3U14qLe1OdDlYQhtSQiz
Z3c8yzh+FqkC685zCMRTHf8jnfgD7NQo8l+mUJdSVOVkDWpVwwd67p/q1/42NLHkyzbcWgY6VTiZ
Z/TJfybaXyv/EWuT7WO+sG68HRka+9Cxlfn5rapX2Hg0Q5lIgWsXE47U4KA1lPPGAjST3R2GS9Oh
2huT3+z9EkvNiIVornMxLg7Eh9gCMc2NL4Lqs3mIBTPO+rmVmAkT3dKm+liT2slfaplRZHf8r72i
bDIJm/VAWZVKZgLQ3P8sYFB0Rn43u8HuzhIZerltMxQBmgj1Q4B8a5yw9XEX7GmiRLJPSYAVWKZU
Vd1k58vXpLIVOWe2Pl+OMs/3hAG/2Q23eo7DPiYzvfsixV6Yg7tAjBuzRsIhEgfVoDo7Z6rrtKpG
etPHCAswoyDQhTWOywD+Opu6o2x2movNeykgzwQz4iOvihxzTu8L8CJcL7YDcbt9XROj8gtl0/1P
OiJBZwQ9SZo4RJco7mvwgr2RcK3JlcnqbVXuJZdVZu/2q2VknjYM4BANPMjWZLVWC3boUcPAZsyy
ni3StnFrcHKNyyh5NWjkhLHyxF8jqP6EEHGZqqVsXzk1VJ69eRj0BY1xPPF8zDNZ1xvdTyXnANJd
7gbD8ZnZ76V+srrywtawEb0SUGVeuca9L6y6IY/tpFsQu02bdvMxNqNP4pdw562EzGRRwgdV7HaU
CDcw7DqkoBvBPqwBvMOPxYiRpmBR8ZMb/Wi2TpPL0QbwywcvIXt8pDzkWd42Eipp5tc3V09j/YrO
vMzsOkj9ZznO2aV4/ks2y+AqMD9gcRW6DRqdKiNZf1QtdMNKlLoChqgB4VeBzDGJke2RrQtPT3nQ
sPiaR7Ioq23EyYfKlujDEkbUl3MbYFwuFuHoEfoLoGiqSTwu5YlcZUW+R4sJVSKwYOCEyS4+bFe/
uMceOQiwI5xz/RixfYdYhWx3rqpIAXD6ir/l/CvikVs+nmm1LOWOp+FGjXcbcKhxyboFNZnptghp
Qyqjt2FkuZUR1LeEbiADUyY5uWQFkdV0KShK3C+9kJkINflZKrkOgqtubSVrII6dWChUdJOnjRtY
j42ikXPg4Pb2DjBQQZddj62D8ijNnuin38PdWTAvO/GINX/IMexF3sYsKFhsY8gyNxbpyFt6iOh8
aAewMZsoW7CQde226onhAuXGnfSu9D3p6AfEgwTmqeLlyjBkN2PhXKLqi3BUEgUBAW5sl3KDseWz
tBp3Eb2w+CiIYgQUDT7ojSs4kM0bh5Plkup9zURPjhVwlTSs9+Cl5QszE2z5sWv+lmFZP5PTZxqh
oM7L79FmSYz2zpoxaGpncKdEfUUk8uscNdqHrrQCdYvWjThrxcZ/0bygohv7+RH/QeeD1n552Y4T
tvVDvjGlJDA3IcYBt7KcsAl1xxBEvepf6wNhxaQGPbVD/gsIPlM0TezrlX3ChCvOtFRXvZwbOZRq
V/+84ewRzoUwmXrJnXepYhQ37tUefKQefJySi7TZb9w7Av4ftpv64gRoC6IO+fkoh0eHIOkT2GEh
O8jZpvr1IIuuPHzsSTkrQ0+FSI8tas8LuG64vhM3oGETcWlKOb1fS6YMBjcuq3+0Zo8XF4dPN4fk
45PB9TF1q/+3yTXIMu7uhlBO7E7eUTW1lGGIR+gU0X7irztC4GPJJ9GNpztB04++UZV6CLOgRfGr
U4Mnu9T56i1lTs0dOKUIy3Pe1hSjyxQQC6XtD07hc/Bu5NkAUrmvODbcD0vw4TD/AE8ObG7/ix3W
TcplNvAQE/Y4fG1UkWHvwJcAWwZ3wptbgnbNYRg6Wj2ssX3HnF88xir6klSjeMe815AyBH/zHnip
1866sUlD6iwSY3FcLRlLGnj3lrGQIXKYCmPF9awfKqLMujSUvgOSA/Q1YyYJ0S9KBsHxwt7mYcmD
hKt1746e3j4aMHmN2j3wZh9TE0D/CGVr6NqzUeqtNrM93EOLYL+PvguEUYiMdoWH8pw2YWrAMk6n
wQkLdHUDXEF0S65FRt+aeQtfihNo8qt3RNM2MQzsxSwUxI0KsBKG35RQmlFvAUB3VR6q/vn5AVLO
zKuLefmZNyI5SLpHcJjNbXYEj9hv3PvguxWD2/k7wTLW7y85QyasvA3FD+SIFHdMCtjfXHtTZdTn
l58SvIZ257g/FobRpFx5YKDXJli3q2NXwJBEsc08e8YHubRzeWFO/7l2wfEBhNtby9ykkyllYjmw
9vG/jlpjeHxu4XLfR3OAFoR+t2N2uofze2+stmzqsUofAM127AAwr/7tFwQSiH6U3V6jpUv+jrFF
4O9ednMY/uR0pO138SDg8PA25vbGBnq+y4tdUwJ6U6n1/RCSMjyi3Nd/0XXf5uFRnpd5o/JDupJ5
2OM+IXLQWghTWRihOsxZS7u5VBDARbo6h8fFl0p1QOpj4TzyWY7gNvxjp/c1LwhhJ5dItRHwdJF3
wrHTmyNdHR5PzCPMjBwrBfXrYyl1C+DKgBLpGJLjblERfEY3PU/pAUvQPSIfwYCyYFlTPzzPTuey
GbD6VgAldu4PnC9nbz+UffNY37+ATrt5B1IBhN3RkZgV/nkjKlecF16idgpL3PMdPahNlLqcpME/
PtwElmdS/jiCsFFl8QdJKkEJ4c8wzzq6u0jFASJcZ9djMKYH9eb6BUpV+Ve9fUqE00RowXbWKnwJ
PWr6fR2HP1X1DQlFBolVyRY0hqEwj5dcVDn9QknjjdAnh8yZWcwGWccNkiYt5XIeoM6iRxEr9ALL
7zBgM3h4Z1CrszxDT46I5YP+mk98ADebZMcjmXcpy4d1Y1anCElBRv/UA8ZJHLG7ymo0zLAnowSt
9z3clLXQtajlhex593ZWLpj20Q51lm5mpwprwyTpUVI6m6+RcgGK0QbzvGoCs8sqOm97/f5NhVVd
6/Cpucg/ftGoNa2U77Paq+t72lgFY6uCJ48WbrEEF0fAR7v03xLJhl2ykjlDPDKCKM5mBkwBvMPl
qXg2YofmDxEkRG3+d52sQsD311a+eQpXJIAB1ZtOcNTvUnaH0e2Arturnpd0mI0srEqkElIZVq9C
qxHHfp58wAx5IomyRrTmXuxt5YJmQTFT93qGFpnfXftv2Gkoft2rQ2bXVAhe8ax9MNQLPXbj6MF6
wFQZVJhJMgSp8ob9byDFecfm0t7wIj92T/qhfylMh4Xh/ioOZ4LsUI0sJEaWtso4fLrTb8B9yJkU
M2TBj3xVk7gyuPWmJ1gYHIJDZjct4Fqn21t8Kik5cMZTpDGG5aWcHWczC1E6eAWeo3I9nPKkk095
HlWy+olx/UjVithSs/Rx4t6M7J82Rkh64ZhbgiaHhTellrrtEvJOSoWj6gYp1u3365ntK1dwhrrZ
ctwtWU+Dpcb1viOQmAYZLESFvKZL9yGfp2zUyOh8Vi9qRLBSNvmFLGOvfEsADw8QwX53Ks+lzJmE
NprUcndIMOTE/HEgeK3h8ZXuGUbTn4BojhR0FFI6aGb0IA9q/WRJ6i9uorN9y5MGh9zEuDqjb6MM
WFf4OOycoTB44wd2S7SVz3jvs3miqKxGdhyvrn9REuU/IGPhSSyv5i30vn1lLTB0CP4l4ZV87Ia+
vtJw6touduHlnh/kdp8iJK4YCu9Jbn4UNlzWj1pj/+7OBwnj9hSeDX7YRMbUOu7aF8+7Q5LVeEoX
LvVcFdTlw9ny14+yJMPMm7WhzNI5tjzTAgo6SpPtmJ+XoS59IFIInMUCsmTPZJl/AKkPravy51hy
9FQT8ghOAoM+757PErJOWhzVLsNydembbLzmB0pm7WN56MphC8TSrag45oc6ooeed2dVW9LgeS2a
cdEekiU8t6ASM1Cz7qsEAi3A8+YqnzuYh4fwChCxvKN74J1I9xAp9ditusXZKrCM2OjKVxW05WqC
SI60K1eBu8nCWF3jqWsG+CZxz8Ly/SM6f4fYUjPw4lvDMwF2WFMrQnRFT1ICmhUo5Yl3yIqfOpld
L8J5zufXY2iuy2DQPNcMvwP7fzfwZqlV1Ewdop4YrHbnH+1q0rqwR91guXhzLPhTB7xIz9O4eqbN
GJHQwECP2RCcHxUVQ0iMuNGgpNI7HWtgIzczmuokISF7WCwSGokQ51ADr70+6ER7+vOAsCaFMDhQ
dutjzZBQ228OP15W4eDt3HQxQ2VNfKdY6UEz3I9rA1haQfUKI1+J77WEXplWuGKxcqPB+cWuqErt
69SW5t8g9Sn7NBelmZXv6VoliOfDKuqihQIvoodN9naDqnN8IhPEU5Y3MvDYmfHVVkOqT/rByLh7
6pXWKRQ5r5CrTMQhGomUrx7NSYFLfEXWUFjzVeN9kvpR5PtScu/V9zYUqmjr9g9Wo75LPRwp1rZe
JOK3xVC/QV0u5lv4jzt/EYdP6ViNSV/Jn/b4JlKPtIp3NHFILZMRFtWpjzy1N+nnT+kGNxC+Ghlf
wwe25i0GwjYCzCwEu06mo03F6axYtnvPSomchYbfk0y3QW0Gzs0hH+pKxMlIHWLw086rI2ryFRiX
AKtjWSA5iSaxEoyBgaL+uhqmhxVqe+iom1hhc/f6GBq+Dvtfje/v72NqWOqxc9zDv5iryami19TP
sxg+1s3RepWz5AAaLNtVDxP4yGMsvkAm40YqpgnVRbtwAJ1GXLulUMgF7faMRrSa2+uLda7luqHT
Jp7Pj9akaq5roozWGQvxbjzGWBUeIHtemG71wwRpm2+yO2Vvs0YVFaqiQCpassrmm3szkkGg8Ca4
3ArrDpgA+XtTt8KH+bgH/8swTowFeXXCX1pQg+0JwP3Mte26r9uNhcfy4jl/P/YhbfrUKNkgbjjJ
SxpJT4Eedze67wNvjEx/aZHpAVnC4tGGI4RDSTjtBQhSS0cVYadQJwEEuIwfkDik7KYFTGYbatcj
wYX/n3v/f5YgAAKlCpfyzVePWDOomyARXzuEn3vVaUrg9zxgL4Flk47p5ClGM/88QbXjKitUyPL1
el+wcntbG8NIXnZgYnaVxId/5A8XPV6AKwnYhmXjfh2Ee1WHOTBo6TYrlPTzItvDioORPF+2Ddp7
S8kkidQ/EF3rH3lRhDaLQ4JhSKfr8rigmD4xxqDd+EHCo7lMm913C0q/w8XMgiokZzxxHKQMmMrS
pvEuGYeu7CTUygLFwbHptUpvbKybQOc6rZyZrN4j+u3NgyVc0wFVJcgyOr9daVBJ3H0EX2MhRdV3
E7pF2tEZ5sXdrb2wZSlyJHgyX4WQcWldmJGAAdfdDQxxpfwkaB7sNCwPPf/PVwVrwhi11o4Wu8u3
RPhqAlq8dyfqC/i5Qvpupzq/REq0ip/KzrkgutAEiU8qzHAa0GH49rE3GkoPNAcX9Lyozs9ifyE9
9d6YVspSGIqrlmDd91Ukpp1GdVSadg24BmISzrc2rqZXIZeQ1yieGTUOoP2qC7rlipoW9VJrPLpu
3dlAmNF6lSMVcerRo1kuHr2jaKeu+kOB93wj4lb+Y/S/xcrOQlSwjBf3AzDO1Xge1s2ITR113qqv
qMPbd1h6AsN16c5OqGAcvKKO/tnTUzWIb5dfHk4M/7pgRwmr11b+acQx6MmFzNk1j78RznfuqlDc
2WNdgWyh2IzGeP5Vl9Erc3GEGCy/J+T8PV1nqjDYh+PPtcUZIizTEFmoffCZ0Yl0GNFGrdaKbruz
GzSy63CN+pm4NHtoicG3MxqzgLqt4yGp8UtB4CaAKHi2NlHWqVxjCGrR0YmnLNOLh3IFDMhh3neH
nVxwGSBWJouI5ZjbDtml3Q1b1o7V+nw6rCmesv5cuWaUVS+Jz3cDdIVGwNac/XBxqFIwI1ON+/wD
GgXmSE3ts/71ZtnN1ZALBN6Bn2Iq34BQkuwxyw3mbYDVmbjtQORqxCoqjkPnTYNQNZj68Fr29lNv
8gPs2tLttzaCgMvhZFstDrLQbvIZ9IzJd9/BfyDCfURGMaW2c5HLuzSsLVHmYMdDvdzs2asnV5KZ
3n+bHzOd1DydcCnnc+sf6m6p65gtGfLDgzXm4tCaK33KpbUQGwLfXO4mtivpRKki06B903YRPBkP
9KC8ayIlMMYiWj+W4BWHwG42f+UuvuLVXi0dZzaYMdQcdg5RBa7wxGrqhQB3CxHTb1IwKZ/r7HQH
qglLgr5sN5ilpPF1WflqW9/MYz4QEeKODFIz/0ggQoVFiA+nXik/XJVE9wff8eNxCyX7eppaymDR
05kYNvDmrHcC2nw0hZXhGZeURtd4P5MP94NvtPtXgsgejaJC6xTb6h1V+iK0o5iSxnKMu093609w
4Z5aOA2+Pj/GXQNZPuGUf1F474EOKlFFF6pRHsg1LSFjBz1cuTsjj9EXDJjAj/sADbz3EjTQJlOb
AhJfGTV6GA+x41vPG03dsHdcdjeNccB0jnkNauHXz89hQP9V4Q+zcTcH7ofX6AaHBP4TxpwQJvc5
HVRXUa/WrsneRs3Noc3z9aV9WCwwH4lDsJIncIQO+z5hG8vkJr3R+61KnD0Aj+svhWtBR8eERkTh
z1WxdV1n2IFfMnhK6ruZbxkX6ROxOilizUbM0Fw/qtUlASlZzVtpug1s53lBpbYIbqVef0DnSdJv
y7HQQFuE5wZ3C8dTbLWC+IpyYOVJxqZpu4GrRdRxj8TbIKBAbjnpD7qCppy+xo2tnv6Wzm3dt68Y
Lj7faqxNP+1G4KMXzO6PpuNe0cLXhyht2UEgx4e2TJjdVQhgG6bIqUKWnJaDrVAHVE8Y8udAE4aE
OgWetzfuUdFYXfIR241jVgyvrpsLhyDg8BEwZaa22D2c4QmQ6eFWkT/1zzQ65C5zhk+Gk5RQ9qKE
aFrRKOZvD5YYVYOeBWQaO9BXwwjWIWsaC9AbPdDdToHUBKAe5aQ/3nNt+PVVPmVCa7P8t0NkNPc/
29jf663xadzDQ+nvnC1IIlRwea1sDtIJ6fPQ5j8gD25q2Vs5A/WvRRLo1aHeVX2qr/4KHJUoZU7A
yb7ibfVTzpnmfHdSRawtshtyt1j91yrBuLbLK7WYcetHlZgtgNhLP6rGr1p5+GKPH0BPfl/iC9Gd
1NSvQsgKV++MkXzSlwosRDAERbuUBnPluygBCa3zLNtjf2QFwt3UWTFIHDAKysclqvvyYWiVTQFv
I3hMuJJDn7SxTq1Ms2wo1NUWodJp9pvSUektunslGBWjWBO8er+Q6OpGQnLoaG5+nEy9wxI/i1L9
RcxEOzebUU+GWctc0XyNDc5igQj6XWGCkjEU/aSoYoUIVwfgMSiZwx3tQIAyvj92jo8F72bpwLCS
0fSQt2VWUVI3eh+6pFDJ5z74Nb38P2UiR58K+MWmu74pKG9uzx05qD5jWG0w9IHRnWpztp658nyS
j0kvs1it8FGH6tGKHoB/iF0Zq4JbSXRsX0nvwxL5fTzx3BIetQ2/zIHZmZRQA5+Nsw3zyFRjSTBf
6NqEVGAMN8NcdPJfuF2VYNxkHjMDVumWCs7uq8RDODmNJ24wM12YPafECQ9arfng3DOjGsZ8kNqG
8Yy6EI6kHtW2K46Cx2wwDAxgfRw5UT7gxibczKSPy/8haSQhbdt1BialU5jkr9YQ6rwBRUycuRWl
wseB7db7LArlwSaKxf7PWoMwGZkoy1KoznyBftTxDGOo/OkGe7zAQ0Dm4TR7AXV4Cgx7Qbc+kp6+
9pEZm/izyVGFYnItL1gK7Qsm+Z/qXKchHUbN4f65zyCzBiAzIS4rQbIbB99mIih6KM7dyK4jL/3C
xfqFSun5pPpK2SjEz7bhpNt0d9Jg61lIUNd9qFJmUKL5h0+7vsxixCNqaL0sQvodaus+9V5IFPmK
Mb+xk7RXgBTWZ6j7vKGkbDl5+uTf1pp4VzsWlx965eVuHF5FjcdRCdkxc1tXoQfq5wrqOtMkuu3U
z7IdZJhoTBR99phwP3apEjU2QgwjMFleYPosirU9LCdD/acdW3+r8G5GbQ+HnA3eQam4qnlPnNxk
ro3TGwn5brWQngYtV9K80yziPurR+BrpqgrBfz80n9lkd8vVSyn5mjEZIXAKJxxyxCk1kchdeMPP
R8PeOXzuvhNcdJEG6b0hzpHEDqRPIOsfax56okZLooMld1hyGXrKGiq74zO3W3rcsWvOxx1CMu5k
iQCWRMBj2PpS9i/Fzw7bgMZAlunlS7CUFLUlrr1u/euA0pZjV4eM3vVy51Lt4qH/yToBSfBVFvIh
f7U0pk5jlPMkTW9n/+TpuR3QzzCpDjH3XyX0rgYlr5JlMEA1bYpa6oVof8roc/iLw/YQtlwFXOW3
MF1fUor7JaOhw7bqRY1+DH+GOGWnEqYrJ/jRdDxx5XPat3AkoyPmEa8Yju8Xwzvv0gteiy7XOZwv
WmOqhgk89+QMl1HqjmS5SriZzyJQTeR5qZ6A+Dih7ymJ9ysE3U/G9IzAR2eRI0mzd2hR8rrXFzCg
MQLLPKmEjzORNkMEECm1KhVQinUbyBXyj1tyD31ei8xdOzjee+L1P1xF/QuEcDAZOFWGTm6xpt+q
KVeNzMgqeXNh9vnBi184zCZvpaT4SYmWr6AeEVFtT1qWhYrBU3NH2dauur9jnpJNfb+Nj3x9cMxt
uFhDUPZgS+QWiKceRV2dT9t3fbK8B0Gb9n5hZFjA1FPlulu5ZaJncQVS4Orx5pSBnp8j1fCyZtar
7wtR1OTH6V62xyc7J9n160qND5LLN3EfFBUQcW3Haf0r6ED5FqfvOVQ/I2t7D4lvzmD1snp0VkJx
yGUaiPVkfsWjehwImS32l0jyopTuS53ExI3Ea2KHfsYGdF2fv65AXsZHxqhwL9qyZ0fM9eAMp6um
uF6uT9ouNR0RZh+DRwtFsLc+fCp0bEgQIWdS773O0B/P/bJ82iowexSrOz1fJU8sH6XYTzGtomTu
RRjc2z8OrIvStCZZZwvyha9vLkCZCPBw/E/uy7vQX1t24mgZ2XybxuE5VYd5i2Wu9Vts8V5rHp8C
jZ6ZYWCHJZZgljKvvyBW1MAqYVWwotbSBgeg0nDs8SgoUHiGOnkoSTzH+DZZZjZ9joMBMwadR3fx
ExvFCk/H2Bbr8OdHJYA/vsdDOYbaG8kXXDikXXFduGQO3uobmLlz6bTjBAh9loQTY49BtSj/NoGm
P9aIls/OtO8UsHrx0BRfjZpU+eFOwsyGj3zn4PU+CgY8n7y1i5ga7uYukL7N19iC7IF/rBtxyOWs
nts+Kt5RrvLtHv/gNs99JB/j4JsBO5/QOVo6IawmvfwuF5PwYckWeumDVxemCV61vI3+fT4NSwe6
/CBZXaW+XGH46TiDh9WfKhqlNjDnm0NYyOqdmyXqXs613sVcyA0thn24eWV2fnuKY+qyfs14spVn
IK7Wnga6GkCtNR7c8SthFZlFWOD6uQ0mlGKXGfzVLNR8NDSIsWrPh2KwhtsAC3fiDS8kppCfHtxy
t1LEH7Yf/AoMiHnPARM4/48Fq2LiEGnfa4FfVBVsvxDmJdbJZ4FpYdMHU+nFWNtajsfAXixUcbqa
tOBf17ervu+7jhoB6rJPxAqgyUGdf46tpHhMIDTCafXC+f19C9UTkB9693T1FqEqmRteQOIOd54t
G7fc6U5B6HJY++vNsOmlPnfhmQ/2fN1iElaVfpZ35u+AiHeleMAfXeD2WSrLEkKBJLlf0oBdBr/J
RZgwgE8LF0gESh32GSMB0ToguxubbJbYN+SMdtscrj/D1feawp15zEIgU6pUAzaXJ15ah3/Mf2RZ
qTteWb87GeBIRdViKIXwSsCKdznH8B9sRyh96/sFBUpk9upKpmMNIgpZR8hzrufdLlvTbShaQK6w
1H7MzOW5zXRw+x0g7veKs1C5KIpaqyH85y1CIIOE+pcKmvhmdvkNtv8bPj4lyVmK66BpucSKk3Zw
RzDPLVnMK/pBByALRkT3GHgaPk6CVK1squh7IUlLcLk42YuNb51qHLyunK1pddJodVvN/iHfSRnl
GYzrDBz5KdMynwTpRanzAoYUzRLidHOwDjxoUTzzP4gAN7/UrrnvObtUoF+5pLxqIWHolIyXRHy5
+rC5wOnOkWY0Ja5fH76r0lQd3m9OKA8J7wQKe7fWioWCS5A2aFuKQlwTLxGkuhxWfxuNeO1HsZxS
vm+Nxc4j4+O/hOJc+uJ1/UEmqyw7zbZfHhhdEq1rofx3gbBYyNJC/wMovgQtog8hE0DUSvzdvbpP
fN328PKPfkgsGetGAwBFhKmmgMCB4wzRj/goZMG7XjSwfYzc+wjuCYHc35rQviyLLN2iFWhbIlbY
Az+NdO6LKKY2Iv3lQ1+HTP6k1ECRtVqZpbdCRPEfUbiKkhTj/lGaT1+y4JOIrKI+k0hQfjiD1F1Q
+sn+ITYTCygvAtxMECN9t27Ed95nBZAuibapevnDJ9of4JaQze8CuAEO50ZWIERkVtn4kpAVMQMY
jEauiFHTUlNB0TwVe3fyGSBhCl+pM+GSqwFT4YiRC0KJ5CGuDF9whAT9E3Y9pkxwETPyTiM4oI97
hQcvWJLEEfa3Rgdtq+Z/DHUBNUo4kuUnQ2GmupvCRZf/uHbFTLZDv1urJbvpWB8MKE8zrfbXOIWt
gya1FpGmGfWRAuV/amY3w8n0WFmEqTtRgYrIU5j/XaNtLsloJgfKkffqb1xZnp7r3vUPygKsRTXB
pkqbhuevKYqn4bchYKvF9WrgYDPG4m0Xy+U6WRhPriaOBYSiT07muTuC/t8eqlTdxaKC+NA/Rubt
JQla/iZu8sVysYmQGEKKkarTJjQyHlutQyXPp5QLZknZbeTcDKO9rmVqNsBn4zNk+UhPqI+p5qcU
6+vNTNy2TS9c493sb5SQrtQYaS15Q9OD1316OHGwx4d13uUt/H6nJp+hIjJsP55TC5fxACwESLee
63FtYXUczvOm9eRXhE0hxjBmOYU7fMPnZjR8M2beN51PNc7xfH90OLoaojZw4sQoA2IHpI0eW7ND
Y2I9t5HktRSoNDrhozvoM6ft3Cq9Ax4kclz0dWvWahWHikZcvxz4vuR5lim5DCo/xcC0JnE5W3ja
L5zf/X9gyG6S6ALWDENQN4jPft79Nl5G1Fb6rliVaDdS7CfPe4NkQUIbdowHnpMsZMraiBma7VaC
CHMdtOZx4Mp9wadvStOu7KQDHL6IMrY2+bo9Krk9FHYEoYlbfYAuvvq6ldg1MTESH74KPpkwGqYy
3/urkaToOLgHznZIDwJmtCia8J9XeFHhWrTWwXxWFi1A3RSPvjX3fFICr5ijzXmGOhxrTWOgfVDu
70SXliqOvgXHjjjf4dQ1NB3L6l0U0Gjz3pwUHOa/WWHN5FZbDUliG1NTrvMfU7VQ25kSTNoi0h8D
hdI8r5n4kE7sg8Bz1BW9VQMepAoU7RM++TrtUW508b1UeY9x6YNNXmEw7UuWM/G/RNDz3RUNT9J7
rerfsLk7NZGvEyru+8N49gsne5YpdbBSJupgma/zb+5MGHdsCqLsvqnW8g2Gv+4mbt+8zUf1bt88
ofE6Hqo+5hN+rnyJdQr9VUkBA3kgVAbSkkzGwkGICy1ODWOuUBy855XlJiIonTlUGQpLCZdTzl5N
9fNgwEPObIuOJ6+cB4cMH9Kh03cxsksyJwNtWvhxPLziDwPpgWjKLYgc/3KodEuJ6u/Zlxc2BmP0
YacBuXBsY5w54Jk5L3hX+scAzQVvjP9UZZ3r5i3eErk0dxM2n+qNZ7hsp2m1/l8HR/WdrEyrzngF
blV5wozoSjEodXcbGBQl5jEgMwpZlncP5l4KKjqKXQKYz8ZwvVYQ+Um/7NJKOrfg8KSfiY8Ri05z
YI70rrEGmt2Qsalv5QWXhstVlE1qzi+g8VtAyogOUFFF5njmjDMdPOtELWfUEOf7DAZNoGOgeO7M
Z+Zk6OkwOfTFcbOE0rfkpA2EgIGlVmVR9P0mFkiqnF2cB56oDi23oy/VPvF3m6WNTiD+TUeFISEe
WR1DvRGxRrccZhHdLFF4M0O2BdWF6BAf2iX45maK9kRouMM3g7u8EnNZautUHQwCqQjWobbUA6MF
cegBnD9RCXaV7OEyH1sugsFn/kLI9fdz6F/a52NCEkI41XpeKiXcQwaADcs+qzSJNF2frkcxZY/c
S4bGy1YmhT0GYLjQkeVV3L8YQBkIfqlUttEH5V5erPhNrB95vscKnwOCLBU3YWr39K3SzTue7m0e
/Jj4KupruA/d7nCzpV+qj3BUcO7O/H7GzZz3CYNHipDE/aMQskzaR28TTDQwymT72ackUrO9L312
+WFNjBhTKWu8wdaL5gzpBz4emzt5oEkF259NG8rTYKyF5Rbwrv8JHdn/ZfEFexFvfvkhQGrJoNcQ
yWOK7owrRFB0khSjrjc0nrZ+PgqNmNPMn22Awp2Mbj5czyDK+qDB0lMS750WkBLnpnOUgKiW44cs
BEoiFjiJGVoOKAeJ8ScjAjaunTN280pPyGj4jl0Mhq1HhHrE+1QcXonZvaYb92ZEb/c7VhVMZbDJ
xGZk1xh43C3ghQZP4Bh9zaJBLFl3NXAhr+uYsZlr1zQ+jsQ7mdBUaVr1dd1mzHCfzikRAIdNYKb+
gYGsiiV8rE6KvafkIPgUkVolBNhNbv/EWRkhWmOYnmmpFKO6GwtN5JQ7wDDWfkBq56RP6F/oFk6u
SHgxoz4OgM6bYJZD/XV9s6RQjIMuzLaA/xShX0lDuutOXVl0DkXqnVhcTxxVjBPB9NQyFYzGsNw1
gwYQ9s1cNQnXRVsLhcLXBulI5G3XX8r64fhsch5CSa7vB+wfZl0Ck3YEtHmpYelwvvhNab2KpGRV
6JwBvOQ6qwAIVC3jj6WUB0LM0PyI7H8ivSdz98CIHUwPlVEuufMsa7N36HmMuEabjzqmEYeccc0V
3EJd7krRlU+EP2qUV0TEUBFZv7KcLE8+BA/gL3K7RZNfkm16i3EL90aVR8UiTuoudS2JSoqgNcwU
hYEzTwHTiGLs54TUsjK72rFnUfDVRcftZNXCfmOehV40KHq45lUCZZi6aofFH/mSYnkr1SBD6erY
l64QPDi279ohgbo75K+YE02LAu06eYSK8SLe9qO1y45717H+3TANGY5xBVeFIHWrynbfjmQZfJiz
orcYG9g6xHi0gJpcQlwnF7wgUZoi/npbKSWVgdKDxyY/KazU9besc/kCU2kMddS34bO4hqp12js+
xBXLS05QZ6ih5s7epRrD/wDqx7WQqcmmKSuNy4aCojZbQ6SwyKHcOrTOAvXrfJQiIEpZsNIQSIs5
gmUZ4yIjP4cS8aQKkUJm5YBtFlPlx7IHDj3yBKrgtCBMhzO2fxFuOgN9GlCHd6Mq/xh6S7nxDkHy
D52f0slxBFIZt3hsQ8umrXRe4A5mUrkuGGZ5egUXAM6xaLSi6G5e04AxbtDu1mgVR9NvA9Ux65w0
N2kdJxS5NW06KwbbnAEUy9Ow4vGW4iMUQPCH4A+RWGF03LD53TERWr4rEFL8M/7glm6Ca2EY1IGy
HPjWLuW0ptVFBV6kejUfe3iqCdqFO+c6oanJr7J5y+dMc3Px0dOycQteQeVaBLazfRvR1PqCOBam
xRbThxxsPZtk3TvIrxVTZEFCpYBGiKAOWIw340Oyx7NQRKi9zticTXAQHPvwbDZxwnInlOfNnjor
oPF+EAGYMU0Oe178pU38mpDlxn02oLZrMtFc3eAH3WEDFTI8NtgrIT5N6fsgMKsjuhLlBvXr1x2i
YMoYTToNfSCOEoEoEE0K7ZMFzNEn4HavQ/e7cnJVMQUIKaR3B04hxHY199idjKdwOOYmpGjLUs/U
kxZNuDYm/Xt+k5ML2sV+cbQwHlZd8O32J4rwz8lMVQ4VjpF5sNkZMymu0kULTrx8EIYdR/7Ut+O5
6GhHBUZnc0RHVjzRiMkhx9wNYmgdCIQ60iPN/WcuDeJb86k4qLWh8tricScwDj8w4ZvsKmFOtUj9
9dzltzZtZG14vx77xRG07cbpml/dXubORyVzdQMoPP+kkc2X01tmrYcGRsvwsxZxdi3Lv2hbaJIo
SnVN4eyTcrpgZ9gSVRGWFgojyZNt5F1gdS76UqAbap2clM7ZU7eAV4GkfOvOskaGSoi7P9DsBkyM
JEanvZHCzFq3zWOGpepCAC0AWxmSMAHGF+64oaUPxTRg9O+WlkHAN5lWMHYTvIiSP97+eSemPHAf
UB+t2RcU5mfs1bUmOdux5Cyq6ZSwr4ZPVAOc4yUaig65aazU+K1ZpVK6GwW5DkfvpI/6/Y21vM/p
PBoA7hjYx+gqJEDZUuns2nPZC8er4Mm2eUzjKvj50a1BJxidqNiym3MHwhv4JXEvpvZyo97QNnF+
eA8EfJ9Rmgor4j3V1g30P97dRyvpThk4jGH9i2tnYMpOqs8W9gumDx4fu5O+lPt8Ewc/HDZ5nKcS
73uAhGYLugmSNS9AhqjIfyw9EhyuECacbXmfG9EiC7FQIbu5yFHpcWwOax0aPkkEQymgU+SlSONo
wsvALfgrt5VccFZm6VJHvPTk1Y287vrKseKbdY2yI6L5TuVgkCqxeesjFsjg7En7mAxFOlCYjbpd
mm9b6t7Mt/yWKBt8Q4e3L8WD8QtJ9SEMP04qVeo4L6d7SIB/wUtrqSCObv8iPsoOP2eWPeQEp+bj
6vM7yKydE60X7wTULiQHI8dfepP3lYOoN79YWrl4TM2mqicroBSUXQ3LV0b9nLJF31C4pDefklq+
RITyJpT80ZGMGdI9XIqIZERVma4OqRUJNnjUuZmnj4pwxMqet9I9QbYvwVLz7B24BTZgurenkpSO
RGGktEcuXsPwOlfXavbf2KWhLno7dd6Bw4Hvykebp+DaYEENeQEP/PVthhL+dm1mVBaLNDSAvBXn
WLrwFy2f5pLfb9dDSfjNYfaYu8ztEO+a+VRspHpSbNvQBDsoJJZUJnl+sGqVN7ufBQ1dN+xRPueE
jkkgl2Qb1XX2DpHJNabRjMPncRrB5B/nmcQUPDldnqMuxre/fjQcZ8dVtTvD9Mxc/dNOs5+Q2pZP
T8cxoxlmI2oJdLlw7LofIHrHmC9QvKqXJZGVdvib2NJQUw44qYLw0LSAmQPMcDRBbz39/wx5s2Y5
Ioco4WblkRdb+O+k69Ji/82zLll+bpjFhljy7KG2lRrZ61Rz6y/fcDpKRQyK9vAritYiq9HCZcNL
G28Rf8RHGhVPRj0ahZ1Or3+PAqOYdZRSBw/i7jnEJVFGOI+hA3ebhsP+OLgKxD38oYxeWxtP0yOV
E5uWmaNvTVrnOuKlRGSU3DMMhAmFAQcfIrX8/pElxf9NK/3ZrNOCLb9auiI161rkajEsD4CtOW6k
UgTFulxrjj5az6BGRHWYkBfzAFzAiIC3hGPMK5pQc5xIejrl4kE0E5wZuGCaodHs+jVd6Zp69O0u
AfmpptxR1uOqKiWi+8Q4FBTGibwsXRoIrhAsjsQ7zgiZNhoMB8G98kfkFiwMbxZPmipnfRBfZUTW
gSimQNYWs4yRqUtESPZphiL3Bt66latTkwoZBHQVerWFBaUw6KkuBkLfBn9xwB33J3Df2rb/TNTk
aTeh1TYNtWSXRjUbNhAMVhdKRHPtxRL5IzVU6DpXLT2GeQvgwOSerLartYkwv/YLh/xtCpLYQBwJ
0wDJg2N3mq/NkQI/gvdJDPiMNNnT5rd9Q+DEHB2Yc6nQKa2UOyWnfJ1GQlBMYAKy+ZWkZb/bRE7C
fL0iSVlbdDwlQbCV1yGf6yDG/jYHEPaaRg/2vtN/GPNyPhwcuEswSuw2R6lGQQGSwkXdJqgjaxGx
d1dwJIYgS4N7/EQB/Z5QmhUp89v6p9quS7GVpzLDOT9NEKBg82Wu/yF8aMCUBNIHjj2sACdi1CmJ
TYcr754X3ZmlTHfQXXtJbZzfOQeoWLVf+NPIlqRxxai0QBLFTo0kTmgRCqaINcS0ltoUrPTy2A6S
Q9GUk+LgWsUUFWjehDkhvV3kr5ZdjY95DcnB6QGQUyXdKyy79wWLiTXz3dorHhThy/3mFlCt6FVP
P5DHxBx1y70JdmQRFFq+Abp9jptwMZItC1IcJkGcGiW4nfMcnubaPpcwx1mRSdjByr7GuhsfqZDa
2M/qRBd7TV/42ds5RNchzJAN8Tsa320PlZJCGjBc3flv9kwfF0SwlZHlHZG6xpmmmatBVKjyo9ky
18KUYhmjIUEnvomNrtCfJUTcOJf99FuOoC33ZTfFNwfztrtXEK4RBxyWoucLL5vPVL6dHZ2TRRCV
ivy16WuU2WPNs61vPDjW2aTy9UN4fy87DGxhalhcnoozU2002/dbBESLmxjA1oATSUWJ2zbt+UwS
ydmxunQgONPbzvLplflWWoUwqCeY7w5KoS0pLkz+iY1tsivVIzhYEJHewtRL3nOmKGwQLzdxBCoT
CO8SPT6h4Cvf/ESjR7PcAmMo8KsTo899kh8ghTlFQAzBAyCgQu5IyKSslQKOeAMNhMVVYcqpZH14
hGo6Lt7I4fLyCpLnTRcNgFeaAQYCBAiRDPupgm/BYdD3pSqSJqhTtJ4JHMSBSO4N4xv7ijnvoQCO
BLEqMab9wtjJ6536kAdRsdzBcdIaTy6ZSMnBTuGlJFHqcXRXbqqTnG41ms5hnoAbJ2DGzUtcCcc9
rkjUgqepZEH3LZzKio907VyaWjtud3EC9jm8q8w230KLRvDffF9kqA7LN81b5Pa8X2Flz3WvUibp
fuVdCD0n1iPiSOIJeQFAbSZc5pH01p5jiYLk4F9upCTPjMvHvV8n6Ab1mlFaEj6Kvku4Ip7iyUSX
MdioFf86F9F5ZbRQ3BUyIMez+ejPHj9d1mjshFCpi53rIhhrs24lvvLm5sIE/mktDm7FxuMb7Wj6
bDuMbXAYyveUGC+tDptlkunvItGdgKoU1KA9l3+W7gsqWDSW1FqX4qRQQwnQIOgV/Q/OU7V/UkWK
NjJcA+9UKlce3Ngp3k9HwzIp/lxqk+5Upumi+YA9axB6FsaAeoWCurvs1JRUn3Ng897Gw0lfPoNM
ZSEx7s+7aUK6EnPwvpyAtjZFdjjeE1QLAKMZykR3QZ/TFA2b2QIt1DKH/Sz2QtmSrbb6EgkrZlnn
A3pEbHndW1dxcFYOXu/Pw/2+ZgifehHxnyBsuDeV/eFPjuIuTNJNtMhSIDSlystq5fqnGGQq/JVZ
64w/CeuQSIYwdUGDyFSGkmJNeaNG8WBxgdDe2hdtZfFO+/je97XlLVAMeD4gixXgne5jvZIUhSJ9
JIgXBqnWMBBgPBsiiO9G9GTYmIkHIbj45w47cIwNaVBT2v8YO4119ZESDSvOFxaxBvWbsj9glOK9
nmoCaM1e07YrJqF7uZtIK22a8uTgHyQhTKnl5PrmI88KeI6SFATedzj+eNyn1zQLhaDnpCgOMX2Z
IfprUJT8bXy5poxxkrOYp37MyLIC/vJB+25XCaidXeLuJJxjz07J6s8VEVL1nU1rlJ6n8b/oeQ9h
hZZknW3lIctUk+fpiO40HtdP1Xzb9oADZUgG2KZoxAq3QGlXPCLXHU5WgEB8bIqdhw4H2kBxETyN
MYEFIZPcKKMJa7Iced3p3w3o6K03aPYHDQT2ZnFY0hhZbeIXPnbzoGIjSWvudf/CZk1NfCR8GgyU
w1w3S1G+rJ6TOgb3aklF0LaHVPDDmrJ+y6SLgL7w0gsY/CfjwYQ/hFlVnw8bXPvz3K2DQlrU2d2o
zy5oZUBWaphW8ZwK9e1EBohGoRGLYViAj+aLIwTx3t0D+OiOyighQbSA91w6IIdiVY89H3O30p7J
yQlRNDyaC8Bku9f0rE6NmqsaBtgVqwOMiOpl5h+4Dap61zucQz0D/Ji0lLW9Z6ZeJ8Rbo4uR/+ux
5RnBsQNmakM1si7x9p33TdOoc1PXWGOJs6OFBpAV3lmuKovF//OMt4WD6FWbcHrjKLCJZGh2OR30
NFiFhMTRqASvaoh9Y9NQbl16VocEiQRb0ICecsoAHlBPdeYT4ei86ke5t7gKGdyLN2YbZljiIETg
97EOg/VCqX+JxK00w4hVi1n9RirnCgzEVBte85jGL8DRLk0xTpA0GJwNiheMA1xWTO4Biwk6ufVH
UkwSLL452Ix8s4mX4L48gmgJSrKNZnPhktkcheRopZB8ZWAhyJGLjl++xPhGUoulV5FrEs235zjQ
1WdogeVYqPcVsAzNzXg/4e8Sz9obxmhZt/KGzFGFCDGehrE/4zVOBfQc5z8okfl/sTPHHoXfaHSx
6JwfuErcpFz6dUvDuDAJvz8vbcOb2MXPUv9lUL8JgZBrhS3ZlL3CIaHzeXFlPWsXYJCPyqRIV3X1
nAeTAxFWLSn2Fi/Prxk14PxZpK7ZKsPQPeu+pMNrbFhHshPZUXAAk8lr3Rcusg37Pgn2hUceB27m
jeXtwuLvP9TUvPlvRz71YlMNofmRRLPnDdV4jKYS31gyEeZgXDUZ7ra3vpZCa7iUcxPrELMSAGhf
2AkdKSWNVFgDK/CVl3olUpWuD88ptnyoBKXG4i8FCVfXJM/6be2CdrL/0oc1iJRd3WD16Et0S7zX
kBkE9Wg3rKQmy7RnTcbRas0Zfy98yU8W+KQyVj4bZ0w7Xdg4nq4PDSPrzzaPgKZDZTpAjb66SbqM
Wq40xXt4HbFkGlmYN7VdBWdbL2tXYaLxUT957yjhTyGf1zxZYqUnDGd4a0t+sXjB9kgCEobY6+T7
DmVsXDR6RD1+jrzVi7YCzPYnp1CkE8CA9BDeOwETKJW0VQBcKC8f19el91w5ef2AF8Sqv3XVpZ4z
zwnKgJ92A7td7K2iVn6DakoRsw0U4MRl/YbJXvctLnE28mzXC9Wy89UAYkQ6HXdr18mnQ6qFLMAY
wDzgvCta1yGnOxLhhoh/Ut7XbvimnAGjNg7E6+RRn8q/m3oVa7lPWZJRbFnERmBWATd7y1Z+nUxr
FlkjUFPqb55Wo0yVhXwt6W8W4SYQMLmuaMpcM93sVzZKZCwZBVDGWdHYYbrhHHCVU5mJ3U/A1zDt
G0iunhX+N0BXAZHUol9rUm3n++f2m0VFTtRkyOba2b5kX3wr7Ao0UzAMplEHxqiy6P4aFhUnWpOx
iC7D/Hg1KPg74LUHuZSMANMgNccvw4gZbwqg16dM/w7Zr/7CAFV3dZnkMr6v8cCS1pzitnuKuavo
E4jx44JodjRlpc/i3CgWZ8MmdwOzWiAKbmMmO1QsFQHsm1LCrCuMsW2ovQCBVpk8ESUDlUoXQjdV
yAWYTi/haNDkAA9qFoeVSFqCVwy/t8Cw1vKmZUB0ao8C1aLP90eU8KLkSMIn6GlRwTbEgx3weJHi
cdBpzE1t5NUf93WBZv56Al9tUBFw1NE6qTIj+T6xt1E2Yl28hmqh/X49jSxLyAVydpSh04PxkxoR
YB1fxzbvNcJB04Po4ILfGKaW938KuioD0mixIFDZGt0DfuVnQ9fHQCMYcwhHNtYp/aNrsSqSW32b
7abREbhLoaRFjpiPgl7b5BSucdNLuNhKvWnhCucyomKi2ml7VXNQsrAuDUtR9I9wotK+4K6O/zxt
0WC3Xiq6Pd6PPKRBRfaZg1d4PNbZvfm/QcCpQ0FpgYAw3g45d5IXkUffOUOj3ppFzhmhC9rGq73B
qcORFHmNgE7O5eqkWwSs5OrRY42klpG0rqMOG3yT5woXz7dm/yL/qLkiOfkiM7Soy4AkXEyN5PDV
9hugMhJ4RBBe3tcDxNRS7HLswbjkwYeTKtO2/jv9VPwVuQNZgi6yFuOVIOuHMSMoP+tEeAURMbUh
0WJtz8T5LMu09j7zmqa+XgHyPFTIKh44JjnaE+4Tx99fyFg2dq7I5imssSVvzlIdZJTWLShMxWXU
TLCxmEv14CDits4NMZ5YCoD3FYDcMOnnToScFfBpdYtb75/aVOV71D7L6zySnucQ89a+WMIck8WB
2TD2N+TC0r7JAWVEbOS7kd9rsZ6+N59V20XWa7/Ku+ZBEjXXENCOvybmEw4lDfqZZSbL4lWvlgqU
OluXS2Et8r1lKA2kNQ/veuoae731EVYp0F6VcMk0eXOZBL0Tmwx/6a8mqBif2/secTBY2LMXITpq
+7voHg/uUUeadewy4hkpw4frkzmwKXH2ncNokLqmzQ5KpjEvU2cISf7hUKwcpRtZLOsgZeozCoec
kjIyGLobNTiS3FVDlMnKFDYRFi2Fpe3Qwa+6engXyL4yBf05twDcCXxqkglXutKqtHI+pWkMTRh3
6yDBNnIlKph3cMTTsorPECq5GalqdhpgiyrDMif1pDum6CTRq5IVM8Iz1ChbK80onB5qfjMyREUl
w1jIUsAjOCFGZm5d1ERiIgBp+ABHgpf0KkrsMNjk5UsEFdOANNFUaKWu3NB+2v25gfEQ4Io/ZzEa
tgIIondvVGRWfTXbKemUsxiZWRaSEhST3xTju5g8iQVUm9/AB9exW91oU5tSSgjr4LnZH1ECGE5m
SJ9/I+/N7bw6jsENMKFCqEwRuJLGRZxtK6K31Sb2T/0JKqH/ILgYnqkswLHCTtJGJ2nAzrDWHxWK
8La2qxm5C8wJ/7vPp3W3Z3D+r2SrYRwHxKAHX0+bSnlArmvzblyBxTuxwiPkaqXoEvEn3Nuyze3C
YghZq9deqqO/DSFcF5ndkWYkA9duGd2b9zyvRylyV08DQlK4DGSDHB5tqZzmcC7ruyWVCyiPtzWS
tQFVwpLcjBgzjTFXDI8pvcgU0hnXp5FeORECe+DHiTJcmH8oETsmnVbNvgc5JNDb5ut9wM+/Kn2Q
gINPc6AyW81KBC0V+bqZzqEI7xc6aXD4tV3JUg2gLBJaKBYnzDw3thWPedaWMVNk7mRGwYlBIYj3
/FrhRAhzzQla+0qOB4U06JSVkUv3+6b36a7aOfSRYrzwAwAtplApjEYaTiXtjD3a9Ote1TDHs5dH
thBITdu7i2GU0q8u4cTHTsIHAndGXiVjT/s+k/B4ZbpH4bPEjqIbeTnf7YH3EFy3WnKNwAgKJrYi
4fEjS7+hCB3Kqz6DQrJvr75PJK9OX/P3QcWxiwAX9ePCLnsgRc91dvIF91UZenW87kg7x44sKP7R
st/5Uv2ni5I7fb4Q8hkooG63IDLIvVKeLzkQ2WBjcMhyWy6VfFDIKNA2Gb6E3tkihABJ487I8uty
hiAEjr76jZ5EqYHcbrfdS87F5Csk5czzPWwWlV+tUgVUkPZ3R8shPgBxYy3DRxmiS330TYE6SQLd
OFzLgjcuIn0ovIi/M5ZgOcYIMdKnprJj6wD7fPXnzrN2N7OgGEQ9gbBBTkO5zn1615SFcWckhqhy
h5MsdThDN6drDwN9Q1iNffEDn4iVLQnlPSgDIYSUIUlxAiHrCjhCsDOc+ytIyPWwAiPY/xv4RSAv
deSYNYdijjrEQUkuSXRY+uKWj5blY40HakBQFWe25KURsiYUfC3ccK1xOyr6UxjPZ4o6Zt8iCFVw
5XN1LcqMDIubVqTY3PeXiHV0CLXRX1gbBlx/BhrsrwWY9gNPOVfwjb7PjT8vtC5QT5b04MFmeG23
KYoV1gYZ0FlR+8apwK4sbXXWNVqUHr6H78t4tLyekJjw+0buFepLlSdoRkmNCb1Jin06cp3xg8Sa
6dmrgjh0nqtnmkhVq8ncf3R09bZck3mjndCeHLNoHE5QdqLhOueH4AaNOOZ7D1nmTflYiXorSPhE
Z4zwSoOLWkHtn8HWzvVcBXsWFU7ZiUMaGr2a76TpNqwZKx5bvbSK76+Kjjkm1pqww8Dio/2VVaIf
JureUhU39+27Aa5wC6iJgkyRG9EswCkOZIas2vwvjOnYjr7+og3WZ3PEBuBemlzABKKOk7zkFkQN
Z+Rm89VzmbQcAjx2ib6Xdu+Hxzg1AjjCg84Sqn2FQh7rLuTFEgnVMUQbkKg1dx4IBKcg3rV6TAND
5fJ5xH0NJ4VpyPTFUD1oKttAQeXb29BwSOIa0pwERVdB2rADZfedXKZxtMxM0iiBlfOez0uqNMXW
dhfyLeLunNWEYdIma3YiK32FiQRfMFwfGOkMqoEW4NL7Pv+TYuMArsPDyBZxF+0D0xfqdqRhJsx+
CkzuZ5DkOBnvElj7GcO2vmboaSxT0WR0P/oxmQ5qyfA4Z+S6AVS2WFVuC7KDdXz/f9vuOIqQbY/T
3dbbKpYQpswiitsfTIFb5+emGnubPz23vNcrLKa43QDSwT1UlFL7tNxBpr09VaJwky5LHPHkgYmw
XzA7aW4B/s/Zes2+vFCIrnteWH0IhwzoYNi2WYa6BPKNQE6dEFkKlqTYQhIxDATfmK5BL1zxa2Zp
pbhdIFW3Ox2ZgY6EvGWzXAvlT/IbzIROpLfgmzyI4FrFUsBcTc0TDga5Iqz/Iw06hATZy63pN1C2
s41EB/nZ+fD5YY/BDJAPiyHoOhaulj/K3NqX495ZSZrcouuVmRLT6aMi18VjyF8AZ6A96gw9OC1n
K4KnUxSAXqnbSQsFFRkAX81WlM8+vedEImldlOCwHasXU5lyxZ/4v8tdmsBOWtMfhqKKrm/BoL62
9mak1C8ZZ/pSi9xM9jo8xNtfaDVr/0F5LN0mDLVoeEZeHPUG9xHVHb1MRKlrqqKH2gviUubuMCDc
m5m6Ywu8MezxkjMX2mfReJPC6tT342jrTl1QKokqIilOuOcyZh1j5JVsPl6aFe593gJtIgPwbVT1
nxMSkbbNOpu8hKbBZN37n9Z3AVeIhxzicY7NlIWFyYgHKPSm/0RtpQUZqt998D13EnIraZC3JKSe
TsG1Q+X+mVA8AefRipdCor6gG+c9t80k/ewgQD/9jUOV2ZtEWjkfbf+4J+sqS++rTpdOD9hB6M3t
lYMMHzIeA3oodyr2Oq/reetktm3w88vTgkvFvI0FxjDLjm3IvcXLlyynDxgQlWaa06pJyccZnXR9
g4eAYiQZZAut/t0uPHoXCu43F7TMfJirFsgzDGQC7eQfS/GaAgql+4ym+Gjk202Nvgd1GKp+CKu2
5NopDJouYRmbryFqnzuhf1bLP62Hrgwe/vXbmgPeyM8ymlijGdIeQYvDySwhx35NxD41hvftq4dM
8xa8srysGFf96E3jrG2iM7TyfZNU56/sHIFnr2xUxsJ0rAVXvr9k0KovctxtTZsVkRsdqamDGwPL
RrrNJxGzwsYiVM71cH3QtOdxlgF+olLkDoFlOzZVdqXg6HSbEETjTe+NFfBCD/1C9tzb3YEHPDe3
Qjz3ZqBdk/S3iXnd0D2K4SJ9RjQW7YrpQPmqvbaQDJWYuvMopv9S4/s/dMmfjQ6xa+iTS962zUZq
7Zcwf9F3VgP5fgxj0l7sW8agiVhQ1dJm+nKD/3Hfra3BHAJTg3Rx524kwabQ5cERCT284xeI/VbQ
/CDTTzkict/CN5hXKWF00NrG9n6be7YdwV1gqEbmRdHR9QUYTYVqttjmKeMWqJU+XLwWoWn1O/Ih
cU8WXrRBqxMRgKiWY2hJQ1MZOUl3Ps7WaVuPDxJIvwIkqnw1EauZ1cdn6xg2GtHC9Xzt30s1ecW5
ta+J6OGhh/3Ead3e/WPsYfVGIZ/dUmYeWQaWPCYjlWpaa6xmifdDdgO43gaYL4s2W0mZXsHIfYO6
1Y5TYdl0pP940gYR3P7HMVlLC7ZxqqllQoCiejYTcP7cCcufVKry7EzQ0qXadXNXGdQJK0R/85Ey
9w73wWhjmbzRRGCwh4zjwYnkzwp4w+Q/m9h/CukQlyNCEo8+4WV1mFmbVlmZDGfRGKV653t0Suad
jfXAt7u+/59A7DS4Mz1DQqzo9XdyAXd/+PaXI0oWG8YW9FA1oxKYM+XZ8StC2NGaBSN4n3ac/UKT
0fWtGJd+YQjMRrad/ajJFjN9jhX8LbJiGplMb0Z+g3FPZGQRO+8BOZrFhCHasLpIKUmibOvXd4MH
0iisSVn2wm1ODaxRma2584lMN8NRclyymOy1xxnahn9lrxy0pPRk3OyiXASVzKQHpUPRBYZMo5ET
tFqntGAnqt34tuFPzXawSCgFIOBfSLNKrTSMt/GxuNIMwKnjW4fEnHvA2pcnjki/QI4EZjU2p9FQ
wu/jFEivVW3+NHTjgeybngeD0JO54FAgW59ZCZEPZxClCFRPsJIafcW6y43MCHrUiF74xUd8QlpG
vTNtacI/2od8wx8IqEKedfcLf6vvXJRVPf4sfefuZvi4LnMmZwuKkCrFjD/Mf9lHKIjvGS9d2R9R
N8P9T3kGPIFbSZR2uT4rZ4AZLGFcWSE+w6O1EPVji45+WuMomr9S4W7tQLyu6AUhIBr/hE7N9oHP
ePOupq2UKF+ScapIU4yDjXf2tHwJi2gG/lMr2gqN+h7n6n67zo14BMLgJTyBQ+b1m420Z9Bzj6Dz
OSm27X6amckc/iKGJTmWP/xKGyeHUd0gU0SbxUSoPHP0txna+jj5HNKkEbT0p5EA1O3ao0DQeN+O
3kCvz+DXONmM2/9lyvs1/6ytk85PG1yUDWG0+lgT42BOvz8xUb0orPeoovJWpT/3yDNVNVWeFwtp
PWgFmLO/LwxljMqz+fVWGVnkZbATEUzf7vniNTgQzNcxdTRmhYrmwueQABvEkxxRkv1doo+o70o7
WSr2/0hoUL4xJ3R+k4bZBpu+/NmZtqohy203vrdsqyluCdaxi9rQcQy9HQBb2/sjY1rzPtsgtoXl
48W64X/57OssjfCJMN1W4ic3UJ1yf3GUsIw/yI9yzw4bEXkaLCPprBItj4nnyBrMEVpvUhKRS8FW
1wNpEtsDCyCzzHwDVjt3BwmFbYvizEyglzxLQnWy1A0m2E3B4WgOzMVRSHacSfeYr3w5nd8OiSNN
dqAW2Avhfqmy1TzHw7zgnOhtUSthcVMa9bhadQ7XlkzvYm9yTdVjH4fLmdkedzwR0feUX8IUizjb
J6hRy2h4mV06Vbza+9b6JlAvmG3O4KLoJ/s3OUOlhm56EqX7kkqc0igXoSaCXaZnOy9dUEFtlFA1
d5O0uGc0FiIJGeMUN8Bl9YeLVNDNyl7otLA/R5gnKLvqhf4jEZjv8NAUOlZJL5u/C1bZAiitUb18
RjSdkAbcAVC+76b9VYRkER+HZ1uuaxvRr2gCVUXBRTq2sSlEDlr4Mz3x6qcL4wWuf4kZtJpeqS8Y
S0p2oVrbertdcuqFduKFBEwsrYNczsd32gZbYRwOHafcw1YMZz7EDB8rGrQUJZ8mHDFvNk3/LR5O
PAg3IesazYXN4TNPZ2w0qgf7NXu/n8KJM4yMEtAk2vQ0UEyvY0cWeU8y1SLI3UPnUAvlzCUyDJb7
SqPlY7IpBGQbK5YQCZFpac7k4nbF8I+hijAHxLTbt4o8YMgihJzgSAmmscK7GBW6HAWsYXPZBT+N
HhuANFE6TCvZqQWjaWCrU7a0JYofE7JfDWtC7ZxyRanziBL61bCHtdNEiUklajlm3hnnE7LJ+WUJ
BlypW8uSf//yW3+ZOe/3TmRBK4vT2uCnEWQBmG+I39Z59RFOVZpdYZT1fPhBZVyLvs9nklz74upn
p434yVhH5zDnAGdjt8Q8tsRzCCfFCS/l8PsIhmcje169JDgbGFtMKPFn8isMiXspnvXbw4J2oyaR
xSxrqg/WOOFtKgnatJfx8uSeniOdUlbOrYzzX9QIjRu4mDO3LnYF/L+2SCZy6qo2hp+9bTA/tudg
Ef9hMITsmU0wroZ22pYnZc32n8qAfO9ulUtGuRqJxot6s+86CLWrBnqAYFM9EO9gJIyRbloRaczt
fmAanW21FgTplBCNaSYOkvthY+6iUdTNoGBiGV9UM875eTd6KBi5V00g4DWENgLp3nOYi6HvUsIa
2KewZzKhg4MpNkgjC9HMiwYplH+lZDCegjvSGPBkhTOTnjIi+zxgcNdxjpJEMxIQL6LVYVnoMET/
dIAE2dd2k8v3sNKQQ71aC06uIr8jbS8KAZLrMXIU+ypwtoXBlSHOss3qPnY5RgwhRAK4xNiQNAq3
bVujfgczxBFywAlCn4YxC2K3gYvHvybButCUXQFg8SBATlsKY2rJWFIcpVeI3s0bRQWv+JbK8Y4y
I5ZI7GRAwpw6fKkh2zxeXUJcUcftacCHTp9kUi/zMzukJLQIiex1ejH4CqhjmUpSWweWraYd3vzC
DIT1E/FKwwVRkcvq3qR0V+AMkV/bbfuFU9PKli92nMqA1w7+C+IEC0ndq26KinBPWzWXcFkQZ74I
sUd9ZdqTtMjQzopFQ1QYqRloQxv2FlnEqKfu1QgUGsSoMYdCfF6NvCq0vhzhA8ClTfAil6lujAMg
Uwg1LDfZeVouDJ7yu48zidCpbbjvh+Yq8QiNZj7Qx5YZIAWsg9jF/vU/+CPY6KAMG87HsSYGiV7s
yENZx54pFVmTTqllXxd8bXzL/VughA3gab1j13K+zxhIxzBRMCXkaBLtqLYa9/s+oreLqYOe+BJu
Tc+jBMun0pPAHtu4r089Fax78+bFFOyIJRzJwiKowp9W6jFQ0F1a0/guKOZQga3/n/UDNKdvCZjj
SCxQ8WvX7/xgHsvid1nSDzEqoORlEW14w38g4x3r8B20+pAQ0chiO+J3Lhou2iZw+UhOWFJEh6NB
scSTQLToDTTdEABIvhxcisvsDIUwjhjWPSrvwlwzprIpSUuQrGI1A+ZPhliStvfS00CdyJZgEX2l
Vwg5HvzvAz+G+HmMoyqoIvpXjncV2MyDYTa1kecXDWVe7wybJlOzDfDI0eDM0n3UD0yV1U+HoanB
TKDz2xJX+MScK22KRYXSNBuzetsCpoaxeb/qw0p5i3K1XBCwSJ5eoHLUlD9tyGnJL5yivtfZBZVb
jooGqbrZ7TiYZBmvUxGINcoOjIYAR7hKq5f21DJ/uT8xVbXU7KMhggKSCyrzKzJ4XpNsIJzkPEdM
tM3cTIygJIqX7aUkj18ktyKLbelVZLNecjodOLPDJ7qsR89wHouEUVelJovGrtv5phbZXOervn1l
yz02lXKc2wpjt93oGsN6igxBcL3ELu7NqAq1EusC5UHzm77sqWxI0GwcbsSCIog8dzRFE1OReWdC
WTc8jT9rfY2xIihCpdaoJ8N90wEfYJAy4NaufAsDoMrCdCKzj99klLlwhHgnW4qy9MPglgOdG+hx
ZoyB74W8oSSpigMRMttizu6RlmH8kjhyZJu079FCw/gdFU8Mk7Aze538ZCY6pKXHaubY6hP1DSMj
H7L3L9cO/4GmTaRY7STNKsuTR57tWfTER432SJ1ib2Lilkf/a6Yr6Wn1ATdEfEJLdSFX5j078N0A
1rQEdlCrrPbfwbZ/yh9n2tGOrqSdXuT455udoIUjUCnIhiFwJDp6uJyGW8oeG96l1/QFpOn7Spt8
mqBZbqnawi0fovVaG6o+WVqBbp5BsFV9f7VYe3bIHKQClfurzTvp5NxJ/Y1M9E3H6bi1RCIoMM4P
PR+9IwbZLLWp9ocplssE269a4oB4pyuZhi5uXwc/hWFg24r7vdJeAiaxyzkv3E04V/GUgIf0J21E
18MMrfpRmiJgpyby4ltyzUVvTRW/msJLpQRKZNeUizeQolV8LJhTD8fdP1ZZEefI9HF+o4rv1ulM
HGxGbCThtF+d4ktBAJ0xrseVjkODx4L/SWa/17PF88vRq6Dwy/Y12Btpm4FP6Xp9hj0mHeJYJW6j
hUjXX+flE1Mh9+kSkr0YYE0ov9xpz9yCsg3bbHr8t0yMJWdRyn6eJafVEvKHSQjC0EcokbTysu1n
bKixa6PW2XuZYLb1nH2SS7msy3SVkxbbfx17evvuq8JCaeeKIivEJG+uHMPFAMggG1ODdgSDoFi4
GcEnBa2CLItadRE5e8971qX8Gg3zjfzDTTrC6G5/24o4JVsqCtoCK2frjd0YwNlkKjWF/qqN2+gq
NjnhPoGvbq7j8O6V0WHDMwQ0VgaVsYGsq5PplL4Sc4+93y4e5d0xgq0jGLvcj8ZXmSi9NgcZPOEB
7ruO781pxCpwXlNjzhjteDa6mQJWQP5sh0ox9RKJyvZoBHB4z/4UU3MzCspu3iXBDnch6dfHAaJ6
QYJYhlDxWXk5KfWU9xmkhu1HescX/J7CpK+z1l4o8wcMfSa/J50JL+iKBVbT3Mm/96OAurctXcme
QC7DxVGzhGhaqI+Lo7l3VGDWb+GznOZXBKyNf2GrfynGzdrEs8D8lERfnnc25WMdOZo8zc4HMjVZ
GpGUGdwZvRFMq0MMnNQWTGxojwgfNuDRtIMh7JpoOO33BltwOyDFc8vY26aY/0ux84IS17WNTIDW
fMuzYmyVijkrpPrwfxgGClpombSRjVJlJo8Z/hFNZmnnpYiK83eX661kXC+Nf5Ne6UPrdlQiZ+nP
jTWToa9yVSicx4wuKgrFPjOFkmlmDhGY93cvr9Ec2c9Rlf7dnTzmYB8F8OVb4CRhF211zh/LJLBv
UYr3ImqLbPKQW602L81H/GIIUUHYRcZ1XMpkb21vWUgOCpIHqLV/RtzvCbvcNfwdWCqKjw9G21k6
8blwTrWWZxbzNIzyTdumk1l4VUvH7JY+SNFg+WfcMSN8DUrrzRDRrnN2ql5EnJmnd9fI+l3lzUZK
uQOWDZUaJ0WTz1RaKGvGkrRWxrEbqoPFzXRY8saKqJjtWHldQgD7t1gmPd/4hkbkXddvbycvAMtm
KFfUzrEcTxO+lN+8RtB/fIq0sz3UXS2A8HmTAR7RdnF3V7Uiq+0ntoOVnkVveZmdR8irkq4TJiYD
HfykRP1hv4kXOQ0haGOgPFKzjesy76OLoxsVqMBBz9PUz737CkXKP8IZ5FPh8RLkhLRbOZJoVYjF
9dZml+jkg+jxRdRMPVSzNHx8SCdFMekKxCckbdZMDM0xtP/WefNAh4ewVolG0z5Jg6Ea5iUKW8CB
3gLT9dMy4w3x+KFoI5Xt0wm8lE5rLqmJ9+19o5iWHwbCOmoLdJBYqLNN6h5hLNU7l9PfcSLkAcCV
bjK6GIJ2XLyGC2AFrVAxfsU9m9eFpgNsVmivFqFDLo7vZXtS7lVMMP5ia6IwN0otPlQ29k66igVp
KafVioi+ze9Qku8Z1c7dO4umC4w6jw3AfFOU9coZVIY2dnv0jF8aRaLydve3JyHD3lTLKqStpgae
aOyM8rpHaLbPcfBAfpP1u/Esfo0rqd3lO9PWapINS/6ZVvsQuHkx1z70fGPR7QmuNw686X9GGx9E
Aklt5QQsWXS6yXMCqoluP3hJuqQU1OmXT6UKQLg+t5Rjbm3ZczCc3lq3V8go5OhcJZ/8SOVGuQwa
A5zAmRG+h2aoTESxRBMrZkf5q2aRzQmb3Cay1lMEbCldFQbMOJRPbhouicL6PlNFRCYcH2zn/Ayk
eP9itX2/3aPXfwOBOQ6E2A0F+ftRnd4f16ZpAcZs25zql6zTPIm6P1TXN65r2P7W5sSfv7xMK+5C
OiBf/jNKu/x9iYzzCPRjRFywLBHAmfq8IqbICoG4FmbCF3RTIZ2pkgoBHHcX+oSb2sN8OafiNiOq
656pz0OKwNtVk6tvIeFwrK/ATtqyTruuEpd+ztjLK6aAJpr7kuUSE7DWLonDQOaPygRTS2X3R17f
B/D/SAl/3zBFQdhtFvr5NBhxHhz7ETpX9c15H6wJh0GusEExARDUXHfRprPW+przp6suLB0qEdbf
DB8x/tzYCy99NcYh5+uu/OGNh1qtm+X9uogZhw9pgm2Z/Za/Uaxc8UgmkMTCfNW3RsCM3gJG4wie
fKPwIckGEkriac94qb+CWfVGUTe09dhmOAL6RmkHdjqBWVUEujxJgm1ngh8xZkhWLw799/oVB0Dq
JG8GC3dSvRDd6XyTB9wwMw5bjgx64TJq4T7bEzDjaZqWukvZvlpZd8acvwDGdFtps4LgjQ7xl+GP
G+XaETIIHhqW8d3jkDimQkc7wGUV+nnCH0ChmxKb5ktDH27FSRLS+w0001ztVmdrasqNO8OB1Hzu
vJqna5mdXeWvFXNfosZD/6xDBv0ASrxr+doiP2PoEehmzAG/u6B/ZtvnAL37OO/pSvI7KW3wSjlq
o0By3KhFO+1/t1H8PijGJLYlalYW4FqAXcMpq36/liISOG6b2sR8xQ9PU7p1qLTAgv+buZVPafD+
w2YFs1skwS4xzfGopkEkF8Cq8fS1yUtYlCD9WX0WKKYSnuaSlbtvfNGZgSKC16+zdoYbO7RYJeJq
LZHhxrOnfw5R4VW0NLQ3b9TcK1jx/bt6qbXg/NdStWvPD21PCN108iqKbRFO4aZQZRY4tWIUU0Dc
3k47dcZB9LZYOWxtE9YNTHsK57bd6tRtCHAESnZhBu+Cy+xqpD3eKzRObU+p623C0+ikFrgS87RM
FwSGcRz2g+RMAmSJCw0fBGGIb7dGR2o8ggzz6J4F8cYzSR/wZDVn7NxAUt8kFIubzSd9DndRo/qO
WzTMmRS21E/swcs4WCIaGHx3uzfds2Z4N3LqwqZHR788ARKyw9gDd2qV+bTRR6zTGkjmagJDC142
r7WDl2UdY1i+yqPSFvHL9NzARMR1WJ33Hw1kJEtehpv0H6dwxvjMsAxJSdqKX2/pM16yCEZtbKxg
U75J4/vVfXxT1jApDNZSOlhBGjoKkGsCTAiUfgqWNMQVVURplEy6KY+YqZWXTG3DdPsz19UgNabx
Z84th8mX8tHUc5KNRZBlMQTHlarcLy+H6gZjfs43gL2XE0YX1dG4GFIUCC3GnSmBn1053MXsdtim
goc3NObo2NhYTxfWKiz5zhcxXwRe90CX4LnPFuAwQdXNvbePcvjXadKLA8XZ6KrfA6I0dN9zNEyy
QAExSDPoMAgbQm5VpPXTT2I4g1n/2Z+9xIOsHR/jtgcAW2O1EgSAFFQKWav86G/dKMuICBMtfX5m
+L5jOLt3ALcAqcJaOTeojudok9ynd36kCK5uzyM6SJ4K8NEOl3BE2+2V1DshCcnxAHeOKeq0Z8nY
UoKJwC4IIvogSGjwNNxDCQC9FtFXJHzqvd+PEL+OjT2X7dT38193sRnkmi4uLmDR0XwL0atLbuL8
V3xFRNom7Z17DKC3sApXW8Ez4npV/g/KCX1bNj8fd5Fo7XifVe3kTd2C35Tbjx2+nvYOFvrE+I2Q
cDunpVj0hdDQNh44AVf2IMh5ou+exN0ilOKd02IhSXY1lTe+vR8apHK+S7w37X/vnlPJ//bPD5tl
WetiXMSEidkCbN5hWNtIhhW0uFEK/cXk83xsiAqFnIJ5keuufW7rC+Wqrwbimj5BPBj5nqF++Gu0
lvRNc32/TkLsA+ziU6AYxwc9VRwfjel6lz36+MmbbKuBHAxtd9Xom0PNYspkbL6nwSmD+QEOFywG
k3GZAbhtHu5ua0bCeuo7H+qSRK6p3PrbKHuNEA6O7QZ4dM7aD58h5+V+gmpRK3WkMU0wIGHX20VA
/1SxKW33GDxvPFEjDgKgHucnlo5Wrc/B+Q+A5viGFglDp49NkEeycr0eJa1jiwf3XuvMC4pHZWRn
QUwpNAZUQF4BVBNQJYmXOzDQiqy29WLdYBwrTi/nT0OOHgnHpXXVOwthIHlMm7gJWXlL/sMl86z3
nlntbYHY+o7JFuTHwtiUT3flp4B+DPWX0/dNtWu9sH7NDsH6bd+2yF+qKlYIeL+0NrpSc3G4CKvA
uiAiuyk5fc0NYPQx1YJhgmheNkI6kvjss+VzB9aiQpzQ2UYkHxTwd7lX8EeI/Yf2NlSNZCP0XErk
ZOWcO3RWvWYWfLr+BAt8oj0Dca0rWLmx+5RLl2A6GsH+VPdGPOEig/+pdW7CgG7mQKG+viYQhYwl
Yxupkhsh6HRgilxTs55PasMqYr1TTH9UU13uHa5RQfyRbCKbudA2vzDarVpU+po1lAxcai4DwdmW
NH+v+fSY6gHYm7vyQvDH93WbZUR5ZdQN/Q2ACObJMQPiZkGRYHw+YvvICvB7BdJHEQ1a3hEmKWOv
ucwk2AUFu08OVk16gzkvwLoGNahdHGNOfrbBpCv2zNNwyYZkTuPvuwvFzI2xddVq5rXPzzYT0Two
An89xbEh1hcEOUK22HqnlDlBJSHmgJrpU19tr++E4AtmSw/4QwCn9LieGB5E5Y+uSVXKBNT6YwI/
+IJGkLrw8pivC1fCsGwiGLl4clPJqhfmU00EGOuFRYBRsuGVnb5tn9Z7y5954a5h7quEQy6YOuEw
GAYZHHuOGe9mZT8mYgoL17rxsSIMh1AeIHcCc0YvRHUK/0L0M2YIQ0c3AJkX5NdMYRoZWlzMKxc0
/WoNEa4w83jeKfrYzg4lXmukYblj1YY9ub7FZoB1iiM5t7fNXj3TD8E+CEV6twm79NWFVxo6N0OO
v9EHgAJQ9DXniJkWpnDYb6xqVzzHuNOQNL+V5Lm5wEu/2ip2/wiXVdD7+ZW5Ged2NKWGyhWCfrjX
lM3HeBEwrB5yWfNxk6+tglgIUrUJvnbUVjuKNYqoC7hyokHO+YbsMCvbY05Sc0hSBI2MGLl5K3Mf
VsUwFbQYrQqC/lQyfmcXJCDBxRPIVSrYYL4W1ncX2iwJ2xrbl1j1vbwd9q+KWRhnXX5NXN3mAmdK
/+FxAnMIY5qzxCWgsJInwKXBRAh4jGLI7m0diMyR9SZQipT0KYlaMBxmrheU87znLn7VCBoXI0GU
Ykzh5vTN6ezox5hyzYlqDz0ySivXViQu0h+7Oq/lEcYqK8A7ZzbP08wiWr0WxJ5Cl2Rjx5xWeZgM
rxmuKdnvJjHqdvG2Q7UqXP6qSX6fxcGcvl7YiG6KS8/7IXnQLfG6Ig2oEZBKL4K/F6MHh91YneFm
PhwwozPMoZ3JZyXv9g7zEbooH7GDFlFYY3f4LiuvQrsrBAIrWOznKnqS9CU9iCGODWzcT5utpH6s
3M93tVK3v8vsDCoUKWDntDi6VsTT+vffW3b5NwKcWFDgzOT6c/lM3HSB26bnjEATo1MjEMWEu/9c
EaYfOrPfHncBydP0LUWjme2seCn6C8ojc56lqLS/q+wwd6/ZCdvDnfImPU/sjdBMuANCscNIDEvc
u7ZAcEnnwE2l7/LRCzApP1Lw8qeToewHSCmSboMUjDzf6K/nH74Oq54nHz/oLseoMw88i3/Q+kmW
KXzrmDJ7SrO5A6d/Eoq75tLbRCudH3KkwxqHavdvL4BsJa4RjPmqr0jhZ04pH6MMoElnj9Y15W4T
0x01ZwylULEM9VYR17ltM5iAk4IQLT0DoZ0rsJeAUOG+++iyuQpT6GrC4FRp1Yi8nldbnZTgIA7Z
zdKIsGUOYLsY/9mRd/D9kiE8TtKDmpzUwzP6u3kbiNNfuHWWEz9h3HBwClFfP6DhyJLNihEbkTVX
6Ns69lUaomguP8e3arSA2Pj9jeSltlfv6+Vt2LIiD/8bSwATzfbeRjKB5nqBYmH3Kluzrt9MHyoW
JCrOeP5Yrcyu22daiSnuBxUrLmXeSHck8zaGbwEf1UC6vW0n54WUm3VRGi3BYL9PACei4S1vbkam
azqa7yyqTWp2GtxzpgnBxqtExGbAceAGFC1G9JEMxi/TuAsn0O8NwdtZ6o+V5t538ROREBa/OIdW
ghGocQmiZh082mjPDf2EWs7yXvDH3BfYMKzrGJDu1a0XkMuNMBbHRBLxJcpz0FqTMINwwiLsDw+x
eIoFxXPSPOUbhBFv50YkOBOBVrKHgGM0j7lC0514HWdcWYwJfUiNB1xFONKJLZz+dqzrNb26k/am
Y07FNp4HJewXDvfN1Xdk+g7jjHAD4mmmHMs4ruWel6RsQHuZrJ7Oddr9By7DGavfIRHhKwS/zWjl
VE+WXGeYu9B1qT+es9s6VKA9udA8kGEHGGYYOo0UKgY8PTy1ZLbYd/4GtoIT0C6gDHynYiHk+eG9
LXXnJqtAutp2h1kHmtnVjSdFSuD7XRW7yFyLzUMjNxVA6ljdxA/CBBxuUEHSX7XnqUcqVmqkhok2
XgfGgHspY//V96Qsh713zv5aw1LcmqHFzt68wty11jK0Y3cosGrPozCbx5xRh/Vzh9cilnGDXvgP
FaUxTmtiXf2aCklFZMJm6BvWWOOgwBVgMYZ2IZHRXLTawaoKfXjUhjeHxJDzb7Escd/nHjbdSLAf
Hs3tOg8wGHhT/d2p12xb70ZLuQpOefPVQxyTTJq6hQ8qTRhsu32u/b5Z+URpED0JEDOwpLvcxMCT
/fsCtwnVZzdQTkdd/qJbZ3NmTa0arvqAVpRAvb52+ARmzvYpgS+DLvWR7TlfTlMNa5aeNIcsoevK
o3OQbap5n8pSBmSUcoPUiS93l1h7iScp+ikpkjp+apt0JS6fv+YMjteqtaqT9rjCZ8c532o6xPMF
NRDvx4ep9+gJYRNZXTlaP/ZNaKkXYH02xUmr1dvlIaFdahC1V8pqUmvWlMJ5+VTpd0+3nlwmbZWL
BCPNYuSh1pwwxUI3bBdOjq7HYlBAK3qhLxM1yJIamVdNH9UjXqu2hvYjKI21KlZ9mPT/yIgJJRqh
OT68E5Z4g9+xyDK2ChXs4EINJXoOvUo1On7u1rAnLkNa+hm5uJrAGMb5K5CXGumHj3HJYA2MzeLt
xB175hsuRDHXIhwmJrH6YoUJwsMaMEbLprQ/aTa/YOK2i+hIlbH9pX6a2jbIwbLDfnHSBIf42MQx
YSFt5THi8vf4U45ySwLs6OHWfGUzGcAQolRTIp0LuKpkLJFxpGfrArBI1veqlbO4CHEE8IyUK34O
hhkZqczT/7CSyTfWIzbsLZU42Q0QVUr7BixOThCm6J2ZyaWmq6KGDSKl9a5GOOou1x7wKfbv8Nwr
bn5ivtElyz7iNxDpdCeJd/CPRxsHuHrDwf4J9LdrOcoNGsDzbw2mGK1feNjvt2uQFTLGxLncIrRk
R1TzkZ4oc0j3pd0DpmGuamhojx200KMLxRwkx4KwLB/fe5r7QgDirVbm1YKCrytOEEg267a+d7dX
0U+JM3rXgJVfb6XCQevVrvEt7Ab9GnG05zcI+HpikBYMT7GAb/OiFixouox1B9lb9U6j0KcWDa49
22Uvy7RRD3Hjb41Ue1HnmkYRu4qr9+cjyBkQT9iRlK/XkKC0WcC+4/MmCVW7bO6MzomFNLDMm7QF
zJQUm/eBn93tvTLaYyeiHjqlmjqrwCtWBdFV4aDeQeo/U8mKPiE9tNn9Rmt5uS4C0lDMH70Oxe8n
cRicryoQZ0p5NNVN3ldGYDovnQxql0A7VXL4De6w+uqejEPxaXgSFnjUFvxt4H+ir5O5d+45akMs
6fRZzv6XvEdOEVh9nRPToakxeV2hT2KYsZipD6lX3/dpIw0Q7Q7oGkqzQJwQKZXUIONpNasNLNNr
0w3S560FQuFQ6tcUAY+QblxZmRrZYTChmmszW2b0nRcmGiCejDlOVo5y0OdHBHRjUXjQgIMoccJ9
UasruDu2q+D1Ct4lLAF5nBClPS/uFHxb1tr6wjypaqyrafUtK4bu49YEkGOhuGiqkuOyskJlp2FU
OuUIMqBhIzzNl+lZi1lAx90GyHjrDEf+eZXPJU7xSB7B0BUKIX1vl35W12zyfIfrGq8au9sjLjm7
aMRnl1h/H5Q6WDJwedIwyjU1pNaTJNQNvIALXBoCgDerl+/FocCWx9Hm88poa0WuZo0As68js11b
XfnzrNY4nyjxEg5Mbj3EL4yqmpa5oDQc2tWDEOt3c/VsSv6VnRiOTy9Tqrc0MiLGo4x8DpSLis2n
NXfb5YqPgBBgPqlNrbJC32BnT3JYOYP+0gWcDmi+TNR4FIfzak4PzMPtzwvtuuu37n3iC4tY9moi
dlxVLZ5ZkkPvd2eLkst6qNwP+YQ4LLlIDP9G4CNXwsqYuy8MHtbrH7hRjDut67l0tpyPbNROWuRX
y7+DaxotJbkIG9ZK9UnKBtOqIpY6qgJvZ40P+NiAzy0yb3vPinLZfqgb12W+4K+gGJawuaqd8/B0
EXoSUO70uqeqeYbS3mpQGEzDMacJ+wX8sloP8TTxt562jSFt3nvsOoL4EeYMxVn3Dogs67ZFPThg
+VHLPSxL8F02CbhQ4L9uefABX1RyYt4TgIAfqdmOLBfOxwHF27S4rqN/tqOJAAUaHmL0BzTGiogY
jkiNsa8EKn6gIyl1aqb2NULikhikrceJmtp5fvDLAkfSg6Isz8q6h2kcpoc2oPZuUt07di1ZUpK5
eRV0g2YRgOCyKQkQfp+EOYRiTSbry7oWJ0rSqT6g03E3piqSTAkzDrLEvYiRFSd+DJ/PQva0rbBp
WHD4T71fUVOXBSeM4GeD7omJhSpsCtJjdHlSO8iVgGLtwvVgl02etR3XlVwtzV9Nhx+St5bRzJGr
w3MPej3OxmGcuamhSciw6piLwv3El0TO8AtXbmi/5rorE/xVddQsdVIXxBOUhkCd/9Ml5mFb/Hrq
F+VUiYaRaHrUgqgbi39L0HkTMOzOtAlQi4GWpY34HkzMGTIEg2zznYqRULDtuDGKeP5xS5oweZJI
q6BNlTDgqfbtf3MQW5jV1dS6FgpkkammjiN+4oBqsxIVicZGpWVTJhVZfEF4jK41yAwrVWRHNjwx
gOW1AkRH2rAKTSSzILhFpxH++CMvcBzZAiZbY29EWYgJFs6VQ+HKpMqyzy4cGNPdrHJF9z3q4LgM
kWMzbA38vpky4T8hkPqyYKZbBlNhPdmPb+6R7gLqeWylsyBbaZWC8K6HDpjFEtFXKio9zb7NMvmj
6iauB6KHMhvLEN6TzOk6auIJMgf+lFdP5QfPWczQvVhKZhay71e/vRus7UYzMf4V5NEEL4tx+gAo
8XjX/5FrA/XQaA0csw/u/aHNwv9pJgnhRgQfK9yR0ufv1SKu1ZoDa6C/fdXHcjIhyQu/iG2myAhT
VINQhL8vKO/f/j/iv7Ttsg3kWFslmWgYTabAZnzeX5pmVVzGhg0wf1I3aotD7DQv+QuCuTIn1gAH
gvTUF4MsE7CV4Ph+ZCv/nmE18mCPaswoJ+umxnCMcNp+X30APhq2Cs9lOuEvn+6HbVcE19kOb4z9
kHTSthOKLFh3w3V3iqAjhtIS92cfxX4Ush6HkIEz9LvhIF+ZJf6+Go2D84s9xwHc2HKaittfpOTc
z/u5n+1+qPpoNv3m6yMLZ8XGUDW/bl2MAfoykQg1NSyg9co4qyJKsTYodhmaueTTKcbs4xviSYyR
HfYnFjVH2qEn5Ltb5MfU3An3q4xYT5VI0Bh/snNiB0MIGjqMNYcZ2pTA2IwQe8tzTFUYnAsBWqlq
yqGRvgQg7YbptOWmN8nEJPjeB/BpuBOVb1Y+ojHReta9EyuX5sFSchuexd3TCvWemvm5LNpugfiH
QVJ61ijr/4/OBERGzNwhl3fmTEeE6fYsNDP59qXH0M+oz0GDDcQ4HTmTaEsUISmm7JRdE90RBFBt
t7vzj44W1odc8IjmkfMH38Uk+a1HbzxKefRwDsDvfwwmmDqKe1YoqPwaZjFDdnfLP+I+ENOZ7rZH
by0FVHCHp7Sgc3hizomyv+5PuSkejCXlntin22sSWJrJiPuxs8h9g4znEdLd1PfmKYOMdtQxy3+Z
aeZKzMt3lCC7GW6tqVUGa2lo/z2enF/gzgidW6kt4NRVUhDT8/MfB5bhaAaqs1IhS4hd5t9L/HnL
0R6WlALCsoadvqwdvgBESKyL+1i0e47rN8Nlgzc9T/gmc8jY/6L7C2rpqFmEEf/RkiUvNcDUZIBw
JU9pqiKDDks6SxZuG6gapelBRiWmsMzyHvBpupj1WXm1PKp0kHRDKo+H05SD4QVGWd+664h8SaZa
Bn/fiEYJDQsmtMp9a87poRcBGy7tFYwBPKdPNTK0/KXf6oCQsCUyP/N58hTW8btsksc9SOqo/mpe
5MVNWRm3sceFOKHCQ9MT0YAYlLmnWJR6Qx5wyWEqkYIzV62mcZl3ZdjFxTFOo2Ag+2yTvmy6/7IF
97p0fmegzD8Ax9Hj69KhbkG3mlzqF/rHKA6dFfNyIOzP6ciYOxri3Pp6ksSBI6Ohl4SEGUN0yPoD
wEzmHPxOSDa8xsPAoqlBLk7Ca5MoGNvMwfL7fYV+z9nNaTvWf/Z1BD+qpRkkWJRWbI+5uGMdBbLS
HmtRA7MZXVKIepfn98FSTz0jQ+Wc1TqByijnlMgbJgZ+wH8MFZEsPKAbMxuD5KeyO0ryHGW1aKTL
eHWvpsj3Z9x74DpeQvRwBBSNGVexCPYOC+2f3aAc3sKbThRYL8BFaJpFDKHcWOEz41MEH8oUGLgI
UZgqfSdgTh3WVufYQE3nucxkJJN3JV07ggBq8FkhvWZrSs6EoUk+5ZLBAjjVs3dJCWmj1ZV4BWlc
tyFCXoyzg+UHUqIL7X7T1FHEPEdr5duEmhjpDnY1dYW9pROhkkg6G/XGSgkK8Y3Xnu0K/GqqcefK
bhIaLXXOOYjwruO/KcLx0EheekU7Uiuh8f0cK5aaAec0vA8huGLCCS92EtZPVs+SCZmN2I6dl+GA
hxfJJJaHJIsD1gM6OJNj1Y0x2M9fzBqYX2Q4+lPMO8QQjONDwuLf9zS8lzKevSXxAZxx3NuYQ+BT
jpgKMeS2euUkp6C2jSgWqkUm2PJ4eNEsViNRA15I5o9knknEA20LAJx7PS4QSAVdQ1tLTlDpPiKo
9zGFBfkVHhuvXzLoAqS09F43Xqf5WPvWBO5kIUetuNwSoQVeC8RUaMyHIPpF60KEGM+Zm668UBls
O47rgkOv9+4ZIlQA7dtkbV6vrNefo1BEvGFh0FljNr50K7CnQfA49x3J0+E7HBy7mBFmZydHGmiu
va4dIK5QuO4F7SUdzh75j9bLA7fqbjDTjE8+Dx8cb6xITWeUA3LCZw/tarGJxH39QCBhSC1l7wrl
1o50oD1bAbh7uObWfV6YPQ5oQDfC0HzFkhWwD82BBfRUUQPaXEo+WgyebbkIFF0w3i95XVSSMh4+
pOObroOL5FS0Dt+92Oess6/nU7EEJx7fjC/1l8asSteUOL3vg8XXPRFgulRus2rg+E7ZOzUlOH7U
Q1leHtFKNEneeWXAavHFxg7MOY/dFXl9SxH/9Z9dDCWaArOo5DH+By8cHfEBnURhwRP4a2KJjNmZ
yGq3iHwYKUE/FrVVGEKbcdJpLHen86JYxKBQdGkEyUMZ76OAmEilwKhb6Vnb4xey5o4KPP8VkQ2g
NSuEM71x81g11peZh84Pt/H3gVVXcDRQOE/bIqwplG2H+3wg6iKAql7Kwt0/2TX8dBxEC2d1Zn9f
4d89zAF+PTt+JvM5zmplo/a5x5Uv383iSS1awReDBrjSiFAhZrJ0DOTxt3AtfRmhe8klVUJuZhDa
IRcffJfgon7XTqKWAsTunKrFxORW8ACF2r0s5flPMHQmHNm02QGsYRCYwObxHbYyl06PNA8hVh9E
p/BwlgJ2FQvww18Vaj0I/E1MTLEG/NdKHTbJiBlVLwW1UsWq4Q3gk7w6Yy4tj3bMkj5s6IsE2V7K
GfpB5CPGPRXw4GMxuQHBskbgI/rvPS7VX7EalZA5qgxrrxKSgxSLPvn/oUV4pfGiaubA0geCNA2T
o1rplQw79qQok56+QjQsR7OvuIqEZFhF85nVTzyUmJr0J5rvaRImk9xghhN0xlnDIvJa9AfhuoKK
+0j0TJHkOMVdDvdAXtqFn71W/eIqQpHBeYHWY3uD6ncSvgg1RDKAzxxdWjlBvXOWsRVNIeKxyIF4
ndrf0Y5co40n3lS+svRQfilrP8/uZmNpmzYhVT1D8WOGA4ppAPiNj1qN7Ft4R8TNTQQ8XSTwaN9s
ZGb7LcMDB2zKURvfsgTp+78xHhk9RyRtN7uUyFqkiXakufZ1slas6ljlgjyjbRrQP6DMfmCJlnue
L8QrJ/qjJkuJzxIpXkEQoeFVb2ecfSCaVIiqrMryREYEP3a25ZV6MryF9Vknt5006wY5s0xlcYFl
eDCiDRsSU6Hgism5Rxs+iJbkHKNJPVCQdd4C1L9b45lHoLX9bxkDAqMrWUJdDL/tveEJAdg10VNg
OYWAtyF7uXsxaXTKMaJq1avreMrcyjyupJrKTVbTkgNsCpYuH40NxMo/rkIMCfZOYoN/itC3n5SI
CLqo9TAFSeXIyklz+plL7/XX7B8WsMG7MQxK+CkGZrzT+B/iDsmk9Cd9O6MScqHuepx9bMLmHKJz
PrxTTvIRs6l3L594KKhhw6zGV2VWl7/wjza6BMnWe4G3DIoe+c0eq2kDgFcIbsU3zSDcIuIbl9j5
BBCuu6pigKPEzJs4/fvopDSiknHMCFSXv7kF+Atd2vR4c6dImvuZOEPokMGMoNpVzGVKqcYOILDJ
INiFefSbgy/2AhEevJ/VIR0kcU+OAaN1HrBDVJMoXlUV/wvrDd/lkoz6ghIHh/7k6krH1NrSSWTV
wrRtc0yWaD5g+1qgbLWsfzJ5vtBKC4ueg3dqPN8lzv4KdX9CNg+E9IFL8GmLH5rOEoKaA7vph3sY
6hqRBEBoh+POnB1PT3aRp0wxxq5nuNGZq0oz6cHXu7j3tGSfk8tWt0sXwjpvThIJJMM20A7Cb+fO
qWObUaSKPO55kI43UoIh2dDjZCqa8qGCaGQfyLZMqhAzZzYRXF3GwwbDfAeot5y6Fad5GykA7vPH
jWk4fRQJigw2FNaOPPrSGTZmJepX01kwqhDQAHFYeDvOUK0ZoIX+ooWU1NABWwZonNRBDJtj1opw
I2ty0i4rnRpCUFGaSnUhNFXPYeYUUsGhLtp5MsUh8Y5V/oHk77oIqx6URu2l6g5+wykT0h43h0o6
fUq4Ll+VcrycTNDa+ZyEbUfHSAWWlgnoRW338wmht4MInkNOFG8cAY4FP28vjWpEWSK8Y1vexBAt
xBCeyiofl/zKD79PPwsH/BqypxEa86Lbt2+n91mWLBN7GJCYTaN9o0NZNVyDFLF1kuNMPfwEefVv
fFQojmW3F9Gm94WCrqkgMAuYNI9HIQGYf7MYke+PE55aJxIc3oIX465RBTPSveivxh20VbFY4BgY
UifSagshO+RJiOh22B7dibKaxFs3DMRSTOcyrUi9vYMk36XJQaRwqz7cmc/lCH97P3Wxn3JwxYAs
UvR/PAZPUktqaosPK6/3htCdXT4gHUEnS6x4DLLLMgeiw8eWJGQJDgMVEj3OCUnDzVw0/ad3yZ/D
UcvMOkSCp0VF8eiQWqztzabDqXplah70VXJrF5w3pqCLiufYfeDOmsn/4NPAAojbDwjJSz3Ffqxe
ZiGja+EBk1Y7b4EZiwspiRK3Dm3stQo3S8+6SyyMbRxsxfCO3J56Onv0vP+jqFoyu5FK596efyKd
PUFQ/3QhH1l90pcR1EucoJ65WiZybyR/eyf1EIZiJQ6zCjSXH5uH3Q7vAPaC9zP4R5TOJuhFvL6K
YJOut+epFDQRIBoZASTNswQXzIBCtIdj3+ohIsS/ST4upfQmB9R8AdZOBlvE5n0MZ0m/yqPfieW1
hTkII4NqFBkgx/epQLiZnS6PPYtlFjF6zFZnR4yLw6M2BLkLnVT63eFDeoARR0OwoBJHYJxPtNQx
kq9Ra06vSQNiGWcsZvUoVSzHtmTbJvm8qMlIsdei6qF8tWgVYfrMAlBXiD7HMbJGJ2keEWGTlJMB
WUW+ycgLIw4gs5znZlwnuFHAHbvLammqi+mqwYO2QMdDSsxawxuEO2k2ctIeRfk7eueGW8knusN+
qHGf0cgmmMRjRNJA7NnFE/aerWK1nIJ8/zMFYJnAJD/wX1MfszGB0k4FGqb9K3JW8MV+/qmnnhDg
Z+iBHK3DEOagcrdqgVTPS4AMYTZTQbCPL4OUgn69aCJjfPssn1Bkglx6L0GadGsHcFbW84z6W9Zi
OMnrk992BLv8BlZM8fnYXl+gcow/H4HDq2fp2OrdKO3gCKUtEKiVNAahGmqH0xhqkay88j3yIBg6
Elizi/6sFc9dJU5plugA6ae8tnbyNufcQHwSn9yZloQga4n0yCWufesafXjDptGTwHlmqp+jQT7u
8jt+/iQIqbFLGm+4xnyJr8ufQfSQoby7Ez+9BV5L0MRM5A5wC9PMGyg3dk5pZyid52Odne9prqdn
Lvw8ilnSaV6eNMro5iRmazYgSxdNuUpO+9/mnmddPz9na0y8Y/tmf4YkWzn11RR6PK8iDMR5zwlG
DMpXBw/kwKp1cJ+SiFJDVwYEHIkDNt2ZJJIiztxHxuJIhB6b+TwxitKwJfu7H7e9yv2FnRN9KM3h
JvAXT5ncrDDcSafqGATi3WH9gsb0LILrHuexYalOcCN2C/LB0NtI1YJqv3mU5edJ4RNcg9z4EpU5
o0RrxQtWhp5MYpux57XtPGV37nEv+gSM3+Bmh6JCHB0mLP2d6jAqu7Lnm83V8ZSDBA3mfOGp1yy9
O0LRYGYBTFcGfGUX0U6WAECiZcWbroOPDrZelnOt2PjiHa/7Sa3RT/4TU8o9aJQnKMKGyP669aZ2
GWUF0lx10Z7qF7JG+/PQZ1yazuEEKt2ZRVM+OPFvx4NYEdPH3jFEHct2rW6FAyht6gYSKuIuv6Eu
P1I9t/K8E2gouJUKOu1ZUQi9VSFoSSRnN0wWKJQYVBrFJ+Rj4NaF0hYgIbUQ7kv5zhtn7Nkghruq
2aglrOluvgTzc4nedkEExs6wZWLuATGAhtw+OAD7s0bJFpoTH8v5oif3MMsFqYG3tMNNmQYOOC5q
R25MDQQkK00V6jzeFazRBMs4h39p6WzCGJkaGjC0or57J0V7FRDzaKlKNeM0QsYKr48MoxO+IPw1
BMfO0WHVUQ6aHM7XMmcEeyEcTQh5jkgo0nQs4th5uPMtzPMItTBwBFMNP5J9SNCtJc4Ift+Sa7lj
XHUDJnlrI1Zx0vuSx5RGj8lFw4K9S5Okjq0hNek9Oj2UvdVYD9LH1l7z+CiwIfw+AXknV58c5L1d
klPSKsmpkuISZIkppNHznpntGIpUhLW9C02AXN4XJiwmbW5zNaUG5W5NQmDLZRElkxBBXhkBfFB2
FBEwhu1a6rd5C8SwwiHXeeYMAMBRIVY3Ra8xzqwhJPqEQkAZ6tBsp4vNefrjhElhPDj0UosA1Eoy
12+HOvUUbgyk9QVSSCCzduhK81LeuTecw1pTCyRiWYYCbAKUvFBGHOJ+3Lfjb9i/CzyRRPhwzoID
0OigexhrDhNcnf6CkwJKS6oiz1nwQHYjalVV8mseI63p+hqIZOA1ioWZf67DXitIKpPeqULb4C4V
pkf2rpheofspU9vkrNzhwKKZTB4PgQh50H8OVZ663BhAtO+DmWkFBMXA38oN8/Noaw0EBxSiVmcK
9doTmUFT0Th1JVd7AA9n69Mh3rFA5zKIi5H5XfL0bWtlHcHOnAmJftIuJfaSlcskPnXEd0KkPUZP
QLQy6pIOy/V/9aD3IwCRg3L1rt4srCR9JzYGRbeKZ4YSLQ0gHRveXBd6VkbOXDvMWBR4/1bVb7eM
tJsjoA4G2JNKbSEl/yr9gpi3gQn91q61/FMytnDj+cbadcSLgksi3aSu6fD6DZPRv4R8sfXAxxX2
FkHQSRLYisSsBVJUBdkpLf20M0F2yGX5gG3wJKKNsgXEPWYw3B2YbYZyBrT3PWvdJwYTPBxJmAFk
SLbGOAoEa8brjojl36mL85V9iX0X+649W1o2CwX0p7giUojK/+1bWtgLr4bmI0V1th6O12uwSco9
qJUSaOr/CMsX2sq+IAJQ3DJUBqU3nF5mB8B4fqEACp0wTmKs4QHe/xFVXKJH9EYtTw4GhVQxqL9b
UV65iH4H8S8xEtnA5j3ojqRhxT55pJHb4n59BUzLiAjXDpoo1rRsU9UlKvEfUey6YxKsTyes+0hS
/5bL1VHmk5JmZd0GyeAA8D3U6xNvg4saV3iWv10s5gYN2NsWV0BnqE365hkSZpPa8F1iVWjRwcWp
TT9v7YrSKJE4BxSVu7P354QH5/8IxvlYp6de95enya/3msBcutlkB5RXVS4AOK3W0hxKR2qxsXkZ
Ahr+rBQaHPRlICBTbFEF2uc7VvyLpkjGR/6MpqQ8ooIX4aq6lPqtlVI8IC6bBhWrUvVw8l4ew8Uo
a3An2EVjjw9TlfQMtz7dihuyNdFDMZE9gVpNRpcZ3SGUUa9Xg4gCSkGUxkRDzWdqE52OUEuhy4O8
K3Qnv27ls/RTNA8HDZoFJ2AKnzoXT55k7GZdj0x1mgOQPke2EatHrlWRQch1U0j/VOC1boM+pB08
/HRPi7ZHvWC50q4/PIJ1fMmbrN56wdsXcGYVPC2wLNv6zFdDzpORZCvu/a4Qk53nNA/batqJAC5a
SZgwWXZ6I4K4JMkeImfXLR+bxXV4H6vwyBE/jkSDyxug7saqZzzAHkGdZfOiR996OryyjHrr1C+l
SnMajynoAyB3rNRdoZKj6nWpb2wNOr9W1WCJG1DeMx2Bwf6gd6EtWRjCEfDES0J7YyK/dM25Sc5u
LUrXU4wPK0IDi6ZwaQ3ht+EY10pC0FwQTJ4c+nLF97TrrnsLTa8lOQW8Du1yQGK7uoA8M7zKajqH
LeT128DYpdfmXDTZJIdXZNvDP37oQF6C8bmOH1lowX4p2FSXBPPzzu0sN1k3YvavRNBDtjVBQg7V
k/yuRaH+8eDvhRJOFc7dyRfyjBsDw7mVAqySagFC3+SBklpcAwUNXxSH04TyKJFuxVq9OX7X23x+
6mvg3fV4YsVZP+06l5730DYmkSZhONuldb05U5+CHF2ISe/qhPeD68cRI5GIvCwJuJuc5iqu2Dea
NJj8eLqv9uKc1QT6wOdcvqX5IzrwvET4C5EnjKWBg0FO+GNad2zRTXyR15+0ocN7luDErkrrNYq4
t+y2cqlGEs5miB66LIr6T0MEg+75weQjdzvDEqBhcqIGeCrJx5CAWiDBZfqjdDo0L6moKvFjevY5
/zuRBx4rx7Lmtf4XossRmNP4WCyx4AmZNGMi9SvVI43bmTlmNNT7gjfOMZUNkmmtHgXKngTQ2fTN
WQUbphtDToZBXguLu8OoCjTr4g1bKEE23z1M9tFgYRlXpaULchhRWt/wibhB53QKUeJtPv0fV/Gh
1RrOiGP5IaGufoDP+Uhq1g1qT56+8/HsZ+onhJy1fF81MLQ1zbXJi6RA/oY66RwGxxnbH8Afx6uN
pb6bAcGD/4p9Q44PldZV/51WeQUG45yBXGcPBL5i6AKci8h7i1xNZqaKvwR9ZfwhuezkK81aPGFX
rSxfLpyQx6ValicnN46374ZpvUXplK++DWqxPLyWUAAm+XPOQao00L03eR1WCe/TUeoiUqP59+wT
zz5KOZkkwnjZG1+REsfL59Had/rOD3MGnCQQqMA7ErA4n4OM9jAVg7C5ZibBrfVnKZUSjukUbbUr
pv7hOd+iPe46nP52kZ9pGPAyllO3F+ktr8je10HCEtACxaVXalg9BP2J9pxzV8ABhoUJ8E0033OI
LB1D83IN13boUk/d+8X+VIqlAOxqrU9Pz72E1RdiwEc6WvktbB3erd3IveV6iVVl98fX5wrs6RWN
Io/ZuE670TPFBWY3zWmK8A5VNNbVAy5hREIq5cwxOsc8cxRwh9g5y9GvfOdh6v28N1ppZYjpRqpv
CiCPMmAhlptEYqu6VdOtJPp6vZFgmbSrBTK0WWcf17dxBMKpYxIMWcwQCS/Bu5qBrNU+6XKANNfb
qccdvmC0w3ya6wOSEC6vZ+2KnWEHAyNxSnRtwWzOFsHCcUslmfLhnAJel7kzRD54ejjk3EvoX/a3
9UeYOPztPli1/Cp1sRZwnu5CDBPK1tPcMxEwavwXm9ePnFh46DRFEsDjT/5vuXe0GIb95TCZdKiP
+KOfJ96AsChx8sMWX805cmRd4S+RgYh2G7yours4pt83AO4zJwG90LkvIvf3O8BFHfZ/XBjsDcI9
9OvzWkKxSDFwJ2HH2olS+MiciNdM/d6VJiJbxUH2lqXpsMGKhPqxnqgvgWd/eQGIxpuAeaQrP1KR
xvMvwUcIefWZs2jB0kbglRxZcklXJRwU3e9S1RACGjjU4rNoOJWPyp3cLuZp6TuFNzFEL7qsQe3Z
+lkSiReqUTokxugiUTDD78qCSvxQVdToKmYvbXvfnlyeWgpxaRFvsDgFXAqVA49X51Zzb5mfThCz
Aby9J7O1fbiVsP+SzeS4T6wTofb9xLfcqU37n2ieO0sEOck2yYOCE268nwL8Io5DUhth0jJjmPuR
6DubN+JvA5m/iI39mtxVB98U/UMBMDugSKkZm6HmQCqd2YRVgSjtbkYmKDr8+HGRCsiTzDD8CRtv
yZlav2war7iwXADUMh4TjHyXbek+p9+MjRQ4JuuCIxN2HH6RBSvritnpkl/IbSG+ve9dKVLi2QtK
3DsMEdhNFHiUHGHgGmzGbUXujb4BHzETjeVh1h4hp/6pLdD0Qk1AIRpduyxq76AeBA3CuOWeBrBc
qjlmmyiaHYbwb9Dd4ObdvUgRKCHDYZVjjwdpsETvDQ7AxuZClc3lyuNlGuN2ADBqfbDgnnalDcHe
t5FKFJdzv8qWlTzP/18Q+23AVGg3PFn+yXefqMKlqNn0ukspuLHYCyw6H2PRTJe/VCekq8czAkQd
mInSTdiEGUdo5c9feO1RH7NrmCq8knHFlafWq8nbty3XWvmiRBAkrS7HFUEq7pme69OMZHDzQo0d
xoXUZDfyr/bboOIA6PbOV8oOMclq5QabADe24vUAOP+HcZ4VuXbAmLuMSzHRtmt/cRcbB6mIlnbq
2IlDKSfr8qH0kQhN5kMl1sT1mfeJ4IIavOhoDlFFAgp1jWZr/F+qXP5BjuZIVmYOg+VCpAE7xG9+
TY/OcMF5I9OvXNT6W29K6NctWtTtF5+O0Jx6eJDm/ebMSFnars7vOZiaYP/h9YBYx3LDS5Pxph4X
yXasS/buNlihRUZWjxsIJaHlA+Z4Xzyno1Oe+xiBNfSuBt7svUCabqCex7byRyWGqiNv7UvrCFir
TzuXjO2rYiVv9ntApQOBsLK2TNrP4BMVd7fb04Qz1Q4W+UQeTdxYsgVgPttw0hQgvPjYmqpWjHAy
DX2+CFuPjfxE7dbKtsvlktcBc7rK0J8DD8ZpTpGpbKWWFIAWHI+drPTqA0YyBv1naXTvNoUgUw6J
u1melcdZxKqjJLc+rP2oFRs1+n3azNrqxtEC41hcQsbzPSKwToGTfGMwwlYCtab9X0Y4+ABHr5Z9
WOtD/GsXg/Yj4itKz3X/rcpfl3MiJcNvDSApE9F6PDHxm9VOAixHzdXvM3qhaV979TE+MAAeYSYL
0D6Q7TD75nAdYNm1Ec+xTOzheRlHZe3NadXVzyAYITgLwtURqzkHdR8grHdrv4SNcbi2TCzPBX5J
GR6sPh1eGkSk61IR5l7QoVCWVVDUfuz+4kVQXtzgTVuG6LcmmbmGOdmIj5F2C2jA6fbOzbP86Beb
7FHziDOQPSY0k16XpceA47MNjfNvo++XEuzvIRSHHogctk+AxZ19J1Jbaw5wLvUBWLgYDtlQfJDm
sFiESwRXuCA7+rGjVjtXdGud4aP0ZLYebpxp2jrk+2RDGAOlGyzz8CirDrEE0JhqC1QbfUBUKbFx
jTEiZOvDQ0L+VrroxYSRXTcmQkz2DXAoDa4Jqp8RWaFvYl2BSsTRpdAu1rQurMJS9ZKnwZAQZsQP
r/WTWwonepdlwJySkB42/UFMtWQIuaN9m3a7kX2bSA1+6s0aTp5zvOImGeZ2Sh9WylR/q5d1kU09
B+31nd9mzZNrjJrP16+n8IaDhQsK6jhCzaWSSNADq2nKrjmVEoFkE0WD/0KkYjSP3EuwPdGmHJVM
xCQuAma3Y5oe/1jjz/SbaGbahAezxQTpaWD6blEpI+s2hwRHeIsjydnNu8ZMX/zhnnmEQOIwFZzO
xojCrZ+T7/otnSm3oqz1eJtzmTriAC7kvke6jFRI/QLqwycGrNBBoM5R4//7W5lP7xFqMqouewtH
YYUnJUUnKI+4adGfZBVOIgr02MioLiB/EScobVnXBG1Z6k9DNAeSpTha5V+c+DJLFfsl2o7JEvYk
h0nVGvbPJjtCR7WOGaG8wTOHtLhSnd9Lt7X2JDly5tp35TBc3AEqZTTyL6UgmezqNfJ6ffehb0NJ
f8t8FqxjJNm3fc2hksznL+5lOowBH5TX43uoLlcMF4Y2CZJ1J64d5FZF2kdClOkwfooi4MaFD3mx
SCj5A7skN1Zc/wTTkzyICEPa21usaZff834UA/J7kCb90Ltb/+7c3ous9/N8QkV/hfFWhqdOWUND
bMsAd/nVE5h9Q/KGhpaPdxAdnJ2HFw/ZrYcaqVT3F8x+RShFZI3Wx9MzzpkYmIoSgBZfu1ZRtXLZ
OmuxOZkNnijLpbVdNQSkFLn21z8BVV0fXSq0FyHRn/EW1SdqItHMRpkHog07j54qtYCWPnXZTHpK
YKJD0PGolAdKeeiN0lUH2R5EToWzNBUzwjPgqyF0CCVsVgKPr44v1Gyzwf7B9g5CXCUqEs5Lp5vZ
vDNWCR85TazUbUFbIxSC8SwZ41i2GWzXBbxEZuRyWDUi/AqMLvbq0VTcJ0yjUc/MsMTZd28Zh+K4
OpYHSSMERAxfwoSoqkfcefN8YvMGB7t54rl8c258RfKlpecJsTzNeDwmqwKtU88puXBICamijVjf
LQyir+XcIE2FToEa7cWypZm4OL9JOoT8VP7M1RmEI6/rQXEomLcW8372EPASUpUJJQPVHn99qzIn
szXH23stPoRz9Bh7SNR6gQMPXdrSsfLyFdz4354ns9x9nQ3PWMkrMTb2iXiD70DPqhgqgGX4QOyq
arpPJD6mCRZq2Xkypb0Ifa7ZHZLe7weGGFNy5LvbMvMEqYA7eS5NoPkUWFCq4yKez3C6QXnhbDcl
mLYMax+RWt7evnORZ7uRMqHQlJ0aaq0prXf7ZmHoBQHWl0l198dsBSsWyq3xWiv+rGNX5yrBH5DG
/iO+2g1XuPvvzDQolpsChL8Ds84uEhHwWec43/twGmx5Iz/i8geJ1zRadqCCBZoa8mZ6JYMdrSrx
VzoIZF5JkD2wugogBxCl10h+7blVtS6OeFTVDCuw0CQjs2k+DZhGfxf5eapvaPPb3HscAkwlRv6G
hMu9XuhpccP9RTHqPj7D3UzvfeV1+y+cvXBWZDLd1fqEPkfkZhUaQEsog7coqYhJQ2V0KS6h/Gnf
gNNc29NeINbCkEFI3K1qBExtf+wqE1eiV9AHreBvLOluczHWFq6ARfMNYN5F4OBCgjdCr8FPgu3k
/Qwj2nK7dsmatgRCOBVc/oFdfwKUfoYZ/KkFnFaRkzFdN7WlY63RXbNDbZObhTatIWWTTINLsvsw
0Z5exYwDX7MTT92oO07wrK3kgBXFpYyrONGFZDfaF6eG70qgh74WpXYqWfP0dejzMUG99L3IcgVi
QLwK6n/wJkYcgM87b4jXsLV8/UR6BfTlzdlEAk0IMpL0gmSMyuIxyWBtt16EZkyltV4ifRqKtaeu
JEm1Nt797r3CGSj4b6VSoe4elUTf37RoY8r0AuCYTO2XIvF7ANZBbu83BOgfymy/rDq+Wl1rFsv3
eEJdX/bLuIy+KfW3jtGZLAlbywm6ZZjKFfRFo525s5zeVUny/cWFAmN0KwITbghoAcSjU344JWTV
hYceg1lcX3hsvdwzq9/Nqm2hlXSajG275mOOg5/VO7poqMHwPBa/SuuypMP9oN9ns7fAVM7A9RqW
10Qv33792uJdmKqUGmMDkYf1JmTURhwmhFZ9c3O9eaVVZsnOoZrEAjBnx0q7Nxv2hF3bTkAs62/F
JDUAMitKDIvDqAQLMfHXLB/QlzAxv8IsfpI+lZkRzAfgx3Y07l5EBuIGehhULN6x6leVU3hmE5bX
MO7g3t/WiR6OFBUfyXHXDAcHeMLMxstLRNyhlFyQUcXh1hwrNiMp/WMwin/n2cEaZEMJhH2FhSn8
Cg0ia53D66tQc6YtYzuIle3vCnyZyY+wDZEHiYtqwU0Ty36VkxlnbdZIAK1I85z2iGHcasgB3YOF
+F/MYngnl/EvGpODs2gDJS9di/Wd8QN9F89FE/esSbquoh02pMTTYX6Bsaf1cSIKrP7K+KDloL6U
eREB4j7agfpWR9dNMmAPM0i1cwLG/8LEZLo/53UcjLlysLrOhWvi7+yE60vsMbva3J/NMuhrRcNp
3cwzg0BC8JPqelxkU3Z6K4/IQ4nypE8sdzdITTulXzjC6uWINdC6dHCC2pcUNXp4fVTRYKZxSKyI
4W2J8ugq7DiSOVB3HHx5HtNZFjObLr/myQGpL5umqr0kGF7bbDoqTA5tbJC+2r1nRN8wi5F/knrF
Eq2MFMzZmbWeqQy2pqp+IjpbaWvrNxcz7YLO3eQt77Jz+6PeZgAGSseruPXhBefR2bzBTWl87Bhp
NTXNG9ehr4DMMupNRhvy6f6yLDJoCXydbtWQxlbnPPqUlo3d9MXUttpUULUEPZXjT5oBa5zC5Rwd
ibiPfKXw4YnCV4JpleDEI9hfVyCgKkd77Pbhti8eQ+hgFrqILEnyDqSP+z6wdGiAlqOYPx1WEOfH
Meil+QKRQ8moFeBLik+OnBMbb2v8+3kOOEQVDHAFnA99YAn/9YLkcDU2BFxLbXqtX4/6dTRuokxO
sKRvTgN3ETAgI4ukiQaYIOUsHSc+9J+vmYbd2zUwJIhSdH5QcD2LKYltxUqvRxpCYQ2Kjwvdc/VJ
jMdsWAITdImwZ71iqAPwSpFDgawrBAL/L/7ETHdKSF9k+P94aofwe18WLqE3c3DJdrTUq9nwS+rA
u0d7f1gpyXv2CqkNW2B8TABsQAKIBaFHHOrkxlgDOuE7IRC/Gckvahx/Vu3tvG+QwS9zpzutgjvz
b5AAER1A12XaHwk0MsDsry8CsJv712X1/9Rw/S9VFc3iCGUwTpu2wP5xs6Po15hkJjdH5eibnp3z
eGRrj50ghZx7V7vlTMPvOJYn265gcPHV7vGN4W4n/DDw2P1uQ/ytTG4LwmyzArc8/61u+KhV4/y6
NBCWbBfHyNLgrqyPK4IBFlRXy39HdTjby7Ks6nw0tV5P9OghSsoYaloD3MkSr9kwuCgmoye5VZOw
KJ2v21flcTyODyICFpKbDRkUZcCC2vcgYbsl7l66mEVfxgm2xiLI1k4eh6BYNoV9an28qbhqiq0z
F/fvUCcAqEmlfH2xgq+yD3hewAFE5OTo/uRJtBpFySyILohfZM0Z4bxgiHy2GbSpNWAwGE3LGBM3
zHCSeEGjl7aKRooYGq88LDvO+ZjLkpdyVMThp/8OpHCG3+PRaIk9ICffb+zBMFUAwUOH61JdUWk5
N3idLusaomKoqrDv6VQgjFUDGuvy/75XLloQCb4wARRdifgcsCVbQSFWpK1jM9Yx2u2Z8SrLZsMO
YlMrJ+KH/8Ua2y7WKQL1vrBEH5KQAOk1IVLmQzzrovV0qsUQA+QTRK6PmgHW+YBWAnFsiaXocQqz
y4OrMfek0cIa9Cq9zg8Ba+dIybb3LXv1HmFzWApWIHvhNRgxxpOJhiDzQ3p9gsZ2KhdxNCwUnlfb
GUziuCNtfCzGIkMe+vZ2C+U6NPOANimYe9JdEe5LXmV818lQzaPd3mWH5Ayzz4XNToDJRjM1OiXA
BYiIvdM2PvzEs7FLV2i07gm/4zsyIRcewWz5b0V7VTKs4L7JigLShwRYtalVILbKTVw+SHnlb0JA
l5fnUg02nkRXqc3mRygRs9mF7UhbytkKWe/kXvy9hllzf/l0iMzq5vuNdiMl2mWRAfRns1hKvcnG
8sRj45tBfRxwwErJk1JxLrcOHmELtkMC3bKYQOiBFCk9uq5Th4sghonHJKvbm/8lhzcg6IHCvjdV
btbe2JVxRr9RptDbIf3QvyTZisIH0SuXKqadDK9/5yp7Z4JqMnC2HkLYWbH9i4JTjNdkFOIslww+
OvhFcj+aRNXQy6z0KLPlt5sHVPbC2osB2rsMYnbSDRjX8N56fh0q0erwZxj0e8pKuAmWVN+fSO8r
S5JDcZfmoeGWhiLCm1jW0FkbaDppTLVKH9j+AwXoiznhPWFlAJSPHwPGeW+U1ofVqy4fXukOmQDj
o6JWijZdpXCrVgBkVLvv1LwSSpu8pqwD0B+0v1ap0mBEbQKoZAjQgSWGMCjmAQwv8ZjRIRmMHEM2
jG6q07iIad5NgMpSSATQnvO5wae2Dxsl383aBP7tKM0njHQVkiW2N2/OMUbSuyFPjZ9JpBKxJTxM
cWR8QdOsq1g2HCqcDVqBLpIYpZz14Zg/2xEqRQedACPzLdJsY0SEkfJ6VwXsAfh3ZA0w1hQj8v2y
k1r+YrSKIiT4b/Ur+Tlb/6TEg8ZbHWxpj0I8bl2WllY4CKUiRmPet8w8rVC9tUGHXS7GWZWELvIK
nBVB/NtLtzYHuM39nl+1sVQu7gD8/+x04Tr0rICQoN/tPNJqohJpZXMJYgjcb6fp8LpKEHKiHzQo
1siJxYt7ApJLHOfEnXL/TEcMbsVZ5wRYyNYN8dIem5O39V53e9AVs1r5ZPuqeTeklXok5hGYXqwb
fODpcZkj+lFZTNyXdxD9eghHF/sBed2XVGcMtAZZCgZPJbFo47Pjib5j7dy0g2kvJ0GyvRSn1kZw
p3+mEhKL2FpNKSPdNSH04I16oIIHgQNLh8DzBctJgv0SSJQjNDlucPvrwigXk4xKYRQQCVGkFAAU
ECSnzcuQpQz2+Yc1AZkp16A9AF/larailI1iHcHzBnhQwcisDPHSsUOZLRasOPlYbqNeT57d2hQb
M3E3N3/SFxSY4otpLdHMMmUzvfFpB1E0Dkcnyoah0o2HdCTf+X1TKZvtqB2e4SLEk6kviNAA5nCh
tFpnflbz7BRNyxlSAf9w1JkCnOaO8lmKMSlx42Et/HCtx3fbHWKR+msk73m5SE1wTLeUrf8Sbt8S
JcyhKeJ5U6Dz9cYVAIb3dmTlDHTo3YoNrjQQRs/7FmCTxqzZq8kfsPQN7Wnw1pCaTGkMUgF4B5rW
v4Fggvt8Axv0FkSpA6x/g6wjtdkEeLa0vdfeGXRtqhBz/nqddEBF2Ls9FCzqVjNDIPfnyNwKas2I
jem+N5mYJR24orVjmNDsgLVjQ9O33UE/pZwSW8b60dVCFLfSJ3SuA1E9Mj5DQdk/UiiYNYLfiVGM
6FH98k27soyRsrz4dZHIz7FOyCW9WvUzpJtO5VJlnbd+22/VrER4z9Cs6KemBpyeY0nbP4TjAWM5
SNFvb6AMivS9n90JlIZ6kVn1+nGDnZ+YWc+kCBLa87nWdSf5HV4fnoGfPzEe/EyTCxSKuQ4eyFst
CjenrgFOZvwy7o29yChZnf7Jzu07JpEgXzfMWOqeKUxJtxrdivAj9VSYufZxV/zD0oLpfDjUNBa8
C/t8sgqCm8UsvGfKu1rFuy10zi1H9puquaI1NF3sUSU56HDPoBz5vYSIb0N9Dy0FaYljpaVxjAVe
u28z/Iv/QG9FsNqYQUN7sc3NrYbwCXvUSC6eFktEZuQb7fT2zo8UaR8dMwrbzax+vqLweevrtip7
HBOvWbPTzjoQ8x4OqTDljm2munJ1haVncdqgwcn3SlEeku3xJB1RY3B+/J0mY2UGN+IF5zWpd0BN
SwyyBjBqzajTmNUSG3CkRqE8nNTIYAxP/xpZVDFkiENh0nki5BTvEF8wTpWVG6Ej3kG0jRtmckun
WuT7qijBY7i8sOCrCqYB1fcgtDkUPeJnm60YumzUWzAhEN0RrJS1BXw1YtmoBt+MPq2EmhDrOsFj
yMb910REH2vlvFhuj1iRCsQIUHSuBmTzo10x+J5Pbnj77eWg7o0Q2+Y+hANTUgGIlU7/RRsKm8Tp
YNv+3sCUFZHU6ioSxsfXCeIGhid8RTextI60wEQSinEeIP0ku8vEPxPhFenAKMe2bNdUStrkXcGC
6k+nhiey3aXbRC196a4WhsHbm64pAgWBlGDKPAF6ViIM+EIgtsFTWF2k/fCnMAhqZkOvQJwHvi2Y
vPQaQLDnupfmJBGJakHCdi1jZwrix1/YXeVI9FthEWOfj7JADz4AVAg9Kmml8i1u33O6soYP3n4P
cyyBj/7ZTjg8VHUbHAJmrfXFppqjdCMpOxcaDi2XP9ZgpfkIryoQ2uUkfZ3MztdeDp+gpncsbGdC
z+tHlmqVZYyWpjcUd/1vSWYwIAPeZ33FeaJUTuvW96LKaOUvN0SgNcg19/cR+DY3I8c0adNC7SgE
gBH48r8qkSmxLbUseB5w4IH9mpr5PfcEEmv4drMPGxDt6bUvt9JNNsSbhadFmC9iU4M7RkM8miP5
27LeRCt8qCD5RWzhzGjDDdernakmAXFT0gDu1g1tkmSR887PfAS20GDdhtFZDu7RpxjxHHivmXQ9
OHDiuqsebEm4Xwn1FehpyngkhQX7FMH8pAZfKZff+C+1i1bD+AcXVUSTUUxJaZY6nwTZJ3RK9G/q
oKBj4+Mc3N4N8P/6sjyXfkAQhtElULZ4GCx58aTEvcd5z93yN4WJ+cOF24dko/HeqnBiBLye83nZ
Zivgbze4E0AQ8uJoKW9zkAX1FDwKb6l939jBu4FzQhf8p2cfFd5NZcHcetaboizBMYHlv+1226a0
VIa6QX8Yv1HQ2/qZsoz2e4BcdVcaDEcclMihzarT9BJZcj/xtFK6r2q6e0tC1bVM4j8h5Rp0/wY7
aIGe3pQm1PEFfsxxxXTCU7a2LIIBuguvYjwLLOXmwp3RzM9fCCgf+svPUuDwb/8DTOIX+0mQGN5F
JxzcUCKxE3pLPnOpNx/41mzdOH3odYgij/firyI6xTRv+b7yF9MMY6Nm73pZfxwxlwmqDGSymHfk
9iTdhlb9vhCD1k5JoF/JCpIlwZuVRfiUAQYzgpd5k+tZd7YuFD6ZBV/bbi7JN1IpH+njN4cJEAhY
7tD26KDyzfrSx/QPSsjQPtsQ8yMRpLsyf4RUJlRrZcmUpnMCWnXeZI5KJBr0NyZMcAdW/SPdTA4Q
3eEAMvQm+vo9qi+SHAXqLq3w7ImQ6aP1+zKuZi9CkcMz8T3oJWpx3sjXrei0gjhaGM0A8Q4HvUY/
NJakFKnbYWzVfmiKEYmBJOStVugaFP1v5q2jfd1qMhhdrjVsNEN+10G4yXX7NPKIG7ccUfOV4g+0
rA8RTStTlPM6DtsKOra9oLcNWfghvjuzKAz9ozagoL/Uh0ad80C1Fe3Nn0IMTV1LPrbWIpLaDtZk
BJh+IiYsUoW4yhMNd+ifO9Z9ZkBrjIP1v04bbpUay/KNA5td9P9YKYjkk2BPEmW5GB3+YPlfHTJG
z1ooHzm1KyRcfu/Hyc1n+QSA7de4E1zRYS/W2lgiuvWov9NJ6jP0/BA8J/WBaTjy/6qIDo4KxNNi
F5nCsifS701kbGKPbKw0npkfjzxkp8SiNjShJkDldaSOZCQFY/7y3J8IebSAW3cDop02IAuABCUb
JGbvEpjYH4qeJH9WLKEPjeU2BocSFUn8yYQLMCjciDYbX8imeDrjSpIv6hKYUbNKGCuODIa9Kr+a
GN83eRy5qOA1FnhQLbDB4qcILj1z9I+GjRG0yNNGVmAPeQL1xBRhSbirFtYLameCW/YKySJjrRSj
tPofBsZ1zuT82p9q6Pn3yGIVrWQnmMHQo7fsJV+ipdRpQtYgCsWeRKUrxK/RXMWcSjBNayoBMFTD
RRKioNH86N4TVVMSC5YOADCZNLYGlnAAX0QzfYC46CfuxaX6lj7wuP+LSGUMvD+y/HbWNVl8mG6d
YMjlU6sO0zerB09gFCG6o502ZF1m1TPThHdybe57ikT/sohRnPXzFM0eor6OKqq8G5r0LWDiz/E1
hWmABnUAI9A0ASoUIrwWEay81Ec6pbvSjBEws/sRtDP38xxgx/iC2r4HcRUfxGQA4Q5tt+bU2LKk
d4UvkCFNoyT5CbQYvsRZjwjO1czkSJmXRspGOLS9cX+LFnZ/m3LX0KczIqufRrowktaKE1BBDSsb
8QN6nMdiTt88e7V6P7VAopWT7HU968b7PkjUVyAMtrJ1TL4xKkXg9dohVUjKvu2J1MpRKw+Qoy8C
wX21jrqN/1PjcPbwdeYiB04Fia6lrdj4Zk3ewwSUI50P3naa+FYkwjb9dWngMfWOu6q3F1AvCYK9
LmeUe+jF0E5gE6sUDnytDuO12ESbnQh2StygyHGcHqi4J1Gl/8Oo6u9llW/hMyD0QBtf2nEAazng
2r5SXbdfLbhfEDBK5cnR3zYECF9Z39Z2dcHTe8eacWikoNUgkZbnYPUhj/MheN8qbyxEYoYtfR6H
p8wRnp071fQdQ/YLFi1kRAcMsvhtOMR50DgifPeaJPAfdsz2Dz0PJlNCIUEx2z6KPjV1PyrBy8zY
IVnFhJFDR/XBoxG6BZv3q9VpDWaA4PKg/4sN7XlZjvUAh0tFsdaWigfslyCnsUHwXKd8u4C1a4z/
7kXK9QI51rlc7zXBPcLMb5+TfWf9acoFuwN7LRdPouzbr1dBDm804h5400yBqRKJJ+LDId7ju2LR
H11zZUjN9VsbuepFWpx0JZjAB6uxm81ns2yVYZvhrp5C57GQN1spBEEw/6xB7Bv4f4Tw/dDQ5LGW
9Ta5nyc8EOhDXFGzbAB4OzQnHvHhCNwta0sT39IVsMk82ciWfKfCmulcA44Ne/q8Ed4t9CYpeKTB
F6j/xiAKNsBq8DkYb/M/trZU8X3GFWmnemrMuws4B91mFWOayDo6TpcJj7eWnAtAEeEuryT8XrPt
ulaQ0vsC6rziD+tQION4FPhXNfEeqn5pvPJgCBEUWHftToq/Y8CAOhnTfqR438ZFzMdBeH9eiIx1
M3mibQQu/xS0M2CZvbnnzC2SojpdILhcA50XGFfw58MkPY5uCC37K4CVyF6go1mZ3c0gMO7LdReW
xPyPrIDxnNH5NbkXbU3Jzv48WWzRzTccVs6UXjwjEBGRk1dl4DQLZ/EiWs6hLAaqGQuz3/p3yzMS
TgOTTIrSXA9aMIfvJHb2yw4FKPhVJugCg0U53FFz5V4HBN62vGGydusPKT19ONYfqhLAQ9CGIlOE
mE5xtQNqwHSP2LJQGFd9X3+g4jvpWvTGRlLkqwGNL300/jBfKmnmABMj2E1ZQpFLFXHuSQW9nj/z
kXJPZlaujs98F3mWXvPSEubzZ2JBkp/xpbaLzqZQ6fshYngMhPAAfHXDU4xDDq7bhSGCN/eGyawx
gDVR/RGgqgUD6vq/zHZeDl0quyp9rq6F4lcvUT+GAXxrCu6e2LrKNPozNER2K6IKs8w7AxN13Wyd
KZ2fcWTEBy8B+S1L6iuvk8XEmdtGHrpM9xA0Tn/6fwo31Qt4yIGIwknZ7O75O7q9ZTVuHg/Puj/k
o0yKeMrID6/bb/2SCLOEztjWcPKRE5m9qruyyvEtqeXpSIRq/COIuVJs1MY5PjNRTtZ0NwZj0Fcj
fCYslQIVNn8rQvTv8AOBGBVJ8K+Qo5Ofkbii+mvhljU71zTY0nd2DfTquYPV7G7OPKMVvbccRPEH
I+4OmtKdsLWvS0YGSCp1CcwGgmY20Z5PHFn101lVXXJnaQXERnKsfMJuRq5ls791CUZNFsCfXdvs
uBUNXOSPpViqxBdqOztipP0D4fHM91sVfNDdnYKi2F/IiWF4N+GHFY21SsewV4JUWlKA2F0w5OJo
vQGYSbPJ6VM/lL7K1nNvUdhfvuvGggc8k/+n6ScnyqOLlugbyolLosmXfCcAD/TbrHY5U7sMA0vr
ggIEjJpqKJK0ccpj6w4vtkZSSFtgZoEPup17X5a8zzn3IXvDRe+4hfCp1xlFjAJOl6AZOZ2BTrtK
MAEYE6ilElXJFQ8ZdXwtbcpqKZYaS6CfPvvsI43pdJDBwyOT2J+ZQVUNChuRQHKfTyM/c+ms6bMp
Pd/Jo9wrI3l1rX283j8pDDPXmtGuaU6MXsdnFmgDMrv/czRLxXS0Vs49yaiuMGR82GgfA/WusxVo
YVMbPOnVipUCfRqHOVLxJboCUubdvVbiZ2+LeGXvTHBaYlmUD2m4iJ+oK0+85/DDvuV9+l+YnZX7
6TfEwsea9csnFt7hNvlpZGsg/o0YrPnhONlmwTzJbfe2Y1LR/znIS8MzoJEpigc4DRSQgdLy1BGa
hQy+hX3daBZH86oPtnVQZeS+6L2PlqPkwyL/Nqx/HJtydaGSEX54lv4TbDpNoC9CDCcR5epB77Ke
NQRkpIxsFGHI+0Dcl/gVejRJawfnlc317UrPXv9WMqneHg8EejaUMvgkcZYR87orOzM323BSeR5k
9e/9dRh5EAVNuLIvVczcO9B+VlvYuYJAjYLvF6IYpS+gIUSeGiafrHLlRvzi6uCb1L0Nn7eIWBV2
meGe+YIU3ZXn/Tb9EyykeR8kkt1fGaIQMdAiD7NeNCh/djxi9gJGFjbyh0vnAlXAEksvr8U7xBBP
PhOT7S/otqH+relix4TYUbuC/4x97L8pmjhcgoad4DVlxxAUBz1ap4xHp1Dju8Bn+Y/npnMGU1kR
Dnz7On6yytOnmV5q5Dj6thrpG8DoAs+bS9iysg9K8Q7HpM9RHuZkwwXIASapFMRPfH3UvRSmxQ9N
vEVpuz1jOl1gJF24K6TLCqht4k5Un3CS7i4I9ouEiCQvH9BJmSVAsAlS6YA6s0bHIaYsc0Fp0bp1
PhnnYLzAapZ/4LkIazviD+X32gIMcS9WNnOzOQ9pJwEnU4laY5X54DE7e+8Fr4IPalnj5mjb/dkf
ZsNYD7CJJAMpvePxEHfW7Uj57t3U2Tsuwh3sQ+nc0Q1Vy72aWHeO+x1iY3sf8dR0BJccYw02IrEs
pjApOf1FX+mliimytTirG9onqYVJU7KATUunb4K4vYirHu9FSwn9ajBPUAhOL/nrkj8kUDmWWqPG
Ek26PpsK98AmLPebR4b817bhfM6e2Fsbdxm3CxadnoJSwQJhnfyncFft+XeyzZWtlWuzdRQYZ/8C
Cr7TEqLVmJ+Ocllx5YmpWSF/Wd7iqXwcomTBhuZbqL/cGnIsyWpGNOb9GFLtGgR0mh5qnumN6hMv
b+fUBc6Bj8d9sOW+4yLc6qXE+Zqxk9iVFAE+zAJETW22LRhpSQXuQSJ+ZQ9KAKlE5e5GgqI5kHEn
2+0OMMe0i1MSqU1F47N0LRakffFLqw0IP2qauqL8S08U/jh7oJHb14hCFPO590oWDi5rQIpHwZdL
BrbAnf789Rf3xl6sFQasGDw1dDfL9vmdorp/p0zZUrRGbDrWWbdR/Sku1/zEUKIb4W0I4zKPGGBj
gOUDG4fwG0dKEAp34Osxdx0CokosQTzZthxcuEGdh0yl3OfLU7rWIdL/hUvjNwwHIk+VNIyL+EAs
1tJvCLH10N54t98ebePqpZpIDU3oemQGBuh1aAU/+p21gqxsS/8U6iDLrgi0EBJivczomg33jU/e
2TWNT1hcGcTaaj0KSdoMgP0g/1O5pfCEYGaaf+12QEDEl+xrf+l4M4np3fDnqdcYTLmCfikIuQK7
P+DJSsKPCWWP/yDCDbGvzQ+QMlGkJdikCcgSTy+xhtkXbYP9+BZMHu85C8FaynjpPcloCdV9t4Kx
7wxVpUsGcFLqol8U1Bv+1osUK45vJVnuz1ziBwubGsK9KXnN2I0I/zfNRkJPYTSoMixAV/Eqzna7
uBYj/Rr873kP75p4pmcRwnt1pYo2Vz8U0kfkDeaz4gHz+PKdC2zlFFOraI2r96uH5cxJ4SZeoOEx
g7QTHLtFqv61mbvIbmIOijU+ht6e4qY8AyRB3g40RNF9qglxpDCH/8xcNTKjLziWi/1eavA9F9GE
f4pXQPWBV8XgdE3ee9zJem4+PmWHr6zXrlKu1k5vglJMw7EYoStpjyPY9ia2Q1xpq3kHvpU6MRGy
+mR7r86zhu4jOPHZ8GTLVBhojqWhbAQaRihzw5R4z7PSwKR4W2isssB964FG1v4R22eTThOSYUZR
mP8vGwh65t9qsDveM+jnXf9kvihqMIsnKZuFKFsShXiHKuask9/0BE5of5tdlflwiANrnut4/BYR
0S2G9d7PgBDbz89uFRD+VvfBiZ6lmi+BJrFmzLBSEmWapEmzG5vJACz1Ygfkx53HodpMkJ+oI8Q9
seS1VzLLtNKxPTVRFOpYmVwcOoLnJo4lLT+vgaL14idtktpPXTgxNjyqwiJBEMUz5KxUv0TiDf7a
2rK0WHQlvyaCI6O+Sw1UaU9ZWOsy3fuLMFNKJuV1IFM75Jv+ywYuif2Mh3nTjCyvMHHkMy/8zuSm
FgM22+maXbiQjpfbZI9SDUb5wq/GQGPXFYVufiIGhZCAM6jzyhrvW/28OVjTkIimCpgx+p4LRwaN
8U8OZTclbv0Arlk1E7Mm6PCF3xZNIvf/Xn7jxeXXk/ljmVi8Z5w19psZBGH3AKe2HiU81ty6DqJw
ecdKyrjAws18wULxYJ2xS8eYkjwvt/n/tcHA4xjFTuwiIDKZif+HIpfMnAqJe++/ldqjc5lbhSOo
5Z15TnMH9vdAMid36Rasg1TkWi59xhaRyXVL+tKsI81XQs7qf+y6HQpwq9Z9ZrhkPFKyhEvfm55f
Ofv3LPMZrA1U72K9Mxhv+mIGEd7/BhDCHNNXw+YZouU3KA0ToVvYhl/SlDUptyWk9ZqJ1tHoe+M3
2RuOo3GuVx8yh0GoY5LE9tf8vlq1sw/RLJBW+pRIpgCxC0/3/swjbjsipt3XnEiKExoYbl361Fk1
7gdu/2ng2ajpe+dowEzsPWl5hpMROcptoJDSYD3TLtIh7n9luwJkGZoN+QYVR+Dp2xZb4zQiqvQx
M7aDuWipqOHdGgOoSvxvGEXuzAe0QmAwa2L62n/sQNcUGMVYTJ8+EBDyBrbAc2OMJ0flowy+SQSf
OZKYrd/suwFtw3wx0i3BZ1O9D45uYQL4qNyJXxqbseFqxkHO9KsuoX9Q8BvG0sc3iCWEpMX6oJTQ
nQ6gTMjGZl0SJLFIY2C3S1Lu/GTxuG803UT57cC1Xw9EBMEB/ru+Pf5MzBCsg4O8X0BWkuNCQlBl
Zg0QtgEvYeMM7vPlfuQlWJSyCsszJKLuXYLDiA8hzlwxHlkol+bMdwImkThO28LZtxbuI7yB6zLt
lcSFXNSE8m77Ek1NQf/xttBiOXKl6No6fQ0+2OOQm6Cv/yXbO5CfaCX5kdXySjBQSU/CoXDzlxDM
S8gSnH2Z1Ml4kRGbwgIGGQu9DylgppTR5wpx7S/sq3nn7nY4a515Nm3rq8Ffndrn8ZhRQeh2rhZu
H6ygCqinYrL1W32AiRofmnPa1kPhZ/zUwLJYnZ60pZW2l5leX8277HbhwkorsorbP2dyZJoWTLg7
NnhnIqSOFj8QsppiYr7NwkUTyB+r7Uj3MbMfs+Qx61SiIlvQ0PXq+Pmx2BYHD9ZC/Z+MMfYgG9Vo
LYt2bWnYrBsZf4ZGpge9xuDxUNEJgVDEOSfZv3WLn/myAhQFRr5gnB14S+3Z4AtmGM9JQJKyaJq+
ufPCS/XxaEDurBy8mGlZWJIeD6SP4YSrqZeOCtmmYeh/OAfYWsQGwKpb5pwmV+ASXkFtZV/JxcZc
6Jrso1mwTK/lcThaOgsA9fvNhnz6ceAxj+EWoqsjZ8y1ynviajUPe59Y2H/Og1fB1RBtf/3Chhqg
HfyYUTlCSE0P28D8Hd/NdUh++ydq0FXvpQPHDwEcXFFcjwQoyziqQe8Wk5TaMf9/rXvVkDge11Uo
xPQAdgYOrmHGFuiASljFNG+FQVWdVX8LAI/kETqstnSnAHo0Jr9YNc1MGdiWUQwFS4qNsv8c48tQ
4RcD1c9okjzX449AtvtuX5PE4OgSED6EzNDo7Bwfb97pM/yI+TOL4hQ/oJzNyDigwuANfV4Pgjgl
n978qBlVSR54LOazJmlhkezhU8itCJbT0nyy7ZoqD7nfasprs7RJJQj5GHjN47MmP+J371iygrn8
YoGUu0Mb8aOaxjNe8dnkhtiPhNEBMWMN/0a8iXLboGy3HIDyqw2E/QX72P4v+skpoI80uY0etpcJ
b4kaXKPrvzh51S+9qIG/u5k37rGZsXs6q5t+TwMSXjlAQtoFSn7OT9d/nQ459HHKHiHVBTLih2VD
vInwFOLLadprT82J1E0u+fw8ekBwaWfXch8LZrdI/5fq+piegGWGA4E27fCX1wbRzprVp5s9aDcA
hMdaCfielfv0kw+clUvS9xWQ/Enw7rO1+vvnYbQeAf/gYT4RT2CKe8UkpUMmEh1SswO/cZZzvUbE
fTsoqIPx8syGkfNphQH4DaThc++gon+MuhAeIsBPem4M+yNQDxV9brjP6Fvhf5t3RM5f8MNGYQMQ
pPwJwI89c1kMDEle2Ob04WgsrGYQOqWituOW6ucSs7BBuMtS/8c1/upgju45enztlbpuobhVB4Wj
MyMuaN0jdYu2pnDNGL5nUHfouM55rr9ug8A4qF81VXxcg2aLbD4G+JSwW5t6xMAPlhhOSVBfypvU
KenfgUXIKSaC2qoFePP+SOQGqqWUTcUyiZTfH9J33KtCL1njXXphA0OAPnShV4G/ysxPQIVWDzS1
G0jITz6D/Vk1YLQfOy+GDStRos79OjX7vtWgVoAw5FRZ4FG2MEzL12ON+dJnSvYXyAcD//RXnpIW
6MfdCjJiFz5fwPgYlAjsxtvKFJWSXooVV4j+Q5alUL3RnLwP9xGFnMyvAipMeg01tGmnapXrj/ve
X+VU1hmu1HoNoCltSDaVB2fRZGarGRymSGIT2KtfH83OOgywP9DYzJjHWj6ihZxS3ywDeLZpQ3gv
WWTMEmNdz+Hi4GKvV1eE6Ontn/ILe00EepA1MPFY8b+u81iy5eL4z4ZkBHd2+okFyPP4XGudFjFh
umvkSWSGBTxifLBZmfLgO5dhQTFWnH1DmzR7/iiJ3JHSGjulX8n0wSND5xhK1AIui3OzSdglRb11
vqG8OjEnKhm/+ZcRejbLFOqZLLCbzLfjXdF//7xShh5dMu3gbdEZezRod6+6ypWC4Y5UEw8PPwVc
l3/yGyfoyfpgGSPNnPkyXcUVvmCDtT0a3j7xIR4M/4gCmYOAbhl2VQFyKGQwSPyALEJDf/Xz/0EO
rgiWAB8u3HA8W89hVHKv3Uht2p+X4uC9N93DXDKNyvrnx3SIrLADElxkmUynGxh/3eOjJ1aJDZ6L
haBb+Sb/e1rmIJZ2LReX1O/tY1qe80tXZa1NEOUl0Bt8uzPpK7MYtXlKhc0ME3913dN7y/GCFLG9
WJlu9lPrPHkFlM1xLvHC1EkW513+DPv0tVDfWMHd+/RJZgDUtGi6D8T/Fa2yx+Qk+0Pt7DBA4UPZ
Y2Ughdb3pDIDtWkCzogrzTGUh3Hwt3OBTvsESjA+zFrf6fWTlAL/OaiKc8u3TysaXDxUjJfiHpxT
fnJAg+zSkO7qHL901Iuq/nYNy5YGA0c5XirM08+bJVEdGudAJrQ4hRrCmfXpas5hGtdk289tUbnC
0ewwXGuJIAyP55/h4z4FZ/+XYQOiX867A29l1TwN5YI3xrZyl+82Vv3+G67Be/WOowJUoSX8Ro2P
wA/s0hfCajZOrGVjF0WhQarK53XcM6CeI/wPvWjigd5lISvCSi7YXEUuDZeFtyv92AYakw+gw2ns
a/kIUWqqgKBbqATaj5g6bB6LQ9jNURKz4RcT6wYue6esE9R7i+PKWRWEWSl+RY5+us2aKh5EIYSg
TRkXXP4tF7TDi07yPIF5heM5r0tvOlEUBShOTfl0BqZnuDXrFWoG2bDMwCw5LnPmRWsaTWAmasBC
5Uzw5qk1zGW1O7VYbq6FvGZh8PVR9lWPHarexnmKkn2W38Jihs1iwIiw7nPRT5N3PQLA+9LTmxRV
d4bkb3g8Du+bXSyXUir+UInZ2e7c5MteeICnFdNkof0h3l1DD3DGdJIxgkg/VKV8ZWC4fKz7mjGm
ieGR3U3hoZzFb/ZhcL5srJ6VA0skiDomb/Aayz5WTeIpTEGyun6Lbwn/rIS7eqlJXPCEDUSTloTy
iLDMXCYdEWs2PpZX/v9eqqcdANvgfurMxOssvCMTvKuPHtKAM7BByHB2o84rJtqb3s2a0ZYcoD8r
P3CMzfoxTEgFEIzL8NlsC3JCHwNiEZwNDhTt40oGnQ0Fw466J7+OMFAzid89C2kBC/8z6v0IqKHs
I6w/6RXWY7K9kqBI8gsDW4/st3EHOP4Pa7UlqVnanl6um02Ogte6tJvsJ5lWu7kCOr2w4tIEgu3k
2EXibR00kb+QD18GzT7CEyD2YNiIt+EGBezUHENywWvkfkdS9eXWbCEsX86mfjW9GTcgN3Ta3RuV
m+T7VjAtS7AZKXe7qUHG5JZbdUbqsJF7oKPUrZm/oQWxzlu4u2XUrzxDIAsuEuW1+Vixcz1REJi3
1UJgYZER30DmutDfEELHlr4DOMUUVvnNR6F2PwPIeSQDC6KgcdYLmpv1R1TICR5+zFjz/YVRy7Ac
l5ySwFCZ/dLcbChnCl8knvDOnWgKRCMP19zMAbMUM916G/rq4/Z8Jw2KyEaI543FPWNXOsYJPEfK
s8Euwe5qJpHKtYNitCytXHi+J3iw/F+3QaAFACIkIigjxBXl0+cbAEOwgqCv6JzhicqswgwromcC
BYg2tItuOPGNXl01owRH9kRfWA8szJlBUzufiud0qZuBrNNKCuxtvVdR0bs81Y90tWqCNs9xaNLQ
uIfhB5zLgInEtMhcf/VH94YwgkRSKreDh+caLOsBOEdnZg2yJ2GQtuqI6VgAknMFb2LPq0c9p1c2
Pzxd/61XFpoEyjXvfiBmSyzxqxe2Orr99VOfhFvlmka2KQbJMv/wE9nSHn/duma14sUFZnrWTbAR
d/LznL2HzemnVSfqsj0fSCd9YAUeSieW8bxirC8I9YoPmrW6a+FN+jxorFykU7x6CmFbtlPjFKfi
IoEF+UeEuZ27Yd50Wpn+iOyGZK9wAKM9SqR17HDA8EWd5jEZtBh2/IoYdLyjmy66bjrs+MhbbZTH
i9fz9WYJuwE/1LzaR7PJtekx93NSO82dyYLQWB8uUakzFYXSEWpp/tOLC7Mm1EA8UHJx5dY+fvIl
TVyAyH2FWNMRr2x2zG0pZHqv7JnhR7AEhhwPr6mYj198fLwloqMW/nYOjQAoPwUc3BHfntrxQDmS
dADnBMQyaaXZ2GCzPjqhQQKTdFRPEJIq+1ZftFtxX+MJ1YRrAb0OtYs5Oamz7J7fn0cnNKB1sMrC
TOfap3lAJUn0j49fB3vm2yoYadYPgcXVeHPPAeAXLYrluAgcx0ne0hY9hUydpRUSryMtTjrTyk78
hoTrcyKOvFuyrZOT5w3HnuqxzGUbBdSW2UeM4Rmq3m3IFFhV4hgFZCjwdEK7zrDhgyTbYUCJcv/o
ZNf0trUpyxjZTq47jfssr0S1HVwJKuVehNzyOfJd/t+i6YrA8i9SgPqaYRYuXx1lSERr40qoiFfZ
6kETI5FFQvmSoiLKON97PwVYLhnLdcm3+X7bt5FPV9D/tmPup13mNY0kfmm61U4Fv6xc6pG8h8/b
0te+svJ3qimdo3AKGkgBneGUaIygGRySCi3Lop5fO0UW3fKp7uBaLrVA02Pa0Y90IGj9y2v8xQ/g
Vu/SQjcYid4sxktsVePbvWpaKt7eZ33tBsEvvQv6ig+/oAynnMIds0KiHyIwfUSknTL917gJcl+H
DlCov06+yiv4BP09iOBdBrq8lcwn6ceK/sJV2T9QV6pBUfyh9GixyojrfWSiG7IBhBbSKOAxaWhz
DC/x+xaJsuIldF0+5uKW753ybcgZZFdhznovU5pn/FwBqkCzSbm4siHaR9KHwBtEXTVlpwC+PV7m
sgvLZL4/KfRuRGGhc8/1Lr09pO+subGX9Da+B8qtM4QrlAyX4X666OQ865dPpGBlkA5vJPscMqgF
DURH6o0S3pd+W+xMRb+uuw7Qhn82jQIwwe5+a1ITBlWH2u/gjN2RRLvjjCNXTx7xAiU3juLMrS3I
dHril1Kbh5DaAjV8sNud7fiZn2aAav9FmWGL+DLXL8FEymNt0YDDwEkG6wQ32cGnX+mKtnfjWyzC
GooOLNIDMHbCp1rnZv9CPNC7Tp5ZsehpkoVnBFKpMxYT2Od/NA5BPSX5beI2arPKvvY16hKuDbhb
7QqeD2fKAzSBvosiOp8zt4+2iC3GPBWiVciBEtujM6KQA22KKIuZmYmV3s5xj10ER0l244cZnoHn
MeFMG1NiO5PBZvwnsRsAuL/pXFZgz7/6u7/4Zaai5sQ32vyDRCeQ5xsVNp14vcyNl8nBqnzrwZKX
LCsCX/dsLFFlx0wol9/86o5sKxCmN2nNbti6q5QhABcuierOclD31FwHwHtsjOc5ezDZy6TcK3bn
a688q+c1CnhJA2b+vQ6iIGOPpTKplZ5jiSJclrElWQSTLLWu1SUjik6CA/WehIM3UgBJWAyZb/uy
zqMDqcckPh/+3asaSCc8nE+me6GD/isDmwt31hMkSwyW3TYKU3dFjuSQ3CgoJtGjyY6x8AAiWsnb
QzSsdk9bRIiNMRGXVrT0n5Meb7as8C8j8uZps8/Yu1LhEFZfH3jyLC/84OBXmbmzDt3f3lVVBqPu
Abbguy2mzfOGau/aMYIdpaNg3tu7KqmukE7w9alZt43GNJ6R6ngPzdpAr4er7v9GaEmDTFbj2GQZ
Zkg8xYVj7jLoo1cstuNy9bM75ux+RKThUqe6hGzcQFS6mVSvjrx8u4rHKk/G98JZiJizmhdGZEP3
jumc/aqDuf9DGL3TIC+dISUcNTwzU3X7agb9gz1dULoR2k6wIkZBUe/l2N9bhxrrTEALff89TIPD
cnD5tv2lnAXALisN9r4wXpcZ0L2BKadjzkTGUdeqYoiLSYVt/Z4PFWVWn/chTN6/kECl5TGqFYgG
JQ5OvmX7Ds5PBqRYxlsUkuHlSxBPPd3CI+WAIL4cD4L2WrzfCgC0MKy099/dLwHUpqB3rpnbaK2U
SJDoa319oyTWSNhxtKeM7hbAXSOv4s+0RJOtLoOSI41bcYEG0ROaV8F2NC45K9CsCDCO7vQmKHeL
uBGW7oYTTpdNxX5plmA48b/XU8QLb3VeO4xf2p3BOHaYp7AxoUIWHCySXGBBW3LTp+nz+YyalFvs
HQcH2/j4jr+rVUPP+EKbOag8m0QUzfC6AfxchcGdAbHtu/an2UUvuoK/ZuyuRgbnn22QEf0eL5wH
q16OUFwA+YLviKW/Bb0ixsQs2fsTQuzXYgtQYZAIbgyRCtOd+1/Qi5splARjV+Q5567vod/CGvFZ
mRqmDkjBHhnz1C9nNRzM1RvpxHLwLkfgYfXWeOkshDgyWhrfd/yIJPGpQ1RYXSeMi1E8tbDSQkpx
cRAV0+yOR/CLYkHCiWyUrv7+Xm9xJclM0Mc+N211WQNwOkWMfVvJL4aidUyFQHs2nPi0zC60Dw+8
k/LfzRv7vstVoIHWIKLNBwbK4+9tPGbtihfLIvJ1YBqv3JZEKSGOReAm+kyk+UWFgOb17uRq67d9
d1xcI6WH6vCfoYdU9vdX9GDInqJHndZKwegjUkK/V1roWBUXVCO4u+e/EbGQzgqASrVhoCqEXeOR
jltXMflrskB+aey165fO/DgPjboi/l6Vw9bMg9IEoKGtzx71dSscw4u86oqtDKkAOI5jHpJq2FVq
rOwEPy10RX5KGHJGpCRJFW/WRVN2s45B9Vp7KMksUPuEdI4XIqhz9rervnc24WvaW4Xg//vCFoQc
RcEKDoQQGAUszNib0Xjt5+1EwOCxm9kdKirz3qsG0ryegUGo0MKR26hCQnsxfoqlWqupQ2UVEYLX
QxYzgOHxbS8HvOYIAfhEEdS3OSglWFq+T6zVNglwAPTstlXflqw6enxwt9X2NqwcxrlYTT5RT2XL
r+rJepAbW9M1dfvUQg3SSYh93Gl+Q54Rd88iDlCD98Vi6qQ1u3bT16+0X297tOklwBZ0x/b7HS6N
aGpqAWjuiALQ2SSTl53gh6LvUCvKK/ITdOG7L/5eW7ImPkDRsfY45S4u8fqgzGV2Cu2o7iQZU8o/
4LQY3wiRuh8JrlpxL9BUU+9q0FQ8ZIdTwYw3/OzBZ43bJVeAwGBO+YBsGik1hV+w0wwlA3RmOxkO
byKPZK+tCpZaXf9Zk/zPzMZ63d68yXVF41yijRqypEAdUfumvNcBUngpXoH3rwb0szyHY38bEOnR
q7mnmbnyE28dGgQXTs5XnFJkEHohc04SW99M8qKed6CqeJYMZ8POuiOce/DA0v2d5tniJOYwqA/W
jRItkEqdJVPoDsfnJIdYrqvJe6bo3pq5vxLGUPmIrg8+jtv7UgkFcpHE6ayMibEj5akLzjQhgcaa
udsPZ8ZW6955g7OYSrWwmJbRFOciaefuzaQCSEizf0lpv+D5ypUDBWc1N7R4WMYtJ+M8UIwV2KcX
DHQ9aUaq4NyFS00PYQ3t+pnioGs4XD1Gj9bBg4te2QutH7VcyoJdKJDhMtaadO0KkBvzgHYL6AQK
MRhP4jIknmH0yhvXj1gYROON7nTbmo53XpT877jW1XxPHn/yDeC569IKMZfrlJ0fj83uTB9r2cVt
68XaheP6CkGEYkPoayTSUjpZXceHc3xQwxfAcMzLIaB7EFfbLRZ7/xJthTRMgWU/GtK56+xd2B9d
ZbTFUOe09Ut80BGQk4jMJ56qPHQRx/FbIhjyn3PD7zs7jZ4lXAfB4X4bGi70mSdoDJJrIlekstr6
Fn8gfjGoNHakiAime7AuE2o7X6YImU0qn79LqUxU5/mI2MEsottABbVFJhKC4GJn3LDJ5RjacY/+
k1u8DUV4BympC67RLPhdUjTNTnbmN4Y+118Sb4PWnsbz21tlP/KvJlttUZgFW4oirHkcbNlP1ELi
0vNuaEOt2D1K01Sv/hL05qGv0zBAT3ayDkbWdMZilcT++KUmG0L3Y9AhFN5msJ58a7DbH7gkTpJN
BG5LIIBwr9U/dl/nzKfQpqD5yqZNeB0Z8f9zWnLYbolcp9RGRH1IOthteG9/7dGiEC+u0PxhAevO
agz2epHpY1RnDWW89NtkL0uFSQ/ALXyeMOGfV9RVY2P2kR2a/bK0xLHWcUi/nyoIF7V7hAa8mh9T
O8vELpZhCWF9+7QriswSfYGi+iGHZqyZSe3wHH0DrCNq6vLOkN29CZPU3ZCvBOldM8Npyre4QRKi
w/Gl/HwFOBFDoiGF9VT07eLrovCsQOLVKlRRUNLl/iuqZGiGur/h1ZM3EhRl6w1KqOdiZHG91AlI
XLGsOeIfCoMJkTlo3gQyXIUiDi0TF50Av8G+qQp0C1Sg0tS2EsdG8u4BcFhbU/hn2mUVLj6+IFZl
/iHgzJmMTl79nbs6JR6ffFe8vxL/jNT652q1SA1hbHAX1KixVLjiIRXTSZtEyLibNpT7eggdLxev
+UOcpFbpoDc0cXHBcpJ7+0dRqsX15dC/FBIE1OHiS6X5eOLNmoVgC9RreESyvyWZE+IwbXPcZrBf
arOcQptiqpG203DiqTPpgpmdnyDdBtVMu5vCWolHfAljksffnTsvg4Ub/c+po9z+yhjyXZShqrhC
05qiQmYwwokF6subzhYz58X2Oj6L1rPeGI6g+jHbJh48+HZ5boiwSYnbdPV95Keh2k8iynh7G2qy
VOXI6MZChjsHiQuP/4bKKVzuMA6pSOttRXrA8jb7UF6r6z3O4LCodCnxWcibzZZUzxCWdZRmK3sZ
6SwUTdCsYQZXZSsknITIuYYow81JeUEEdwGywtdQCRw7pOg8LeTkkhbrcEfMLxFuBASBBvLNqD6g
Ls2ogcEe7L2QkeOfBCTdMnjTBvh6moJyvPV/5vRmYa2TtYZ34ZuvGGfUWmLR6BEVzRhrUaTZqQ/V
lyspEda3Nl8AEN9eHDtLHKuBNBCx0Avzhko9aUnG6pCS0JtfcjRe5I6cX09SqIDm5xz2Pyq9hGQq
Hd0t2fpkAy0nGlMt3KS9geZ7pyCqP58wzkj/JlOHUxAxhH8J6RLMCSIvoL5tIImawRKZjEUGBAqW
+t3/DQBkkK8+1NKc8w3R3H9d8cRGoiMONGwgOi4F5+v3Ics3/Q87Eursr1ZQPYgMgkJXJ5wh4Hl1
x0eqPNXJXGektRTOIww1M0whGRI/vWKJMWXiiQXiKkKrgpfKDhprDNc6YBLhQjVVexdyqIHN8ThG
GMrlFt/DAsp7K6DFK7NMHWy66bmGI6GBnzwIEwI44c2LXhZGG035D263Pv/bs6nlyoV3w7hd/p1/
a8PYawkkZnc1FxSJCjt2GIy/snJdcmae+8EXoAqcnWnvPdO+WH7Fw/EqEXi5FD5GprBNHfJTmdJj
QEFFUY8ssHvfbUDWiF1md8V2Tk9itIWE7GGwnCfHzs9S01U3b2VOWhWO2WPFGh+jxwNlqVud/Q/x
KY9kUQqZMd48WYrsfZi4aC03laAmtxXMWUKdP7abZnyO0rIobF+oF7849fbCN4zGXQRG11vZorlV
ir/Ip6VgT6PlLQKkLR0P9zbOMCS7a0qTn7zhglpy3ggDeujzmmuMEpsS2I+0/EyC016yyC/biU1i
OYxwcINK97P4ir7OM3HmU88yzPz7VboFExpRb3dVJTO9bgoy4xwAuf/riARux8rl8QViu3qLL4OZ
BpKZmNzVswA0egnFhoQHMu4/mpm5NTnm2mgH/PZEfAF+vVgIbwHjARsrkPAIaKYEl+5caw3J4Oc7
h4IQx13qwgsBtQAh0Bt0QNS1j1eCW6NXectsZCkM8sHsrrcNLXK15F0Y77nLDoa8GeKfjdGsNNvz
uCGzwduCkqxg7VVdLyh3LPu6COr1f2dzuc8i9vpRZyJ1iuqoS64/VTbzCWqV47O7RPEzifs50C/F
/tKLhvJ2Z51ptilsz2HGyZLk2afRAV0useeTP2Wr5QfrxpR5i3lagcDU0nCQHMnilnFim7RHI4MM
T/qwpxijsg/CWzMt6eg5unQ7ORXTNexMrPXixhw+dDZDRek7Cp3nMJ3OsYMchieTbsi1Q27jepIJ
PTKrKgJfmRhYCGq7yrZYNHgweZWpyAC21VMBZBu4AU3tqJRjvgdlwV8+irECPZ5NQUqtz16gEnGT
yB9TqROKtD29uhdRpVC+7jt4mrrcPstZoXrRqh3oRtXizh5C0pRmnOEmlWGoaHVWXec6HmVghcoX
6r7yqaN6YnJYhXLE8wpvsBHDmKvrqUciuk2jTWwxC0wUYesGV6wkwAHYEveOueYHdGedSJRMeyOD
f2DjMwWnyivawGJ4NU4MCaPyhNGdhbrJQ+Hp6H3FBY61Ucg1xpa984YbXNegHkpYQmkYOhYqBvK2
/T4mpPWI71cGy7CeIy5dtnbg87bx9Fc9ol5YWTmBqVJYMVEjLY6lIFHgH6hwjBpTgBUUW6X/XSt6
HqWgqegqf0KctzxDxAs9dC4O6rdOGRqvvRDpbXsrDArPF8U/w/WOhM7UdStfppmxIEYTkibV46/9
Ey/Fs+tR1MJMBreK+EMXLSDfM7b3BE56XagmZKkA40IkC0Tfy/rkfKGOxlEfG7O9HE210ZUJMog1
pfwh6R9mgJq6HsSJiRS21vn75WnYCqDllotVINAHTwFcQF3i0K9rt0mvlHaLvqlY7qFl3b6d57M+
daF2dIMv4UH/AC0Q1jK6cnB8nqGHrFv2y9ODd6orFpOgZq88aMUH6jwzaoXPXqSMrb4fOxMecz+w
rVDehLVT6tdoqIX24hPeblHOCv6IC9O/sfmA66WvWeuecRFeUx9OyW1xhUirKC0SuGz2ADjwKi5p
v+NQGvAB+bUs2PMqyjWjdGgXi+OHsErdnmvAFk3Ep3ULGTa8b4M+oMj4Ap7+tw0HiayRVlqm9MbB
4S1E2jiWAhKMUsMkeWc5LW5UJxi1wdcwLvinLJp0ZyMMY9AKyeL9n4unCvIQ89JnMcV6/5Gx0oEu
k0X5T0+xu0VmrQEUk3RxTRQJc+fEsDPjACBIqUhwBhvfYbAcLCxj/z7uIzF0cRGyP7VAfZaf9XU1
LrfvxdrvVuUuWQNxJVaVrUoSvYf1WJchiGa1Pf4trMfAVWe2H7GAA49y/pDZUU3f51MFY1XC25ve
S/X7C/69E3LavVF/bO/NJ/w9jVIbDdD4wHN6haNmvLS9S10eTCjorF54qY+YK33rVEWjquR0/igU
NI1RHCi9uz/vVM7aoDbsfoAL8BZFUuyWLsO9/f5YCaxznIs070Ucp/Xs3WEHR6CRjYGTbq2QP6ND
9P3E6hurWHWq4bDSsC5mFs0zhEh4sbbuF9yxy2ErX8kivzZAiP1AmPbe6iChjZsShIOYrdTFdjqc
gNQwVX3JYjS3qZ9HgoiQA3tU9FIFxRCw/YjYrL6WAH9IXzMiceWvxOcSV6A0xp8759IAt3dNEACi
DC17czZ2vjYEXWoWWxY4HxF7igcJPiisl0mZkltdV3Liqe1aWr9wZYZK+VTRVnVR1FWUYvhMIPaI
gi4P/o13imvq5eoPxFZ/tq7mcMEJx/qqfEqA9k915J3jD+ALumVk6ua6wkQfqWLr/HEdMjpdN39U
M+t4ViGK0Q41VFUdAXJFhREwpKvcg2B/1oGKRR8qKru9xW3md/hBRrbAMppD7sI0XB7dLXD3wn0U
HhQDyZNHn/CkiNnQrbSXONebn/u8kxQ6yzFjZ9kVA5eZbZsuUj4bF6cssYNtj6zNgkyrsOP98PUN
OdytWWL8zRMDXtQewyBP8NLdul+6COxgDFurWw+FmldAFKjIvAei0mbfKneFDUa/UOafTgsBx3Qs
WUtelhYEudxXNlYfg9jWgQdpP3CGiXt+da2rbV2r/UsQ3nf/rUC4/aPcCO2NM85/4jHN8CuLXUmi
8Z56t/wKJpRfYJXvLk+bqX87amOEI3AFbjXKwtk47lAGd+sXDZs7iBLq3iJRlP4RDCo9Mxk4Oily
7MmKFP8rbJBSlr9ol9aIvpcuoeHKLxclzvEXHvOEPhMj0UkAJ7KclFjMwV+uvTrY26I5BANZr+ZO
NCdB06v5RVHSzTknFogKMF1psKE9kfd3bDLGny8XxWuveRTxldW95GC6fW8fgyOpnx0SxMlf1Mbd
BTp+OfwTD4vx8NiqhFiCYqG84AzyGmq7Vp7GDkmdwfw+jqJhlq1ptvJp0geQaiwbOHPSPYqp+Gv+
KKjYdHAXaciOpBDWfdsuO/Mj7WtGm7EuZiv0Lu1VhkFKwPdrE95mHk55T8y3ISQu6PsERHWJstwd
w9ghXrigYYJO9zbE6UoJ6KdI8qMorSiZ6W1MYdtYhdywspQaHyWR2Zo7N499dQ5F+6XAaEvayC1A
EWdcuG4LvGBV5mZK6sdS/SWgJqOTR9K7gdugCAn/fVjmd7FvmfwBs8XNM4yfTYDl025OjFg7rRhq
G8Xa5MgGjFYNxb0AYHgis6JvXeNWN4OaL32Tec63GDg6P4nVBvURvb82JVM9fCtS2PdIc4/28OB+
lAXO6+uVwQWGPE0zRNw2m76mq8NRirJrma9n4/9/SmsuhlOX9WmeuwTCzdhu86aFkli/OmvzjT1G
PQ8CO3LSBW7nRz84/D8wigQQqHMOnug/TLf+CbIKXlc6RdN3hQP4wBfY35VGha1emM3LUTWuUeNC
6AfzYdK9XS1cvR7t5Q4affFxwxeRCdbqjqt0UhOD3L6s4b3AB9Jexwo5ZjfQDxAu9PA/1D8SHmTW
v2IlX5WhAWikJHWVJRw9Tv1SsAvabUFHLrNTa2Gu7J7NezBNogUnbZpXy88uSFB3Jf9BiwzwRw05
qBOC+PuSpPUj5OXhTzAOOLsq8b/wLpddZRHWBQOCfeR7LiMj6m7xT4oMQeNuymISxMQzgPdfXoWH
qMoHNI+kInG16btAxpn33aq3o6DRkC9P+XmmEwXTgp90ZhQop/Xldh0b//DF0xB6thsdkr5YPkpk
ZvJ/2Z4TOyuAalzohucYOD7gf+eN/iI0cVZSqSB+Sl/SrJsclzLQObZlvln4LPiVV7Bc2coFFWUc
/jYbjReyEHN4OcKEH0AAbhHF5oxCBBNNZqTx6CauAUon3bI3CmemVnz0KTeasLJzP8uf57GqnkUk
NIMFatbtMB7Djzof3ETV+JNklccKPqTG9JAF4PRIfGsaPUdN1iV9wVhUl1fyCIeanfvb+Q+d/gH0
mtf/q8ridtZIMXQw+EXMemaZ57hLU+RaEjw7kRPbyhQixiEFb3yyfV0vXSZ9c1JS3BUlCn14hqol
/XmJO72lcJep4ktfcLI6UB+Nkulnp5wRTmQqLkafGrVAt2GR38GQQJ2MaYNfHIuZF1A/1xqtahn5
ezFOkr9ScD7kjOuDkwHLUoaQEMWFeeKhs57QLBrJ69UNyYus+Z295Z1tKqm0897oOkmAFTc8tVUj
8jFkq/cr4caAvIbPltqypzEvptXtmUXl99F4JVeFkvecj6mOBk6ArDXbsk1nl9BNHFonx+hAgCSy
XasCOJs+I8jcDeeAhcazP83WW/+EXdejo7GJv6Ru9dVT+DS9a0gKQbB9dNa4PjC93XDcp+5vKV/J
HBXeDFzHLiCv0hDJUCJHJaajigYazLq2ob5JJsdJHdhNANneSwShO+qIsVMepSNoTHVNRBDuenon
G7idKC2qLxF/6dseMtvxpRjkiF2zqrJ59furk0NDjcEq/Qfs53ItL27N8XM768dn2Sq6s82V/Ejx
EMzO4V6swTJXCPSFjP2mSyNK/g8BO9OVS7S0p/srA1C1J4MPzOTlThgBZMgmEn81znBpf8Zv6rLB
4z4aW3KSlV7DdAotsMIhLGQb211W0H+NKQmWMRK9fxqo8M26kDZ/GqzpLn7x4THlBrZjCDZ+VaUX
NrxCXf7rGPIQryHqMm2Laq18NQp0VQuj8Wc93CSXsTWzKru8il2Skr1aHj4ORtwnGKRgpgbJOgaj
jrAKBL7X6ju8JP8zxFuIarfm/rJCsH4+5V8evvtxM77Q+xvy3MDoD+W4ga5omGU/k/uZ65Vqfiud
2FNSQ08gGtdJ/K3fzUWPB+cZdG+TiZA3/QAa9bKjeaXwcC50M/4vgVJMiZ8bvP8LOZJ9v+T5298S
sx35MPR2dlJvx5ccKGS0WjY8ydJuIbO9gB+IvEb+BNKrodECXB/XFwGbVUvTS/PGLw/uPkxx23Wu
V/RXJBpxlpenfyXo9RwT5kMVcaUvDGf6d2Xiq/fyGb3LhVR9cb+LbQjgTXUXi2rb0tY4BmNSt6oK
6tzogaCKpPO1lfjeywNZDZ3nKMEwG3LdgAm/PtjHq1NlHBTYohcfKl34hsM8F5atkXe3LtXUBI4N
osixuVFNud8RYkhaXCF6y+Rgb189JarkwoAvfPGZqUc5mjQpeMJKEwoC/SkTncrCFuiqRRXZ7HqV
H9igJQGNJqU0bN+p0syfydK2TxAQyxXB6BhjoLmp+U46beCiPsCEbPek5+cfknwQLfEYpVR+Dk2b
cWq87ptAhtAHEqAvyePbGwpRDIzBXX2UbTQkDvtfdWxIjK8nkA01UVWxiABxAJubRpJvox7/M9IZ
1Y8oTpTM0HPSY0ANvLm89/H6BJ97Uczyn8C98tPT41gHoGQmVNAX/1uka6wlPrQml5/LrSYie1XJ
wi0H90z+bOB4jzGo7yg+z0yzv1D22oSIH9FNZ+R1k7gNLKphHxfr3u5eZETh7Y6c/10qQlwuA0Yn
BO2V6I1wK+3zvG7noGJilSXWbTftkCjvPW6qqPpuScvDS+OlTz/+cbDjVD8U5D7NlOJF7cluRI63
o4zNSdyKQhLNMFSo5AN9rdunyp/1UVdYbEx9jtvUouMtdAbsw/qb5vA8732JjgumfhndrotTDwIR
Y1s71lEiO0KD65Uj/8Gdm731tqgX5l6k5Sq63NNMuMLfxppTFqn7VjFBcn8RVKq/AQdLpUsXBRi4
oj45gpCLaeET/nvtfTRtbb6Wv5RVPBPuUdjUtzfAXsUarEoeL3e6mypzY6bkDqgXBHph2NTZepUS
NcJXlSmWWvvn255Tp9vVV2MZsAL1Ptkt8MofKEnvtAza+tXkGCYqh1427lZWj3IfMi4kB9YClDRP
tztmfV8iHo8KsjlUphSE3/px41rmuiGMzcUZFDnTkUsKx7ZtZz085X4DeuIwJXEuYujOZJeA6cwR
0Nsr3a64BBWCW6QzjHsQ6g7dZttLgrUHJ2SkxRkQsb9kxiNw5AOaBENuOhlg9LHHN8k5w0ow9uz1
j9+L+W3sYhl+pNjvO1cSwxpdi3DRmXukgPEGF45x95ryfM92Dk+x+MRiBzh3ZqS1d/hcP/mVf6yY
35KMPs8PQ6Z92L+qWuFfX7yycpiiE69AjSms5G9aT3DtY2MKNdtrD/qa2Y5bKrrULSV6p4whRWbk
X+sHoq3gAS3LumZ/dKOT8Iy3PZRN1WwGAtwIWD+hFz81BHejlTQGa8egs4vfh0dn5rO/3VAIgYqR
vnogfqsL8/nkaV81BxLJYPNBdmAk6ROCUi/quLXB0jJLDNvsLV9jRcrvrjerL2CK/T4PRsFYJi+I
KteXpkD13UcLf3SFRZQXcOSg4h4DjR6qeVNoOJLxe1z/VhfBhMOoI4OdoTIssbtVl5M3GuumsclN
uLuNzAKRxnoffmu5IxbEf9HuZZm4DU51xmKthajuaAwSF1QwvzM1ygVxGIhBzOaGE5rhZZAELOkG
wKLK1Xsl/MfKrrUY+5ZoFO1LeB5sFpERKMY4d0oMPaO36eNgaerZeeGdQuVNORTgJ85Y3xysG7fZ
d0GynJQkf4J+UwFyLI1inrPVve1sOiQ2d8PwkJHS4uPCeuc1WhnnO2/mhJfl8YamFEQYoc6Mz+vW
jBfazk8gc7m3fsOgSw8LobhBwmDqvfFhKnwJdDBBs+eoE/uvcvnKZeIbxS9Xjc61sCQ09cq6Ybbu
dSe0k4+16JUwB3Uq/LkhxfLx1vyUTvEJ29C3ir0lE3QCvGR3T/wH/R47Ma5rkVlGV7g3fDxK29aB
Y6JXLzarE6v8LSHT/gMM0MHqZMHCL2YzDaSB6OMQo4Ley+uRstQ8lDdgu4ob7t8XlgVvcvqZ0RNJ
taemus7vTnrQ/GAoT71JEB3ivEJ0YTZnOnDA6nv2fekhL7H33Vs8b569nWs+z6MzcT7f7HKvjOf4
PtJSlC5i2tw1dcMldqJw0ZWaG46V7t1bZuUfQ7/9QIU+gpDrOPAmrO6+J74z6UK9WJzrxXWVEZzw
cgtT81pIdC0w1z+VvuqtVWg0owjhRuFwAdyFt3KvxHC2gFE4mbh6BuHAapCcGPlTXpJt8XmipHFd
CQN/9DwTlMdLA6nmQNkgpDNabpsxgnlEky7pjTMsPqmo/TzgR6e5b84ij7HB4JRHh8FW0sdIujzV
AfN526CM758InHmn4Uphokj5JaAAszd/U4o0lfzWU+vNQKEvf1sl7OmVb+4tVYE9AGlCKtZt+GVj
Xkz9J3SnOf0v4tsadK4/MQKr4rFTmgYmXnP9DD+9OqOnYqlLC2M3F0zAKCarNtD5Pql6TqB1I/zo
r65rORzlfan7rtuvkh6gNrHzs9+R9lONNgQfje2GckSxQamN9SgzWlVOCQVb8aygmd2eEBT6wGd3
Ve3pOnqlsFPsB03Qwx5vaRXxJ6bt53VMrU5gi2h9JOmcS/wLEVUSkdG4KwWJpP1GThckbAPEWm1w
lNhtH9jMxVmdtYZ8sz/ImbTn+ijkuVmPm6mpEW18JGRgHM7+Ad7og1USPXYZUrn/qZRyw3OAxnLl
fnBmpRY5Wweadbx3qDbVwvPtE7gWegl3Z+eLPjz+8yIFoe2PWWj2cr+uEru/X7BPLTR9XfiBMJ4t
mBi5IVlefKDwLG01RuGfL035AMsW7//+/Yvgn72T9d3Lk0+hmCegyIKalm5i16/mvpzLOIFnSji0
LU8PzigW+jmJb+eUBQ4vEzo1Zw5xnNqniT7oWwDnM85FgwSSTDZcOfse2RTCLN7c5MpCaGwQVG3S
+cAvU+8u+QwxiFVuSy9QyecIRcNQeQQUd7gJtwrqGuWB2v+tdLq6bnwxcoBUjRpNlJyOGIGvyDBk
bbFTA1DtaFVA+4TpkxekBx9qr6voMusMWpgmDqJ7965V47ay++C+ofoDzX9eRk0mzM9KihfyFC5h
U4GfL2axRYL4XwFv5rFL9BFwOyhmdTvEBZe5NNQxwdRYICNyjxje7hWg1/SSp9Fo2I4g8zMK7KPv
Qp/l/Ez7qRqxm1OpPIKksj23G6ss10gOZqpO3uah8FvvBLF3Ljs9Zd/n2dLLoMQPzt25WWnf3wQK
lCSnHn7m5a77crrF7KrkE06W1BvVcz/wDBoxibw1MEIfpwMzA3CHg+yYih4bS9uYQXbMm3jWxAj8
nuH/+La4vDLJPGZ4UZD5h/IwclnIOuZNyLb3Zgc2ImsCx+1sDTCKYbWlUp4LAwmdkAz8cUxdBbTi
sQ3FGT5M/jalsnzD5eNFgSJYDlva8j6yGqBBNRGqo2yvaopPSFM1x0f8mRg7habPI1HOxJw5AoVc
rLgkFUHWegZGB6wOGBoP4gGTEBFCTx6afwKVgN+WogVM7JQ+u0ykzublm1cmN1g/OcEss+RaMHyN
mGM/MShAt3a0GVGW5F0N05Wn25BJy7v6FqHDEJrVMFR7kJDR1TyV+yG0+1pgrmjbqC4owHl1uw9s
o1g3FfEJhxkay8gt+GloPclsLXLtGGmxdpC4tI8N5NEIW6SMpK8LwO0D9xS8H8JQB1AavNlaRwCb
4EtX+ZrYUkc4qXkrhLBnLUk9M8c/+5Djdfx/jdttarIttCKY+vMtYLCD3g8bSq/95Yt4ERRbSjcV
3GwSFRS3jPxc9gF5TcbgEmNz4Emp3FHaMSN+4Y95+TYahWLZPiYbZpseGWf+5jGGeUw48Wl7MRPQ
/QQjO6RQZibmFtuMtFWw/DnNpTHy47k4YV8Vu91KIDLs/dgjVHQdEBOkyt1o298K/4kCiWo5gQ7U
cbB/2qFRQCMV1Z7Aq1RT+dJjTSoJ7+u56OYtd3QPzUrZxws4YbvuRuLouz8ZUI1xMXdM2q85tHp5
s5BdykrIeK+LlTFqYTZM7zaiaOx64ayUFUYqpiXuI1FtzSkts4zIUES9Ar1dHNYZTmgVmhFwPV7+
Hd+Rq6gKa4KIlgUG0w2WYMPB3zawzGwcFpjfxqEaBcxgosg6RT7uD8Pg5FDmJEzAOB3red2SOFh9
L3gWsc5jiehp6DcSkIIbKLcJh1i6krNxJGYcPQ45MY7vTY3eFOwCEQKmXzu+HSEsvpbA7CDLzO1G
8TwDjsivXatLhx+L9pfcMrzknX/n7A/w5aUnw97hCEeuNsHFbMLpZab0VsSF+nS1ZnJ/S6g45YP8
nMOdvqkMO4bAfimnEoXqnoODj2A+7T8yrjKO53FP2Tkd2VLUQhZ2kVVbIVriPKQjXMaOR7D0HB1b
I18gmIzEzQwH37X/38LEqRnFvOyXmSM3eGEVe3ytQDnE7QHocR2yAtvBNwRft6GnLJOSP+/VQzGb
uHL84ztAmOO/7X1N+X6afE7CvYBzSauPrHT3Vqj0yq6j0sN2Ll9h13Ys7MB1/Yw6my1ENbp2CRES
iLLKInfjFzvv7KfkDfSzzYXOH0znYIyL9+HCG9vZfvoK41SKGpWeSveeyVD2hEvN132ney8oq742
eT8xdIxLplYCICk2RiAJA2RfjbAKAZ+yzn/2BnOsssrwWDKbicBfiaaM8PTLNvxajUjJy2/ApjAj
qh76DVMzwIVFO4IZLfEUaM7Fh0lzw+5W6WfrCB3VbfPGnJpbNDOvsnHGtmekrKoI9OI0vsN3HeNf
31SVH4kQwa8wRDPr9m6Bhps5K7f7kEnKM9spB34ssNS8qQuLpBjcp++dUK3IfJ9YpIEmMEyWUlmt
xqup0L6dqkR/pf7IBI25feHsf68qKbjf62rSaEfr7aFfv12wNAfABQ1alJdQ8UFNfi0Lq6r+uf5w
VLx2UcEumMTYu7OEov4WWWsxPWKfaFqOg75jaZzb4+FhklALNhRGMdtPradRe2/Sv3znJ+d+rS6z
ynKAptej6rzSN9PmpaU+I3Is/wrmeJJfgeqRy+OuVpTL5MBAjuAYf0XsBCkkphmmOYUoHmx/Vf0f
FstMwD7eM37CggPecZ6GZGTgvMYAzoPcraYf/0V6Jho2U9zbfLmWyDC3AssAXVtAoL/MdJCaIXwS
K3t1LeonjhZ1VE60puAcoZSUItMahF/50LYTcYaKs5OlIvmUa+q9GktpI57GZiaFv03WNJrLkF1X
LVLmi5al8bPprJpHghOPbznJhUNtWob6718ZuPuLH7oMCGT76WyUs4G9mnNt3K1BggXkLn/RmTiS
PEyKvTd3XMcqblE7jA3nof6bgf6ict7R4isw51Wd40PJgTH4NP8aUXamXP+w15eTWfNwNqWMUgpD
e3/zkLfruW3awosvz5nHi6GTzr7PuuQTUGabBxHXoXBLOMBCOdTPUw9LQICUso9SGLrioAp0ep3c
cjYDmPBQdDWp8DaR9p9m4dRyl8BPparnvwVxmPLNgeqR3Wb5AbZYVFnNzN1w63DQ3mBoApm6PCbB
HLC1c9OtPmY7UCpDrsWtkXgMZw864iCDp1znjkjDzXEvhf5kedXn3w0s+RMBgHhPk8PpZopVj+CO
VqIfWjwFVN8ywTFJSQJdVhjbR2DZVw6mNBxsf03nTEwfQ67GKMIpSDmY+GKhfqPg+7W6FJpJxHqN
mVQL5/jI727pbdAinaXJjSFWHUFURs0u0d9GAD9OHZXtV1BuxPElduIVW3fy2JIhPYEuwLSxbcAr
xbnwqXuR4SvryU7t9F9UPKuK+UPheaPTc3E6JFkG44K3ZPxX7zF5uCfl0S8O9ky9ddmUdZfQmSmr
q3BIgMbdKzqc5qOfoC7IdJrS6jSfdeRKvyAfOE47EpMF34TCf4nCK0LZBS+hJ8kwVxEpIfKk7Zwd
6BXlkeS3caBa4hUCJ1lfW8j31IChoScMXdIdYy/9+2lLB+1o/ibtRy3WG74+DkmfSLtbJ59plOb5
wGGvrX25lfreSD2DwK8g0WvD0BB5tUYrHqQkkRIsgl+tLr5wJg2N4S1ohwbEcNnmniepl5kf7cqo
vtdOy1Fc0fvxYuEA2Uj3cqCadg+eyLX9yGorAjgLJqUAYNQqcjR3r87uBTn5EQxsx3YWedIBTMVg
b4TS4qFgMIZgdZJatLbtSPK60vqFLfrOWBrpwQG+y18/IkfsRIKDip6EDVdG8fgzfU6cMQ04eN1u
Uo4XemtUanXLUNpEZOgcGXfi/CYEYK5KYzzOmmsXCGiMDSmu8J4/XzyndJa8PIly9UysKlt37C8a
eH16po91/CGLEFfZugy9BVMnR+8/G+97Tsv9ca6tXHq80SmauLkKnDma5WbaCvvR08w+kCHKKbu8
DFppDhOdgrJDpfUJ/YoL4RH8X+PxKm56LxQSbjPx6FYaT/+UmKNZPyHHfMFFINr+nJfD4QcYeSvK
1U6CJcTRYDxESGMo2IpWbcbWToq97PsmxZVFgDWa4rZyyCEtFd6MFFcr2zqMs33JNnXD4ys4gaYL
rSQL+9FjmTLy8FxUfM62A7v7yrunYMKTpi+2SrYpz9hrdIxwRGpi3zVTBWRKJuVQ6faioMNPvRxN
ahoy/WfsdUTCxeMZvgRRZ1XOGeuLFOM0N81x0dEosqpAVu/vrXUgJ2lodYumsVGExCTJHQhtosvh
O8l9+c7EZZC6gG/anMXwHqXBaPHkL59i7yzyTGE47sxqRw+6UrYzEVxnKH7Sg14VhoYs1+qLTSFi
CtKLRcLqRyKOGqFrV1QBFiPWWvVbqMukQJQznZ5/C5qzSpBsGmc4o9BurZN+bU9gN/r2Ybv0ymK3
xNvHcZRcmR2pBsNL8ldRVtcJOuDiKXQqtOO1YuybVrUvt1a7xyje+Ga0ughe43140vywALdEY/QE
idL4AtBgNa80V2y15PJ0dVnSQgA7EEFbLiSNHWXlpf+a0/X/WyhEbkzAQf/yI6vL/QyK054QbiGQ
e8lY/tR32SGWgLJW40nito37hJPx7W61rY+IANsmQtq5Cc950JPYillhT+hbUjHP6ZP6/4Yp0Tme
yAsJD+6czDNXs+wFKTlu/+S6zk+09u4eHTHb419ZuZxzduHEOCF3kyAy9oAZ3o5ElsQvi6axCGds
fEt2TVPyvUhzu/i5EpEuqZK+Kuz0IZzn52gm/cjQ6a0/OoBNMXZbmVVrcDB09pyXSs0MB6RIIW5M
S+uKMplyMKSHRtQjWEWyGFSvxb0g1ZvsW1grVwNtxkrnmImdUsOlRZ1Dc9kZRaHYIKsIsmMqLuZP
fRp63t4X8t83KRl/tEdnEsw5moP66LcMNBvXvbc+qyyUOtOPj/ufxTmbJtEyKPQVbfxwcZjDxcF3
1s7KoXo+a+09n0TEwiH2u6Iw/m4dXZU3t3BeUub/h7RQ1HQVSySLhdbZIU6ih+ywTAC+ulM4I860
e7P4e/JgTOh/dQEH7AZwUKJt5L5vIJZEh5V7i94FKMdVXQ9Hp2BZYWA8r5sUJeCT3Hl0jIrpHpqU
oF4TzTg0HC5RE6bx6gNC0b0ZUR7B70hADBUopyQSzZ80jbVas03DgiQMggfzyTFh/ZBfQoXiF3ZQ
Oy+vEQ1g+4HcKyVNTkUS3qyWGJXo2YGN0zoyHrzuqxlpb4ZhK6xY4TVCkfIZ9ivL9IvO7UKrJS2K
amfoQ7bXyNmPbEc/UASGTTYG6VsBLZmYmVeSvKgp2UjWMHexuDFVm+dWBJOZ55dZvzFEmec6bhD9
99Y39VUgZbzrugGeFTwMLX81CE7pODkEw/PaX7A9xPgaW9R7o1wwx/f6Zsy74VxFUOtHiwXcbAOv
zztUqxDwXrVtcTC6uIXdHZU3HGlYA4dwHVtGqHotsZr8oKVwz4YrqRFgUTQXNNprbcdKkZYdAbhv
yBt8GK8yqEBSP3I1QXVlZEe3SvssdDH+iH9FTniNrwRiWgn9vZSvrHF01jnks4+O8nLv3skkqKtV
fa0aA6mCS7Epoazg+3bZCsQqP5/FUqomgxFWJtz5h1JhEdXk/4xDGMljVdHxf2viXD7QhUZlthgD
WirlfZJsDAm+IoagPckJeFl+jSpzYRr+ry7YFPLD9E6Np0PqnPQtmMpvke4G83D/phFAHv+n49MW
8ogT88DzP1ot2T/Ape8o8h248dm9gYfeywPMOAg3qi2c/XJtDbrKV/aqELPF/gIoZ8fICoJNAVXc
t10duK9d0rSJLfw7M7cav/XAt2rEol9i+26guSW4W1CZTB37RS0530SsUJ/CabvMFA7blONg7N7U
Oo/fDESZkTtxeruGRORYssfeHUTu88ehp2ry2w+LOLUKNH7wsQSUvwKSImVFUiJoojGVcOO1P7ud
6lLs6DoNLPGyBab4To8ta3Tj1aVwOVrRNaDTfk+UQ9repyGbK0rZt8UaFYuFAGB1Qb9c3X9H6aqq
JiCkmkEHMuHbvBqbXmSvTzPMmnQWJjQGsFIFQ+nk270F9ZqRScEgVaRW+y7vRgUh7AkvxC/tsCYN
oHsn6FVjwPvoQGpsGGhUdQOwCPVyrC+52zazvzJmndJUAa2Ztgqdsn+BYzmN45FRx3jcnFzqnmPi
jfwAa6Z0WO0t606kzA9E32r1g6uELmvvuqFmHoYGRNDoS0XarjbKrTgZkQOnXvTwkCvwQMqOa9oL
8XJ7H1d9KycKlacUrFNJO4Ptxnv/sB5YoEy338AZXVeQeodXX743P3zmpHXHoaWSPM6fcsgSFxup
XaiPh4bDP/Rh7N7jf0wXjSco8J2b8xP6CRESom6IXfUqsuHfGKHAnjCpCDOfVyeL0xs2DJBPqhcN
b+etGY5/eG7xGXxgwtJTMN8bvpUByHuCkqPqfV2c3cOCwOYVTVT9NMYrXiX8gq5JnuR8HCpdVb7J
tIvgcZmI1WpunMeZp9eA9NzkaLVM47FmLtmshPN5aflaTw1cpkU0Ie/eF9X6mEB8Y6TnyY3eYt6o
b812851kip1WhLgVmMK5wgvv6IV9ipF/JfVkkzsz0Nodxh7XI7/5evgHpig86lvF1vJbjSuqU0/3
Byw9GWEWZP8S+dMduV3eqoUaCKe04UvlMmjMD+fkMEqJCZvtZ1mg0rNI2DpRQOcVFjki0aHHLyq8
cfMQDuNVLpX16HOo28nRI4QvmpgM1S7SU1toGN3LBr61IDI6525calJ9524vp8ElsP0cpAm/BsSs
40SK0jCoUXgRdSQF5BGPpNpu0PrrOJRMllp8T4pXWubt2J1z2j2Z9QXTZ193NLW9AFJFyyvYpVES
i6+vNiBEIW3f707bht6ImsEgtolKntiAKiJw4av76ghn0R5of/stkjjNr1CENITeanpKiPfbDbaM
I08OLUviZiy4Mo89wINe/DUivbsyOXywN8UtrCl0ECe4M2rNDQGFCQmrqZP6XwbuTgaULsgjfUxw
wrTifcfunxeyouwVjk8mVgTTHlQnH6cRoqb5xL9WYioLWccmiV6tcaHCojOdry+96L4woF4McM5Q
O7m14CGo42MoQx4OLUaUiQP9oljg7uRTwSbX6WCY/lYlzbV1BYv3+Mtx6j4dUILJ//xPaefQO+Gv
tK4feE3Z5WCBLPPrsarQiYoVcoyu1qFT/8TahabmNYnHYFQ7TfcGwcqWsaYUgbViWvCEKSK7Zxm6
Ca5XqwWr7k+nk72MjZjrFXFsjjYsBjBtsRHbgrg2KsZLx3R0sj3bT73oLFHtGWF8Ky8LBxboqI+M
EQyefjNSUkK8bpI6GaEaymVdUSAVu+/0jgVg8Ts2ZVpQW2zcZb/GMC79BRkno1k2LtHL2qwR58vj
9gPUgtyHF+4noWoe5ZXIHx+ceCxfCaz3bkmXQdtedGJj2+eh6zIYaohCIT6ulmlHSAGgypplh8cM
2PUNN6kmUkM6xIaXkHGos1OPyuOiHZaZ+Yh4k4wpfjE0vcLqzmH0SqhSxxwhmUP//I+hJ/Gi9ZTC
zV2RAxCFu7MprbLU7HZAtetBAEKMtmRye0uj20qhCUOg8m1pGqTRQ5iCgCmpTCEIir0K91li3DyC
CAd37O7+E+0nk1SaYOjn9sCYK7lmRs8S6g+soOQBMKPYCkv0JH5w9PmQTObT+DszoJ046Hqy/CKc
g7e3FoTqL3GSUbAlXW/paKKsufi79rlqRgInH7yWINjc5sezKZvSzPoGW9NoqxmH8ElC3ZxiplZc
YgSXsl5EK5YJNYXYROJFplU2clfOmgz9YskOx9sOh/CTLpRcDcQZK3ja19HqZ0ntuB+lz16Af6q4
kuxxYl09tIcFpdOCC2tX9hmMaVU2qFcD5O74CEfmOvB5/Fm1NgRgQT7Z/VutsVzRFtvhGC7A3Ahq
RZq3+lSC4dSbJZmz+DGIRVwxCdjajyx2YzhKCj28tA/YNzxIGCTuqx3a0H3iyTQKpAo8KS8TsTb7
LvPsvc3La7m5w2HKtuhxvT9gZnRYKRGE20PA5TuYN4KLhOmAPvE1+qLHGqqO3afN9roeS0dyiEDt
Ch2uGqgyQfYJtXe8pzbbo13fvLjwdsq6JhN4fPzOqTbhzIl3pA0HzlLXA25wy0NU8+iED9wkkitU
/8a+jTmhsrRfmZZgouTqOnSgirULzQeDph6AQdZSOtVih0R75rq/2LnEAt09VY7KTC5fcJ+z4ffq
NvzvvnbWXbInMIjBDc/qgwsyQGXm+GNKzf2z0Cr8aOueKLn4Wt4GmbMfASK3UVtj9KP82aXvUYzD
AlNbmJPNXcYzaDWb0sdGNGk/V6KgEyJpKSUzNggvMJdceNdj/TP39Ld4yK5wrKDjRyivkMGnBbFz
+NFY7HMB8gzjzAj0XSZFsU8MSBOj0hn/Tsd/ykyHTJYchd9pcgxCJ9j21n6i3+bKIPOlwiw/gG0C
e9cDarP+UVE8JwQcDkJwmKx2Sc0nKyCWgmx8eXrA7u62BHJ87pAu9X8hsMPEYbYr+hqK0Q00dpae
mhUIdysYxw3btjZBDWB5OUGZeTJxPobPsVyOWmZn8audh7cXFM0CqNs4EyuExXf+HJPFOWW+2dDT
hufy/G+x4/BLD7AlJmb/JGWxAmRAZQwDYNRZthTjBDULIw1PnjJhq6jztWAo0VeE+8vxe8oq2+qL
QTV7XP8PU/P7clNIO4MLpvYCACs+z2ruBSGdnYYSxrTQM9/nmC++YVCNaWDfAJTlfpH5XnAoaSTB
b+36sq9i+XFN5UKpSt08lvLhA5Irl/vlzhz6YELiIzsdb98qiJCSoNM3RAhqTEcSuuo9CzCUUJG6
XcHFcgbbdC71lOGrDUPdkbMi9RP4SLzBqlugaJf7Cl0TVxisnVzDmr2BTDfbU7MWRYis80Ch9mBs
ZOkBmHF8/sWj5hq2z9RHz2pXqNN905ejqE11JSdi/nIEtt0V9M6kyyBqa9QUm7+oAIBmvEVdrpkB
F4MYwLJqsLEJJMz5rG7xpvwgtjoTyxzyzzzkrpkGnnpHOwhkG2gyV08KtEZuil4Ejz3HHllGf3h+
nnx7Lo46keqPrJn5Gyv0Yjt3SSO9s/UBFEIAbZWsHUFcpgaji9TEZU2JC0IunmT8aBhAdL1aC28R
4UDu3+vRuzOTAnY6otyyRoq0XgPnUe7XDA3JISHVrUUo85cCA74uHOCob2VH5hGJvUJP4XrXUpZX
83J9NBiWGrOY8oJd0C+wnmRgpgnNnnqbkCerNbGz4Sjy0n4Nh2p0XVmjetn6yT7m+xqhNM2OxUUH
DojKle95g49Vnor5HEiDD0DiCPaq58oaF5GOVGian78/C5p3L3Gl2mPXaWhRbtj92Q3rhzN3DTfV
CwBWHTIVsZzRHjM3pJwnZ+N5VBdlPQ+iIFPRiPfMfPpeesa3dG1GPpB4Ri9b7Y/+VEOR48Zdt24a
y3+FfUksLkiEQFQOmEy3EoFMU5Kme6fbObUjY33I/pMmnk/TM7zkUNp6QEoNbbAt7b6Lrph7+ZsI
mdtOilp71hxnemriRfPZ91L4W39669XeSsmQlWw0uluUmGHyC68DxxRjqzPWrPEAguBLX/e3l8Lu
1WsgPvroBfdYd5IuimRJAyh0lpGs4E4sAhrWn+WYD3oxcYvWdysh9JdyhL27ZgvttOOG3HLWRsWZ
MKQaZNQf8rxwJ0rkoxIjLv6PryOGLgm9zBa7koMKGsNoS3edtbSBJ+hJqC5SfemDjuHA528j+5vl
+hEkavDljbnNHTqvgRGEXV6XmXiSpvzne8lBbQuavwwUbnyz1YVYRx78fT2mN3Spau8JEgFGjiIX
80NFhS5H4iI4I27tMYlhOk48SVHGzd0Xk3kY/HriXsVLhVZLhJ76FVPl9em+7x97VpTIl8qsOvhb
M0AoE6N0/5/JKuBwR1VHDNJ8cnHXlqhr2E344u8Te6eNYC5qzV/jTcsz95oG3f0JD7vImz+kG01f
0BFf/HVgT7eNVgpj8MUxh+IA+Xxo1cu18syi6YXdeBPeabwt3ClQOhjuvUEyo7CmZ4eVCHIp0wWq
UclrRGTtTT8wT/eSkfSwojvHVCJwshp0Unhd/EV2fae7kSQaJYFZckpJUrwUY5tMcGSmRvR+g5V5
5MAmuraPIxpO47GB6pOJr3LxPHV0VeKQmNCbFkC9HW00ZvWHRYksuBUI8vghxy5CqxxAwkObBVYE
lYS3XvC9WF7VW0Xk0aqiGtVEjLQN1bWZMRFl1gxZCwT0mj05zGhgsY/t/4yT9fr7pF1UhL5kKZG9
E4COiv7YLKCtG14TuQT7Hxjx8DsI9hsKi3yX4ankhUFLE56xkwCDXYkF6NXN8NLFZcm+ZgcFqxgC
qzZ3YiBdHE0lhXjMcFyhJ056rUHo2Z5bSu2WLW0pahzD/mDhUrl9Zju4mYZ0Z/f+SA7yC0kJsYgb
33Jb99kmgk8e6ycG91u0rgXdB8JQ0l4bM3OKvGavW0pQ407qvs2mLYG3SQFYFww1KWz91Hnnu0tW
ooYVuXreyB9nJy8VVRGXrgSs/kDEr/nGWIEBzQ1xqhJxzbYl8om8VD6RDgo2aJ1zKSg8WVXY4tJk
E/uSDt4SQliq8YJco/wWkd1UQSSji1+ElZkFQ3UUQHJCoQbG/uo7NRY/LJsAjmA52KX1+868JlHN
44v02nT8daZR51HWu5juRLxwLlQ9Vppj54RzyXU+9ENcUvgZB08Su36pEQ7ogTrzUeAK851fsmw4
qMkhtq1kBGdLC3ouJRNJmMThQ3930nf0qP8wDRzHPUe8XmY8CwJZBxuX7uzOwXNdKktyyswumjjV
dKm0VAjm7G+hY7PQQFAa/YZn/PD33I/uLj0v14Bly0iMbYaQ274ualGZGiHhNc6PnmNS3IdqzaEh
e29sFXYCYjVKhkxEVURnnU2l+FB5O3Ss8ZDoIGfLadvqtqvGUpAEE9U0v9z9bxDDNHsbkKJL6/Rg
LeQKDJ690Re+J9n1ZccAfVQ5x0aKvCKMFGYb35P0IxIqYk6pEAo1FVaUM9Yzv4tGZSeZmti00ei8
ixk6AJ/fTmpn0K6SATaobRAWadWXX7Ydm0oDpeAcOAACP7aA5jpQ1e7ikPKmHWCPLqWN93kAT/aM
RL77GqcHJm7KFohchZcGLrRm6wZjmPGexwC8idrDlrZD3g0vjM77YVrZWuuIm8LD1C48QqdsZ/UY
2jSuJrmjyo4iC4S4H6SfAdKowrsLvULiMbgazdZ3uMQdP0sx1XiYnJzr3KrG/pYitjVjV80ZyVLY
Gvdu4culnCYstgwRKk7c7EygsQ+KUrdLtOmZyfIuIgiLCtDmegUvTijg+PVk6fa3z3/HI1i67N9H
QQjcu07gRX9IXaYAL6L935RcJrD8u849r45bKqUOGccvxh9G7D5FOJEOrgrG7kVmqgJLMe2Ax6X8
f24VBne6J3hXsnGnodQkGaremyZCaR+TsISCYveezbzlw/QkymGH+WhbTctGd7EvngTG2KnyL1Ay
JXc25FzmTc99M0YJDKfrRVWlDQV4P6LD/v5piZlwx6NfLCO+cMfDJxm+Ics5WfPhVSDyamIQGbp8
c4UIudEvHrfitDp4gEXQTD4Y+pjYBHvk3TTOmTJ9gAaibgrt3wAaRx87roDwxBLwXkp2Dfx11ovx
YP36K93beFAHfjj9+k9aTdyUWjO7kVIn7odX9chFruRjlxpyb3QwXZpk8A47SZOZlkJDVdW9XBKL
+T5Q0xtvQ3hv2sTF7xOLWje/c7eNXgcFT/9Yz4MT+A4OeMOuP4pjKl81Ld4AKysOUujgdtszer3w
85RAYBhApjHrceRQ3BEmwX5s1bxuhYjvsSgzB+uvYrktb9yt0tPY4e0BLp8KgvADCWvbHJyNUQKH
e3/EnLx/v6eGY6BFtmiAqykriR+vR/Yu/OS04LuE5DPtG20edhhjvzQbYNqEyxu0d5ccs2L3hPUm
hFVOSuJcbo4i6zbJBWKabG49KPteTyavzvCcqmbE6fwulqimSevXP+ucr5sm9coPMM8vIJ3xWsnN
JaJoF9orAWq7Y2G6lIhnEx+KrU7364o964qCGYInsjM3JLonTcgCZGaMI4cbjGVURg4jMUpA/pru
fjEtwTBHnFoklBx1BG5XT2lK8aHjxHfODthbx2DLmZpSwFR7wUP5XXJ6KbbPNuHfNCnauGI2qA6D
Vg3M+IiMp75OnFNOpeOJMZ8Poq2eN8GvPl2XsU7OW5eECPOgQIklZrbN7OWBIHAqw0Yh4kKlBVVc
HjsDaX7vglz973VbBZnZm39RYUeY4CU73WnmOi3I9whs468hYuO9dYu/4j28Z75QNd+j+/vg7Z7u
H5YDuIPLwt6DozU310Am3q6sucw9dRYyCW05yHDWIXYxrM+rTrpSu0rt60PyFQTr+XEQTHx2lBps
ss16yHqFFbNCkKBebHD7DaV4DMM4UHBRyOcrKafmYNuG/pduP834NZQ63KNWki5+4bhAFoPzFYgw
lUXyKK/6Jv/eXaFSrFA6dvlq07TPCSveCPPHnHN6hTn/hk9/rpFRVa3V2U7gVzY4m7nTzTyowFoF
Fv61RjtlGQZmAVYKtYR/yJyjAZJzXD/ia7RzHiPTIFszOq7fWZA25iagXrB+HlqxBMSK4AHdJA18
yaGquyDNXNEElb6c8ACGTh5oz0qQTpbmxuY29E7XzM7k3RjmmX7NF8WWuQgdNN3VYa2Tg7Kzr2+G
XQFxOk66m4/xPk1d4Bc4nVYoxwA0VYEEyTr0nk4+Cw6y0tJtOOtlsm7/2r+t7zMMtyTmfS+huTt6
BpLSb7/cFWXs6XHOctofF9v+Ey7d79ReW94JLbQwHdetEe9anIRG4sUrd6AVDGl4OziQkX33LKlL
Em1uv9a0DTgQnGTMQd3zvwJvd9X3Zf6M9l16S+I1OPXbrpY2S7yv8sHLegTkTVotwRaigV1EMxeN
3bofDEqhiTJDaWHj/vqPjIp2xu584fovr3BsMtLPmhyUV0ik3EY8ipW+2R+niXhSyoVsLuunM15/
M0L1OMTnIUweow8R/S8BRyWcbD3QNgkAleiuehNWaH4397JmBS1bV6hmzPKjwZyy8QAAEorqM9n7
XaMFnVS464qvemWAnfc1hPoNdgpLNIDkKUDw7hgOc7sX4A7dTHT3uo6O4xvBo7BhV62uxHMbZ+4L
2/IG8bpI4sin+x0BF0XFILji65JoqTJqX4NRJM9vkDU6H8eg3tykCTb9k4yf+FsqofDMsjY5/9S5
DFfDe91PBsL3GrSMxUfLHi0TZMHijYrHvR+DRou5dr4wuV8RkLDjXNwwBYmNNX8bpBWrG9fBLx6U
T2tKIRgx8QMKX91AbPBFWujO5UVM4nsAAIOt98ZNQ2adjGGiIve9j4fLZ37BFC4EtOhRa2z+60FG
Y0gt1xhir4pUzRCJv5hiU81MV+k47vSu03MQI+1BgDO0rNidrzx0wGXxC4jJpnKiMVUolkXpfX6O
CF57mwFg7M9w4oKrsZKL7CFYjjzs3qWhx6gMaVbvGiz2MFhO2vjzBUyDg/O7Lrwqv+D8ldQoBPQV
yp5NyKmc0EgLbXHbaobxvZkGV4Z0qDTBRdh9TAaZBaIZVUf8BOq4af3pTkSfWIpznXBLXHw22ByJ
uoVxWm0VQSLOtXhbwYFBS5w1gLadcLqpjSX/PqauGXHZWNS6U2MdDyKH3qOV2LekQG8A7jA97E/c
je2wIWVIhkGAKvUMii8xvioNyHgs9UcaCWsDf00cbjm2jAqd8S8pC5s+e88YGDA3HJ4Oa+twv9sr
pM2k6pMB/o+a3M6CcZ7WdxgnFcOScYqicl/v0wsgvnW34f61khMX5B4uQ1dKTH4vUBWveELduDaM
M/LSKPF/17WUuPMnDEiPQRZhPQAl612GWtuR4EClPA+6wdzi6Spqc5ZGW411qXo3VNgXNvgRQLMk
BWMzP7VHgxi1zyXhSLGsPdmdBty0CE6yJk4j7h/MJuhnJADxyF0T4yisnR0z6UEIofrnTYVTVcwZ
SHB4xoZ9F7oceuNRuwVF2Rh9Rn4qgDhemt/PZmh006Jjip/2iwbu5vh1eDmqXe1qDH9eT3PCvIKa
z3BLgx+Bws+gKEGAt9EvNCdp47BiAS+Z5aZhX9zhfpWqRL1c11g0yeVGFm2TCimf29aofFYbUoel
+yqcrUugMxFiFoEDliFU6aP17+EAneSlpKQrwGl91lNHYpb2TBz/zwCDyLm4jYJLM8df4QjOBoDr
cIKZbS3MGkril//eOOR87Ah7cw2SiDjXM3MHK2hBAbpKYiaqsuDKu4POT0yiSycr+4roa34lNww/
2W1Mqx0hgGJDnKCiEvH/HL/1/WNCALLL1Qi+FRYAQ9hXN57VXCQuFqWGbxK23jM8OoYpVIaI4Sn1
zjbwRqBzXIvSNfbLfgG9EePIGQ3pTlWVNJDqLuNzQCLEdbfTznOaI7W4a3nkpK1ep2FZui3YZFcA
DMq7IBaEfLfjlA+0VSdgszqqrauvr9WjzuPJHQqGACrgHXNuahZNQ7WWLCK9TgDYFLQ5CawssfsA
cp5re/fNq4sxcb+j549aChASXwFT5mnFSU/MU6ffeU0XEqOFM0kfQCor9h9bavbXab6gHNa+VLbE
dhqrQZj6qTykQlWHtqn/a402QE6bs1HFfmfV2JtHeXBnbCXN5uhJoHK/CHY3M0LZ0pvSMtrbGXO1
b6eKe2b5WrxGKMY6TZEprWlCTEIE12p7TyvxRatoGtZXdplfLEF6GLMWUUoBGb7InzEKMWvTJN2U
UaIa7JuTVFqQWXkRt58xZC7ETCqEs2puAZRG5pn9E+7ukAoZtvT4+ogMUHexinSvqPQw8H/8acn6
F2r8La08lzkzDkCjkBvxtHx9topX3TsR4roL+oeu34el2uGi7MgX3UUpCTldRMgKGhnPeVacEssf
+kynG/is7YkwzZyqC2Pla6KB/BuVyoyShLjSopuUKg3o8tFidIrNNO7RgIUPrzUOegL25zeaDMvi
fJs1ZcVXZt6YNVPO+5mInwVsQqaK86fr0e367PuZKiKcpgqYUuMswR+Qqau3OkekuPUlpo5EU1Y6
xgFL9D22WUGERmHCeDZFkg7knXNgSzxVVlRtnsEnKMRdkc37VjJKcOiUKNCciwM7Z6OOrNnmoFlK
/N9ix9JbLXAVmfSgoDkYxwqNV2bNTBHPjLspTyWAViZeI9/pogoMEwGzaRLBCHU4iaXLK1RHeByH
bRTMQaGYh9upZYSYTxsJJXGo/eMjrq6Oa1G79M5tb4g++8o2nFEsBk6+c09C28haRL6fTkqnRl3W
/ULrc5Jih/xzSeDJEjUQGS4WWEb5M/KW/V9L88FBXEDsVMUqped28HUck08wFZywK5QjWRKO9xtW
dCWJejQBHuCIKCZw6GGHHTlV6hrE/nInxJQD/uIf3e6XDYYlwyrG4c3xSaIuOZo9GSdCSr12gCjV
D4d+A36aUGv+dWXYC3nqt9JgirKbE201WXdDf3jYxDzA8oIQuXTK3+SbyAQRaMS5hGEahLm2jjo5
GFyaFMI4lUz/yR+usOKW9YTtefr1XOkCMMQkbq4PvOipysIihGYYb1aVbiZcZDjfIXFIIIcQBiW6
OHam0uhRZbQTqjQn547Ul4k+su7x6Vlsem1ACcum2SelQlEGj95RaLaetLHZuCkX22xml+3uu9OW
fzUulB0moGAsYE5FsN4exvrjH2bM21uQ0eqywUsVHyxkz6J7SdkWps/uIPReG36hStR0iiL0a11s
Wo7rXE3ngmYhYf1eHMWBMt5qwLN+7GapH68sdNlocH8T8BSmZlRxVMTFBcWfDriraOlTcYyex+s3
wPMqh3biXjCuhlGKtaRmVNLcCSc3zXN2S4EbKhpwP+A6mvS0CZrbQq47lb5TQJCTtsyrj/wysQBB
K3w5oXHljCL0YEn0DRJUsV8WDdFB6L7qGDat3DzTjwdki9fMwBpk1/R7tIIAV8qhfcc3w+eTLiQB
ia/kCE+dOfKCHh/NdSbKYiT1H/MxS7CSDocSEm9VEMAZ6YG3gjxrVu8A9rrIjzmPB6MTwWQKTp81
tjINcRElwzuvFjvsf5FogfLe/R0ilbD/ANzzZTXIAo5BqswS6bBRk4XUnCCG94Vto/ysLehgWrr1
axCOQmL5IDBNtfkmx1R8P5az26ZoKxPo+a5dZ6yFO3UcgXAuQZn5aBDzRc1P4lqFOYZfmHKrUIWc
3jQqSnlny4ghOgpLwmFnx+LgmlLKYe4OryuEwJiAodpe7lIXwWTjifx9AWFnMum5qXZbcjv4ApC2
YU/RnVzYDIZ8r7HItbec6N/FusRNIhsrudOyGKKNb7ReXc51vrKlPoF6bdmQCqSdMSZ2iDDRRYta
fOqAyz/hA8tmQtj5YeKHUZxGOC1XRULTOMsAz+fkfQzpvr7HVzG0kPlp9Z9tBugQO5FVMXsY5+72
YkQ5Q9wMz1sHfThKMRTXuo/qXDLorEy/kS3ZQWpCRpBvafYYPllHNw2RmeC14l08oXU12EeuLFEy
Ahz0iF4vtQLIqCEPaaBw7VKL7j+lBhTDVtj2dnWWM7OZsXxvWj+Xz5ARb7nP0wY+461CsgDyXF7B
MaZCWrjvCNOwWaXUz31JJUGy17pHDpEKXmdqDHVkmtJT2OG188HeZRo3npcdv6i7k3Myx2kTs/BX
kHg3kDb9dqni22mxmzw+B8wzPbmAEXNLYkCq9bINl1fkdLEqVKjmP6OGdKaxd4lUxBhiYD7resQm
Ybqe/NlDDRgsXcVLBlqbtbeCPFILgrrCh1NFc/QmWN9fZAQfqI9hg6+PTNUxmrd2uR98owfZVLPd
VWrEhW1uUyU5r7lCluwTd2YD/wXCa1L6pZIMTYTviXAiuH08nRqVVCVKh75wS+ZjpVAfzcaVMupK
g7hz4x89xpcnPFP/ZHIIApxxCx0bUmIROO/rcHOyMeaxJ9Z7S4nL+KNqTKWzdVkm+wIURSJr6c8j
bPBeelWnCFQSScxc4P84a9ihu9DW0FY+pFbO1e1mO/5bfAVvYyHnYtTbk8SOCgyN3G+IhB38aWWu
4wFvNY2gW396Soq4YwtV+uP9WEsCxSNaUnhfCWzulMSXuVPJdLxgR8albQ3RZv59m+DEuHqlTEjq
sAqjKisv3N4NRhD7lYwAwX3mR27d/X+hC6LE2zydoE67m1kEUu5J/8xFnpKvBfcdY80pIXk/rzQn
47RLdbkvurVcqAsLyPJH0xdhz91FpXByexbwBi40onfmI1oMMPjgujWbwwlihfjpqKfp+d9uHmUm
CIi6N0H4w+04WV4Y8DdNUQ+0efu50albi8vcE7VFS7UcjrcN1wrjDScO5GrKgMZ6zedidbEMtM2X
No2uBvazGrEoy74ATEj2FG0iOeisgOyDyz7c1daCyWu18ZX6bk3cIUca3y2mNTrvGWVTd2h80DQ2
kW8nGL3LSvpVNV9nYtTDeVyaO2AsL9YUc4yIjZlnD4yn26lETLjc7TI6EwgGSRucU4ty2R6w4VP6
JPbxZUjKOr5gvGlons9lfS1aGLU6ixzVfbcaoGL1OpQIM7ytYsi+VBlwhsa2Qb7pxV5LKnp+2Sv9
r2L7lFoP6qMkc4SoJrvfUeBqCwKeVu+Y8MfmdBaoJ9QoCAMHIUlVbWzEMm4pBuHsVP7k4WEKEN1a
3fwmaFs1NS/OT++gZhE0H/XO8Yg+yHL/DxY7GxIl43PRwtJivVXTUxsj1UtS7uili2eUwpA2P028
yqyAHLuvpW/MeANHh/kz+t9ywWcLHcwZTsvEwNwpOnAvhNI0Slqhirh6S/VC7BAwyu+2rR73dnI3
pyU3KSgFUjoFYUvUMPqtp/V58Fb3bOu1onEkRJ0OUuH+PbsRS2J9UuckMJBgUmFRQIeQn+s4kP14
5bK8cKtQBoxMgDV3pt1UrFPR7WDM1KyvsHWdCnpf+mrqwP1uOKtq2gvn/4lQZObWMWxUyGPc/oup
IyGel7ZRzj8nq6ue9iCcvLj3QpKQjWDjI/Ak7aBQcEV1RF9SuMADy5vm2g+SH2j67kdxfKFrUVp2
KVJh2Ehdosv70eKPJg7sr7+D6jU21Dv1U9VBIihnBQmb0Gj0bBAdnR1q71LkIWzXFygKCnCygT+e
2IEE/XtipMREIZdJXbRVca6MJL/UMxndjhPwtbXw4VOTB+mY/yR7pRV/OJGpiDiqbIU473w3x8fY
n2jH46BQGihpNOxn8cjAGhk5ZePkW8YGdMAHcQF3McC1wap392E5SsbhFrarb06ErVri3dNzH+gM
wVIqRse5Gx3NSiC/6e38guhM88D+Sw6BlI23wxs3jwSXhO+wyCDthJjM3xKY40zsHskPtqcvyafW
kGN0gXrxyUDcYau1yUmvNaXkTeGottbadiP2p3DpPT3YUE+VpI/6D1IWHT1x5kwmM/fKZD63wEFd
hyVRmybPIMB7ubCIojhTBsc3LtVKdhr7pv+WeLvw7e2c8CyiGhw5/Uhzq7Sb7k4r6waTg3IaN0o4
AxJQ0KX7348+LhGfL5crqkFjAOdU4vtmALYWWL3Ta93Kufv599QIbQwpVC5mLy3D7zX9vIEvo2Y6
K92nMYHLI2lWuwRIC3+gvnd1RxxBknTrsgnrJJpl/j1mn2apUwbq7JajQQuyNehS4Sk/tizHmGHz
Qnyd82JBryPWAozw+Q7fcVAm3KrUezjE1NK+L4OecKdotrPNPDO+TwcvckKLmKvEYWfQqgTngABS
fTZBMLfxGTjrTmy+X24qhZ8grl4Eq/bKaFkufb2Wn05WokTHzIY4yiG1/Bc99yZFMSSPtJJmqeFE
fTcOdhxQNTbWNBIWBsL94yAJ892L1Z40AgAhXeIVM3cQ+nq3aHEOEmRgoi5NC38ACJP37fm2iUgS
trkgHBE2uCP1GwCZGKPXYU36lF18p4Mg+yuAe6qnf25pgIJWI3yDT1MK/k0yY2eXByDX5dtVDuDP
8ElNMCwl5tyMCzRaxOWGnyZBL8sUhY83ir1FiuFsT66XTQrIBKqna8qmTQFIHit0BT05kmPYXuQq
M6aT/HoCPH6Hz6jGbkKXafRYycssApL3VKhl/H29F+WPTcDSeMqb3ibrw+cNF46tarJ5LZiTGPVI
3xSuWqhPTBO7SFnXRIgW2NUqLn2OcJr8jsP6dJ42pjg9ZQnYXv8H4/4esOMoIoMIrUqhPRDD9ps/
L33wCC0+gjpjMkXKXE3V/rY86IkSXWpp+scyl1wygmzEAjDJJwnMUVBEsU3iRgttELhF1kg1o5hn
YiqSfL1qBT5W3UF/lbCue6wg4tV27EzFdt5CJ4Dm0ZF3lQb3NpNuNF9xmlEU9VabRINy4kBX2utE
wfrJsa6KOgs2exfDSJg2wlVByVDKN8gHdQtoXMv18tdNWa06n0mnUgXGu9qYD5bylk1Klk5BLoWo
ctJb+UoJ6xCzSHAFKMslcVKHMEULClp4j58q9IjmVKNSN9xhaHGpALf+BIpy3eHqsBNKdRvyWhTY
OcKbPF28JlvdjSNXrX+vU1UP2XkpJ8i8RH7Dp9RVuLJVB9Sum/QBx1DzTDtPalV07HOpmWleENMr
IvSj1hcastP4FYVgN9aq0CRSbpEufzRpZsAc4vmyVtQ1Cxz+v0yTSKFODhfaMl+enW5e5jchNZjK
z3gcTk+Gg4m6UdozQtr8xm3QGKVRRCuRo6htnjLDZ9nZ/18C6BLMGqfq8jL1LkZ3Heyg+xU2RuLK
/0n+EiXAUmwQXo5FUuK48E/N6Z6qQSGH91gXSaM913gzVl5kl6gNh+Gpj4KT1gl6fM5Iibz++bR4
VtUeVjFSOMy4oXA74fgBcWkd9e01/NbSNCy8Qs/GPesUbW3Ggt1m8o7Z4CSGqSvXFvJ5xK0de315
pWfE8lOfdOPpGyZziBFsiFtpmLce3OPWXPbXN6khcatJoaLIARTq9DBUH/2UwT3vafySK4E9alNd
tjC1ZAGpG7Mk3veMBkK542nGr4P1UMqRRWNMbrrnYnJ4ciVkl9xkS95kUZk78rV9l/ex9022F8lA
6diJ8K2kAflzasPS5pH7iOdiXTGWp3lKRtR6TsBX+AsrMOh2kmEs1AB9CYw9UlZ7e+Pqg8g/1t94
TcUXkqSaCMCWP/nY6plTHPtwCIyrln4GszjhDdRE6NU+7l1Kx3UWhOZde4EQVXTYkvPczrPA+Kgi
2fdp3C6qWb6yAto4hX0gTEyIKDGFhO0B/hrq1sBz2ojjkYQaGYHon0kol4O1IsjthkJb/znb5VOO
43E3e1/Kl5A0OtD3u797dYDF+X5CLZSzyTfZKZkBDknVtV9gniivawCsyeblxqX4ZvcGf5/H7QkS
zaqt1DX0w9IkDaY54hoyqQvzNnsd0UM3Rsptqq+QLXsdX+huGDEcu0phFdoveKWAwX4xfk+VivU0
jpPpGEBPSkeOIFFapT3a2E4C/6uCWTCiHs2TPMXcRATLRo3X+/3J2oVIK1XZfocap9VUgZiSqq0i
aK2QcWRyvDecgYUWgM7APLjapijQsP1WIBXmKxVjHHnLWUT745VFNbpzhP1W2b1gdVJ9/KiA7Wxl
X1GGYIKNL+wIhVZtnH2X5v54VBt9vSpavQFV40o8EpYfOSp5p3FMgmwMrwlf7SchQSzwhyhh/Pdd
vwd/fzgJnYTNtOv5Al0Uq//lf4zezueg4Df+3Pe87utUcxQ/3/3Iq9W8Dy8EcYVU4nMVzodrI7Sw
X8cGGt2D2u9Ma+tjirTEFc9ew2Mf0d5UP7M10ho41UK9WaNiM5n7P1u4Cq28SfhL+H6r7h+ghugp
8VzIde3yZ32HvRr5qnA9Ruj6MYvGU8uW5LQbqunujcq0FwvdJYOTiDKNku56emEWXYHvnZRgAsML
ec7EsY7jZz4+hg/GWk+NxMjCb9cFkl9YmirpRzhOflj6ZmHa8ytdGZSpRXrG3q4ouI0XQbwy3e5h
7LpysBG5DvfgK8nVf8VOY1W8UY50xBpVwJ4FIAge/eUeyHPI9Kv/CFpjP9002oFS1p7gZ3F4QpLg
SxsMx83nVvEFoPKEXVSpe+uoWbUPwa+r5Fa/Ds8fplJkbNdWlAOX4cXHvYKP91VopcGyY47ZfxEx
/9IsR2wfQzM9WeQZj4Y6SAok2RX5fPYvHJMXKQ4PCSUC7liNr6W72PSwMp/oKxspExDWXaR16+3i
bfRQ3PV0cS6PYSBErcj1s59waVZ09z0WbXAYbBDZ/QOhk8JM4JmDu7oa2ul8hXRrA/Q3ZUy23dD/
xU3Oms5O0CexMB6sZHnaF/m++YQqLbt1rnGdCkF51lhQ6N6Yl/JXS+YkAFCJEsMRrQR/TihDISqk
EbDRpAVA+9P8x7TiVQUNxr6trqbEdVqxkJ29gcgwLZ6aPi4xXiDWfilKoFnEOIeyLOqqc7cCnfyD
Z4gtXuohFOoeZu2z3I9PU805mRyEOjkWlhjD5Uk0vLgOtxQhTT2xhgc5lsMmORFHd1HHm5gmi6wF
sj6juz+Rpjco6nayfTLxswKHxof4Ab6Z7qD84w0DWRGLo0yOTei8cE2HZAl0RIgu5HUbPh9Upix5
fhEXDwWHFWdSb3ZaBSSmQZ/i+EsVZZ+fUghWUftiNATR0Kn1Chgod81A3fgZlXxwrrs8wY+WJt5m
IFe+A3TCAiPaYIRiDAQ3MqHnWpXagz27kfAdVgbKh6kdD5xXz0M0OsGVQDdczF83Rx8suodsLOFx
kQDbElSxHmQG0xmYwt6Z7xwvrKp04raYk92KFyGBkZkOh//WvCuEVWMgF1yfMjqF+asEnR0vi5MO
rHN3wSO5ThskCmYsH2C7ieeMJYEpCxtq01lsWsg0eP1vimScctl0bhmzDmQ/so+N9Rqc5/eWxKUX
y1FTNntC6pBIL+WyWjgffoLsEeHYBKV4V7oE/8yazlGwIUq7lx/C7+gHzkE7fbko1VbY5M3MaVna
7RxB4ReVpWibnNq0VXIi8betjM0bNZE+NwF2KWOLTmIvO6DHwRQrWGq0mkJu4AnLStstq/QybbsT
bOVH+Mu1wuZcYX1DaA8sgW+tWNERqrBQgz/5Xy2JaiLGmTQha0TdWIPC1hOUH58DVjb1bVyxUjhA
F6vEEO4c1RYz+S/qOAItXbY2xR5bUa9SSgsXPz5VugUWugCydfZfNngto++Vp1njO3MHpqon4t4/
eq8PnGgC9BI3jCDJgYfjztUWEm7vYN5Ld4aJJQKvCd3/HOEKT/ge1lnwqcjZx0Lp4C+JcCD0HQBW
A30HFaIfhzF6qWUdXCtH+qddNhUHd3eFRXRAoxcx2kTyFqDF1xYuu4YiqUE/GRXAcL9EI1prHgbz
9yS89cI7OB8zzN1IESAbdmI0Lf3e3nw7gV8MTi+Aoz5VKAN6+15AfW1aqLXXaDEEgdoa70RyPe0k
O+7H53b66ZVsSCHrl6+V0MzmNNAH4mGq8QkPz3JtRlFgKbgoGukOdPCkN8lD62uZ6eBeHoQbIeBM
jRf1EmVG4xuEmjqnRKQY+zQi+LN4YhaV54/37gJFx/kCtL+mTrBG/940Q9yIYN4/IKipJpVVi8++
BslncvN1zNuwpdqlA6pc6u4Q5ijc/VoU+L/VdmAk/QGgB17NvZJmY48ZsBR7L5PezuZptIS/Eqep
44vICCDOd3A5M5EHwXq1aFG4GQZopn7fn+dvKRPq0sXr9GNKUW0OoPyxbJDmsKus3FaubN2G1+Tt
q97Z+PJL6T+uSLIwHDB27sf8tezTWli9jjdAxVT0lNURjk7whAB1GGYVeTUuE7+NjCnG5lpGMtZ5
csGz1DR5uVwR4iCRpxLUlfw3L0JgR00O1KpIEPcE/Hczn9DP1f4oBLZO0EoTuo2/pxp19093Ip8c
wEnS+em5k1GiXc1vYyJdv8PMud2X4XxJ9jedQC7elOGhEQbBpDlh8BnWmNa8tCUziawDy3e689Vm
7Erp+k0YaJU4bVWLM88OrHM5biHvplaJcHRlnY2G96Il2fxtEO6vdNOIZtGa4sqRi+qA1fEkLgjR
25+GHO9yPfyHecZTv3hQwDI1eTc1iqIzmOPtkm8Oq+GuZ9Lj47hd2aSQ6cLJMA5h1bz2Io/Ca+RL
uFkasIRctpqLlCAEnm+w1qKV1WHYK3elV1j+SMoryID8SyFoyNr0UZZZzb1GuEABRTu0Kb1jUU4p
q5UzqxIS6mZaCTMQ6CSuE1laP03QINT3egbwP9DadBp14RKlc0uET+1fTs6o+vY64vQjRZmMsxmo
A1JtBtfus68xTsJdR54FpgJhL1h/LBSqkGkxkb70W7SK19Sb2CSPWl660KwPFnnVclV20LARzfAU
gdrSTkN+c0JT9lGK1qiDGZ8H0OcNIkzJftSr+qzpJWIRb69NPkwx3hcu0dveojgWz1An9XtiKhLY
YaQBjtBfYIAxzCbow2ZfI/DoIDN7A7V6trSSl375njo1/C5UXc9skG6LxN9ofCOCg6f3WD5yMudU
zR2N98U/SrDwWWCFhcXIGoW3+1aYlkugUzkr+7OHn3LXekqhlhmoeormxSEjzRBlqqa/40qZMo1P
oSy0Fa+/u6g7VJEl2+vCau4ZtEm56X9FDOjL33rmXvsYMGY6EDjJ4tPUm8cjmt3Ca33kCg/hfIsY
5gGZzGSwEKyFslD28+PDGB1F+yacIFIYBMB+m9r2YFZf+dDctqlGknaNiNBOkp289mv+rForgUl4
7+PavoZavdSy8Cj+8wjOIuDObHbVpCXz+MQxqI5NtOfXqZoel0FJSjlIeuepTP3Sh2DZehBdwtq8
dH3htWjuMncrEcVZFl1ZFQSHD1XujUyvBZTWa/6cUmdwWwZOw+R1Dj9ptghA42Yv8SiWyW7tfIyK
vP+tAjCA1FYduR/10l5ixJWMkEUSaAAY/78r7llYUb3G110iOFVjJp7UVQiv/Wsr1uxB5y46AZra
NjO2WmH1qMOERdS6HkXPpH8v/AytVDmPTxE57SHPsPw/baPEs0+Bn8fCykW3R5I92HULqi6XONL8
/spbg/Qd2i383SIlYY48xJloyHiTY7WcF/KydgaIyx0RNH/uMUMzN4lAcOBT5FKU5u2vyXsBPWKl
3+01Eizb9He1y3QTPQv4FM2bgW3fMIAlPv3tOWlFrz6x4qFNt4iL8gOXHwwlZIQZWoazyJTCYV3D
DQZgvhc7j8BU1vDzJ3RnZZDguKEEt0t7XD/TdOaWwjl3wPtNmPXuQ7RH7Hic5N5JvCtOUeAnM7O+
UeV5vNPR3f+bRJWhb1TR4o0oQ9UmZoytuVnj8KUTbdcvtBFulDqvSQDXGapt5M+cBqjqg4IoiVei
VRqPodnMIEjrIrh/WTh9LshqokQhpVm6QKckR+n9jmwao5dIyb2cFhacHvcc+XXbGsKSQPTYQJcp
WACdHieSgglR6ybI2ExLZbIpjKyi0I1cEtbKIfvf0om7Xs5NsTAhcLmfrfv/gSxw2prpKgPEITbx
81TptZZoHCgxUaa05I4JjexaYfbE/MHm1fW8zEmLcw8/H0cHSiz60xpQIqu1bohQ1jQgSrbZEf/J
cLmIJpXJhOvyD5ACz2AkW00UftZBBQrH1CxUY+Gzt/WYoEkHC8XcU8+y5LBrhxuJ0mRjV08goxra
4roZdJh7CHjsFeDfd4Ks36QK6MpPiPo/t1KM+mUmB2emIDY/1KQWG7wEj3xy/xmWe9CVeHks6WAo
uJKwkbIRR2b+E09xSYj+UDcQBILvd2agrIXs9tNNR1tdbHz1IdgK48Nj5Rj4WrrgksJRn/RVxEHy
eCXBQoeV9yd+2vGTXinDhZ7ekbvUnsrInYmqHLH7+x0v4o4qKmP2OIWGDuB4hLoVX3wWmI5RIz+c
AdZ18PP89f7HZ+uENhIkGTSuKhGCb4Weo0qc1a2St0+FqfSrY5p2dhmU0yp5yTc31GyimK4ecutu
z+RJNOqo6v6zLC4lZFurfKYrpDtlCevSQDn48ORffFnbeenXNA1WVYweDqbRak3YHuv5mubJ0uHt
m+mWfO2Xn8EKj9mWaSW1IoqoySFQYEGY/2hSKYFBbVTGe8f5N/h/C7izH5MYNg7uCbCU4zFtc1EN
jjWX0P426gSh9YcOSrGpuWbgTLk00r6uq5+LFZ/D39NLDuq7s4t1jEoABN34UiO3wsFVFhNAwM2q
ryVGVlzXeLUzCcwO5OUg63szO6WiRxriXWsgja4Zbwm0SNEErQyvQ1tK3K2U446J6G6oDDbTzVRZ
KNJu5HVN/UfMd3+zM8Hi+8X5po4eTY5wetuw8wlJd7uKfhTplVsnjPYiWCzOqd1M9NhpJ+rTnO3e
LwOIVTUjq2BKzhcf36a9NqdxWd0q7+QQZKk55WXiD8Zgqae2rtIQWLuyCS86amd2okyqtaaLwUI1
NqGARQJ4z1h72zjXhlBYvwuWfg5/Z4dY5mMFHdJrjdq1Kvocgvv7hph6jeKuc1F8BvqJVLrVHE9Y
PUMUFJSciX0CEsn/y9IipzIJFGBa9IOW0fhele/w3F8UrsTYtJNtPfJ+luZCcPkhpxITL4YOSC/1
eyIDmn2EmD4BZVfziY15VflgWGZYJ9xEacLulEy9N+ck9WvHVNIoIq5APbgsPjU1NRGZnV6Wh5Dq
4TZ83gFNggBVOkGlAIh93Jn7gwD6I1v0XmYS9gTHeu6ksEe+7o4B+Yi44Zgbpj19WPZb/ATm1FR7
vM8bSmget2Sxx2duUv8eAAPgO/2zk8+lR+WC8KGfw1HPscIS+2ttZdg0wTzyZTer7MG14EPIJp4D
YhKDKQNvj7cuc92UkrVYIZM9RsOLdBILj56BlIzcAKpNwYV8yQuOerZ9NVDqpNhnR2ZKj1L28Mf5
YDfo7qfbzO7AHTlJl4cRRF0fDob3hetmnU2f+7fUwvlblBZiLjXZOlyqg1PtY7m5yO2Jyqa1JoNl
dtIGTJ9FmzQd+Jyi+8QVL3nqw62hu5fBuMpzxkt7DX4vZBBZI3+y3zo0eZODxlEwHUvgYjgqE6Ck
PeK+QEVLF6uWuXwoigc0Zv1pYejhHMTnbE0GQ+Fu2N7xa9iduVeM3Qmzlwzy/wYPjFhV8bTY/pC9
d9RCX1PBTR+/tSm1JLj4e4i/LYSMNYunOwxbtAojyn/dlgILS1BoF5V8LpV6K9CLmueaZGP59uDZ
C3KyjTpjLlNmPK45v/jupg1RHKhxboIeQp7UaY4gt7bY5q/PemC7b8VmhlfTlW6DGCTnL8RWI4mE
T8wlYF+vOpVJW2HuJot5kAUuq/g+k4hGH97/CrY407BUO7QNQwl8PZsZ3bdGNlrc/XbQO8/grhMD
Jir+Gjc7Pmj84ZDtG8KjdJ1EuEgNMGnoqLwUM2KQ2dC9daWtZBL5Y0R+hyJdeNrFN6YpxMEs3tbd
j2OkxcalwV5nX0bfIm6hAzRPsQvhG4/q63ItMFa0V7Jc4k8eCYQI8GvufOMneGn7XXrBI1fCQCtw
PgnY4wHEv7qYljQyr/g04G7BxFb40FOPETDaUTmM5Uvwq6ILXPkn2uWvXV410uGnKPykuXJIUfR/
2LWEWEu3DO5jnoHeB0SPTH36hSkapljauFRjTcTH8883/Sw0Cg2mksf2NmLvf9TPULll49gjPdUV
jyqierQAEilT7GlVK/HF3kq/6Wv0UpHSo94hGRam56cd7gb4zy8g7NygZnfXZ+e276HYrDGCEjJ1
+dWi4D4SSiL7+7DpvnhwaRKc15fWe0L7LkwZ7+1q0DYf8g6L8W9ZsmgeAk0zsonrSE7R01wjj5BB
vmEhL8NAUGhQnBRwZOkPZaDC5uinqAuNebzDt+Knsc6zLpfdhc+qHBIh2ohzjiTZeFExP1k1ZQwh
ULpVfEv7sNcuwGBAzUgIqBoFsdfXCR/sxNixWx06iuX96Q77iTbNlYCLUqmTGGgy5zwdXEfOiHcY
Jj12FFu9dlagW4PnGKWOpbwoLQST6EOIdlQB9f0jEeNl6xvZ/WS4KDpKwHxWiQbMTEMYmjALv/BI
L8yU66sGdAnCx/OVElkhbpPK+NyGfTx/186UC69MgvDSpYL2m30SyVBNPyPOh7M0Woqng80q+joX
IMcgy+Wf0TtWZo0/reiG6RMrMuTwG9sb684nVE3lHHLMmbtlSK11sz5kXfK7s7WVjFSQDXcLjJiy
6CsdLOE96LscVUgajTQflsEw2EZx4JdV7ZKtruep1TmigT60YdaM4sOy/ekydOQq9YDEuSysJOId
NOYkIdAjknZTt86JI51cNYbf+YcUbnxHISMBG0lhQyTm5DRooRHxswoRo3IILshKYkCO4CdLi6PU
lVXIdXbJTkBqm4cQw5EgLhq218NHW3g1NVMPoBOFaAkzpY52MOAZ5TgQsj4Fjm3s+Q4bxfzXLhFd
NXfQAmTc+/VKfqiJcy8k3sKkV4V1hTYUTAK7rGr+cEKuWzHwcKoYDqnmvTF04hLbAflv+azSCkB+
e38YhLLDzssA7QW0EFyyDxAAjc8J2xmcVgX9uxxknR/i1K3mbyJsWukd63XUP2IyV1CH8OJ4I7P2
tSbpCzRv4rW+scE1db1h3p5CUh6YHM74e3uMnWC6TxdOldWZHcQY3Zk9tDSxyX7+Yn5sCsE3TekK
50xHSGoAjzu3y+kJLatKtYqxZBlsi7hnA8916QDgtIQF7gs5BW6G77BLGlYksuWWTzQgdri219TD
nLSPcXkBAQwVPynb8Jz6I94GcIWuSpT9lpKHnhy7IVHZuX5hJ65G6RiGJjrq5+Ud4vbO9xgw1UpT
a6mcMT9MiDqXvYVuB2pZMrXxY0hXvmqX8mue5SKSEeUsJRn02FlNnKQneVmGi5TxeFFyIgNnq3to
BeFF+wuDtf2v4SVAhQ4mLzq2zn4UdjLdEL/45Wq7lSaAahyf/rg8WsLhaxKT575NGJXbbg7gPP/1
29U5O72QsN2VXD3op6v0Dz/7YRNudDihuSbrk2JLZXOF8e0dy1vstSVFkSVP+m8hMBhWIa9nlR5z
bKcAnDT68mEWhVZHTwbSrS5yDPNCQ1ScQnwUC+/54COvQ+dfntZKMlEna72lH8haPy+xs9qW4TU2
YzGf9pjvp9SxjR/QoJrzJ2Kov6zonXHEc+tXAD15G6vUZYVAyfR83/k4j+xUzVb5xlVLRbocF+DR
vSfxiHHBBklUVs+EDglaP1YX4dY0wJznvVJJw/CfB8njjFUnH1yAv9O5wYYNSG3x9MmKOwiF88T6
Nm3PzC5mSNS3trYi6EEJqQ77sz/jZCwQmH5dxLmNMy+lEIVZ2tiQFPF0zbs+JxPth9/ImiVNYg0O
bBkkQyUSmp8CNhJPo9ZFnar+hWaFVZffg120K4IP4CDcUkMUiOEXtYo1bIKGojCsAF3X9bf+uCLn
zBEBHET4BKx/VHchKWDc1rh9AVGR/jfu3oGUce0/aOPSD6MH3++pQ+H2d0fBWMiuW/aATh/3YoTT
UniCJIyLlGlU+drN0a57HwcVB6Z890+rATC099qoZ1Lawtc02sziaVRSUt+tTjXfljYKMvo6ksvs
fatckmarJfJUiJePK0D5JLrqpRadxKKNJGvZhBJpOevVGNW35tuG4CHUL4uU2v8qlYGsy5KVfV0f
d3lPr2yFP7huyJJ2ssdMYvhs8HqvfUq1MN+3HyGd34nBPSYmfxUwWotcS9ZZticq1lYLwLSXl8Kl
KgA7Bacacr4hvCl5TsSaMXrDwlUbnAL/WIqm4Pb22tBAlqHojoPUT6qr3CN8CE9ltMGsYEIIf0n9
kf+VvY6iyonXdLDPwSaRt1fmifPoZqcDAdbN3qFvvCV0TlFxfik2nM3n7tR1zvVOMt0kAqBOBdBS
vr2X8xW7zMAQuq09gmZba2w7vNb0KnWeHV1ZRyKzFAmaefV//KmN6C35hc+nZZCrtaGpqg9WWdrt
3+ByUCCwAfzFcU4/1Q/hIZYr7VjT0DMUpTbxhzrg54gHKQbNV0qnhPxi2uOQp++ociY9Z1fo1V/C
O67HT7U8rrLaym3fdxIxtYNGe5UcWyfzC51wBMAZ5/y3UiMNiqfMxLOml3aYBREW7wy47yVC5Zsd
RODquNK46dNto5HIprLXer9b1xPAnEiiY6yC2IkM3EKPuixNTf9aCgCZiUA2eNFRGsmSQNbDfSqu
gcgs0Nuorj37c3nf8bmSgSbgHblZ2fjqnzLpnbxjgR0tr3/tcqlKtaZxFXL7aMcpWW+5fw4BfMCy
OZjkLqLyZn/LFbjmrHTDnuHfmfMhw8gkeefxpqC3idUcCS8s7mQKmy4Wr785smorT2yCPcXNy8i6
NcE8hd+mae6/DndY6MVy3VSWvpnIY4ujJYELspBjAgTH4XuyV1CVj1Nh1SA00FPYZsz324VX2jry
kK28tMHsg5az+yjd9BJokqisWP8jX90p+IjUNzKrnw4LI3N8YEGPn728rUFJ/yiwLfRb18yqrea3
yfUZl0k2I+UdxAT2plo240N/8QnAmS2QOlAlVjAvoacXPtkj5p6qv2bdk8hLrZaNznb1+b0gdpx9
El3Yg97uwZ+4h3MQyLV/EwJNnIYelBgt9cttzzpxxAMzVPMZnY9xoIMrM2g6HMblSsqKgDiHAJ8Q
e1jjfR9kEjchPp11O3U6dnSAfoGjdZ4y0lRwiESRZROTtOAuyJu9z/OHZjGFQB9eTGdVTzXPIA15
MafeqlHmLSbbTQlzclXMDcI1yULh9TxfrgKXyNwpN/1Mw5HJsg7c2i+CYZzZtp7dafRewHShmmEz
XMukAxk2Q6bzzPG1FD5skT2Cs5+W5uvsOtE9qOyI0EPmXOI0ymEcGhFJIpFq8kEXD7ftS/VXH6x+
c3pYd/Y1hr7zCZWdsxPPoidwu1OEO5vTyNRBiwqcoOxi3lBGXE/7stsq49vR1dwuNTQcXgmbratY
9GbuJqEvme2+NYSnum6I1JMVLjDJDgoJEHHGllasaf9jhYqIgjzk7UAB1J4EKXOIU39P+Fge4GIJ
7aOpyX3INuxMF7lbv55vMqOjbcO95TKXhsybW6v72kroVP10iCc0lIgX9E+90f5TCfU2XGQqSyUu
AP9sw8WMdkIQKmNWwzGKzwxCdcFdqLIuaLhIsVaX7P9nlYaphrMNVms8sr7b7MnsRraTZBfWp1QV
ZD7rpCDjZ/c88ffclejr7Lef7NvBZCy2y1DrtXYTkt0aJ6rc9OujE9CMKN3bXEhjFYeeeqXQgYIG
IC2KJPEgQFUx4E7pwCtjq9m5bUFy/Zz3zBts3eecIKJiF8+YjyoDIyCZuZipJawLdhBThzVhgcTd
mKHpvibKiafaVizJcQI/OC4U7mFkoZuzhvkSpQEKnu0Qu7KYCmyQV6T38D7Ke4OdxzKqsE8vbZJI
zzfdjvhhc0s4PC9tLt+gVApw0yuRv2nrYd+3H082pGU3CT5fSjkBxmP+zGCd90BT5jrnT7XkDNG7
lJvmyURK3KpftpUxjihqBd/ktWr7fAmVajOlLcJ2JYOX4CYUb7P/TVcnmotaUTNFnqynoL2P4i1j
beNShoP3l13e3ADBwkJcRPCWnHMp7TzBJkrBLymSau50Id7ZKLJ/SvBX3e6pzC6PXDCGamsXyEeb
bANXx4E6o3LC4NIwBGnHCygENximaxqYVhyb92jzRzv2ZiQ+h9IaIvqz+1Rt4ZT/cn16tZH5Swu1
6nNsszTey4/lmrpMnB8Vd+Ld4MbmXvVJTzRk2lTvAdst30zpjqg3nHdhWcpTZIIkpYD8DbcF5z8p
e/Wg9RgN09UBKjSX5/cLvKzmbYn1KZdm76YwNsJpB9qZ40Om09YMQsOqPF1L6X44zTmZk5NihXUr
5E1sGYu1ldsQ18vU8YB43gfKxYkT1oo3DKE39yOP1KmxCBeScRUK0T455loVAa/bihqT13YE7orm
6WWD7dmWoEJNiii99mEgN6BxR/aO5Tmv0eZMvKJLqD/AHuaVgDIlMecSo2jPLY2/DSwzXBnNdPAw
PulEqD7aSH1+QeBSJLmM8GYEUvfmZYWNu1Ip7wg6xzknA/+E+oXxffp7+fIco9i6lynWHbpeKF+8
eSYx3ZuyxzQtywQ/vkDvxabp4dY+WqQ3RhnwKHCyBltQIYY32/TcVaaZ28easCcsJtzml8awltBU
VGMdA1pfaf3Xqylf/BaOPjuB+AUDMIxudacsSaKkN/bbOWINCaVTH0OYzvlrwlBKBaS6ylW1/C7c
D7jAeGg8hTPhiSmxp41K8LnTHtGU700tona4tc6JG+o/5wv+PJOe5QSk5rK2oAj5synwrIzgR5xw
RoVdzYl/FFeSCwbkZ38a69iN7zLVOnrBjjvi/KpmwaddXR/oyKSzkFuGZmayWv+37a3WMRm8gewi
HwdeFAEpgNx8Tt7kqA1PCzDEEYfjwZ7kdgW+jK2VH/WxN3sN924TNAMNDr6vl+0LE9v8qU4KHvv1
5LJDI7Bwv8u39SI/ZPmYorZgdi4i3GgU11b+vWhZt97w6I9WWYaeBJFWsi8h2rMJsOlmrGbudVRw
RNXNLqM42qCEXgnH0ETY3HtEVTYpNm8Ro/t7/CtXbqarKefW8ONf0Um+QE9zTyrU0UP5gYFjc2ts
twpsUaXck30HZx21UoxchEvxsMvZ0MqzMuUSBRPHj79U8+Ajd7ED1ic83cq4cu9EKmPHQQ7j5ZRr
xFQLGdU5ew93hXK80O9GpiYejmnjNKMEkDg1jchqHL6y8P1AwqCTSTahbwE4XlFAcFAB7AEhIpBA
sQxVvshzL1NR4L/N2pimzP4Cpq2MjxEwKv7lg8Lw0QNay0wKeX5c9ENptJtsdRJrWec+rwQHDbvj
kIq5H3rWgkwXgpzOg9+DMO5e4NEuN3v2T/LeuMlpzK6TVTjzvC/nZoSq2iIcTDazMoNO6CneGAgx
4f4C69wqzhZjyw2cy+LXmp7G++jZ0CGPNkhxUiyDQUTx+S3HX+eJuErEHNeGF0lbN3wJdQtifnLB
wtd0C118SzBHxvMZ9iOp14RyBF9eryTbu5L0b9KKKt00/bljb6AuZoyfkF9bxTUE6ROncIYsZ8SG
Eap6CM3xrg1Ybleq3KenoLkf2j+QPDWas/ARn+JHp8IqnmmhVdFaf0BL2GMwKgkp05WDtoyiJtBs
N/R1DUQgRD4rN3VIei4Wf0xOsbhdVSmKBQrDKAEu7VFySfe+OxG/kSIdS3P8QycKv7GNNm6tqRG3
P7LrKIGpgB252NrHpx6A60WaRznNl3Rcve4SGCQo2tNDvHSnHJu2I6YlFP1rhRB0Lcl+z52eJ4ib
fI6tXUCynrt7BVvTOZp2LNX7xhgDB2ZzOsbX32HbCUdxzPAgotKvqSd6zn6u22rOkieXxxa1RmWO
P4rVS/P10MuslKLFfJ8gLrPlAFvHLr6T3exukew2W/aVJNAJDlH9hfQ3eo7EMBijTZfJ6L7LECFZ
tKtU6IF6I6tmdQ9kcAUBxNBlB62ERQZtcxjhVl0xI/wmzXtwKm/nzmVCmPxnoHFsuhyBo9uNZyAy
2Rug3lKlL6JQ2f/g8UAnCQEWHncF6Xs257e++rvr2tliiPWjLsqcoR4q5hfo+XO4RZSaj+5IQnct
2DwPmgqmC+jxNo5UtjzvuOWy1MJzBy8pjCnEs8uCCD8K0bPJdTgTwHXMewWeMha1hh9lESbWZOra
L4A7ZBpC+2cw6gzCtcy/5f09t6N1XZirU7NbdeXc+dMHUbKQthYQUGDGkoc02bt8I679ZzliOTc1
PiRWJ4d+4q3qrEW+7sypxJfmGDbyQhHQCa7sITWA7WoQduyeBefL0Mnrum38bStOsz8SGjcL3DrZ
WLn2R8/eB+9ZowM489W5A99DeSBs/rOPuPQe2w41Bqrx+vkQHVTqCu4EJkJU4zbLqBRGzGlg16yD
8PkYQFpyOwosghuwNpnoY1D/7OMlHB9ho4pEGfXxJpXpXYXJ/U+EwFSnLe4YdVeQ8hD2FgSec/ro
W1oa7AmgWwpR5HHZCLc08pz/NFYR8c9Aip08pclBnd2nMGyZ7+f1xyVwdy84cqENdP5+1nqDtNCP
DDGzx3+0A+LcDs8VaqbIkGk3Yjj5yAqhTJkqKuQTs5bBzOXlRAtEegz3wqqdYIUPuWl5fvxU5yqM
TRqs0CoyWO5o8Si4ygxJDKoRtSwN5M/D6YQJhbf9+dhQkOQFaMt/68rPe9DaBy2HcSoec+89ahHB
zFt5txnnDD0m/hphUo0132UV+IT80Nnrp80k4Z3RhtI0wAmYTj5/9pDKhja9rhWxzcEAt8Jvwmv9
JGJsNReInB9zD3Lrz1zObppNxStujI8UvSNSCTcg++JHHMI0gMIptITIcIGd8lGzxxORCauK5fhs
3iAsszRvvxWVtTPUO8TO+vMEMBP5eBdhbClPVVahbPuLBnzAY4l4JaEbn2eGVoN6hk0I9rTMOyz+
69vDahPHuzFQ/lf+16LgscvUeqYuzhb5RNxRrF20hcsBo/7MKY1AswVfCfHlN185yxqjlbQpPiRs
/4JiX+tlWNSktYXWgwHiCbXSowr5JlpDCbascthXk1I39Qyf071GulHd5I/o7T/oLW/rmK2Nwx14
b0Y9W+it8gVoop5/OdiOHj6w4eAyMyoENSHWv30DNz8eRynug556AkN6tGyL3zo23lB+yfYl+g/o
i80ZigRmzV774ksqjgOO3B5X/TfUxic8RVEETTeF534jcL30WyI7wILN3cF3lBa21KG//ZDJF6cg
sivOvmmxGwef4d7HZNJoAeAVLm1f07C8Nw3RZGz1iffTcE7NJQwNb+Ifn7TMzGD9+QuTAfCzsHDO
Kgfy+SAxEJHBsZIIcWDnLMnuekMYtBplxMXkhWcy1R/HLo4bApI4fn7+q/AtflyD34yQAY5W/T6K
QwNwbfFrh/mUz+U8Gxkevjc6RcAYYFtndwDTbX0qtLZCpAei6iDcjG2dJ6ees4kV0Irsq/gPtt6O
h5nmn2eQ3mW9uEgz2l0DbRCKOSUOMWbDc6Xai+AnxQbqQ0qoyqG4+E3KI1jVaoe6HI505yVwbsba
u0tC9/4wQ/1QLytUbQxCm+kxmMdwCDOZ27Ur9491LwrggGQ862R3o9MTj44UU+lsCa12rAD76l4/
09Fz+SGl3QHpPZPUaJEZZ/XCnSXWge8PkbaH4wPpipCVGM6bojpsZsSMbVtUTzSixuFfw1EzUsIU
qHx6Rhgm1e/mWx4SbiWiHn0W8QRYoIlO4Xar3x38h/oMB2/4fGyljJoSgxJzufDH075PvADhEAKF
Vs0lCP3eVib07UnDy6ypONBQVlD2M4cezYWLtD5gDNiOPXON7FJw6qafrbvDNLAhpWfdNrLtf1YA
aTzAqRbzmMW87ns8DPwxyEMpcggsJoLBTjtEL1KXi8IpqWmK6RhIgsBATdBNkCDyTiCisbPwQU98
2R0YMhu916/wkZQLG3js6YDDd/ntCkb9hpuuSGGuaXRfMnpNFh5bgFFM7PuMf+edMT8wEZrPLuXJ
Tx3v45lRPwWaKQnMJRR1ovxi0wXZPScozP0rAT6OT8u0hFQf2m15VwGouQ3FipbPld0rxAb4g8g+
9H0Qpt2P4mE3+sySSldjTJ60pC+jYIiQ9+u7E+vPqUncDhk+WB5Irpg02gNckorbdcn2Obj2hGWl
ZnFIdTVirMCVLGRlj8UUBCk3uxjmR7g8x2fCfnr8AkVAOnH7JrWD2U2gO7k+yfQ5oyJAhJtqfjPd
U4x+hH+uUDnGsVJez4FiRd6UobC3uQwN5RErGpKmBSTLLLAF1XZOJ/lI4xlL2RRzt33cPWnYuI+z
jDhi4k8+Pf07fHWMbmbf4zO19nhsSDYqtFcbHQ5GHGtE1BNPMX9ROLF2DhmZMX7QTyacC5N4r21y
r3VTMtYz2qDIdU7scPlX8h066ldQFKy84N9N/T9432pKE7fbfKjSxYl2C6Am+WjHf1QTU3OHDwxP
sw1Bf+YUrFiVzdxjGyucn8ameAPULfxSwp4PZjvzh9dledgXFpW3mQUsBLg8+EWn3/j2DX+K99xQ
6fNaNilSXpmqxtxmI5I0TFh2YN+dXzk5RMwE6hvqnxa2shCAvd9RurPi1RlzV4Qx+kGHCqUzJhYO
eQatu9yD2HOcwnkafyC0d8cyF+KbjteiDuVma/iy03pKcpePoE2Vh89jKW/xog9rWf0E6g9i2HXH
10zp+Y9vxSyrcv27mLmfWzyHJW+lbVnhKNts3u3cdx/7rFZo3samodmSAZW2Q0S32ooayPqh6giN
Z0764R+yTiYmA/5LZV/gmZlfXvfkp9t/yQnEh/1HfoWEf+mdW1fVZXfDC/iCM5zF6zFORHHxdatk
+00g+2xqpt6nqTzeu8zLoT95bUBxKOgZOdJTvvrG2/cHMcBEBzTqt7Jrhl5w5Z7z6FeiuRTgOf89
abnZYOaFkrMa7I4ujN8fRdZ8Xxr5FxwY5zKj9llzYwvzoTnEbI5yWIDvV+GpFfvvXn38aKTU/pN0
uxr1y3UuksZ3I4+fSuzoGmrKl94qivLK2n+oSxuq1sIOth6yLQSKHSN7IwT3cf6jnrr3c1Omki5i
1ailrU7v3q89xir+G3pXkXAI8CpIo6TVNbt+9AbWvIZ4f1f44jpygY3LgHlZJXYqrtr/K0D1TzzV
LKo24xUbHSfEVfe6qaY6kklagHZ/QhZZwbwtACkULS10XuPd789iJ6vqwZKhAY0s/OL0o+VnK28j
c/tKr79V7P8Qv0Voe5usxQBffnrqE2EsE0p/GMgKg80nVar61AzDajDqR/JJhBv8elT2OoZELD6q
66egxjq0dVb0wqBLt4zx7juSVPNj1x/f94azfnK1rW/pbCy6KqCyGxgzQp/vIwXR7c5f19AgSbDm
Ko1nxq+qrqWApE6VRsAKJFwc6ffMGAk7ncDNaLLgrRRPCEUeIam10UoftuhBe/dUT/ldktkZVKmX
LX0orM1WeBrpwIr8UTgI6Ja2n+00r5g2Phbi4VqoRmhGwLo1ZxJml8VOYl5s+X/IAjfTttIi3GaC
6yLRFSCGvmq4KN6qHQTBEnpgVXXdzmJGvYHGA+B6znx1TSeqUMOZdS7gpiO7eTyprW0acU4I5nmg
1x8ctlj/eMgcJNiAlG+yd9akVppsKyxT3BUjtsKSzMPKncv5dD03zWNeFQFt9SkA/yOReScBbXXc
HYEhApqHuhLOrgxaa+K091VdXmjAraHIxS/MloKgqUMinpuPHmCbR2mzFHw6iGgdYt+Bi965H3lo
udZZ+T45j2n8DlK2Y2YJXDRHLJ328c7rG1IvdhpR+5Ko657Dv0/cIEXa2WbtK2E0tOlkc/ALAjq8
6jOigkNcmWprYWOqrmWJERbdTZO86+/6u9cA+4BWNKK7lO9sznO64e+MivIaSqNKA1lk/UDOKFAC
Xhmzm7fN9JIDuhZute25/mLh8Y6DtXzeoQJW3ZepapP52JSiJpVBlYJT2VdRyqJfrZcGN3/kVAvt
xx/nC/I/thuqu9gjsnU6ELDF3Bkski0dDEkc7CY6ACcLdlmwcYDBEMECZX1BC2Z7PIgET9HrooI2
LmpB+E4kSrEvhiWAmYgOkMyjJGeajcwAsGfxK4p8zSCdPOkV2A9twynX6OLtzgVC2o4uHxP7exvC
6BqJ7eyQCvefV+phhtHVcQ==
`protect end_protected
