`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: University of Arkansas
// Engineer: Tendayi Kamucheka (ftendayi@gmail.com)
// 
// Create Date: 10/02/2021 01:36:30 AM
// Design Name: 
// Module Name: masked_decode_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: 
// 
//////////////////////////////////////////////////////////////////////////////////

`define P 10

module Masked_Decode_tb;

localparam Div_Out_Width = 40;

integer clocks = 0;
integer i = 0;

reg enable_counter = 0;
reg clk = 0;
reg enable = 0;
reg arstn = 1;
reg [15:0] c1 = 0;
reg [15:0] c2 = 0;

reg         r_PRNG_enable = 0;
reg         r_PRNG_load = 0;
reg [31:0]  r_PRNG_seed = 32'hDEADBEEF;
wire        w_PRNG_enable;
wire [15:0] w_PRNG_out;

wire function_done;
wire m1;
wire m2;
reg [255:0] shared_secret = 0;

reg [4095 : 0] mp1 = 4096'h048c093b06160622095300e604b9021d0b3c051b088b016109e808430c4f03f101be00550771059b03aa01270a2d09d005b9006f00d9017e05c70aee085e0b090a03054009ff063b006507a106ec03ba04640c210864098f0882052b09b5042e00da007e08d308de02a10637047f0ac904c307bb0111021f02650c6e02cb0b3c0c5403d20431013409f800b908e3068e090f09490088028b0ca80520057e0821068207ab08f903ff0b6e075f0ce6039800b00a0b00660a7b050406130418001e04310bc30516081e01c90a74002605f705270100059f032d043d087a0b7b086706fb09ea013e0c5e057a064a08ff009e056309e5061e03930b770ca102e70c420b890bfd0c89012c038907a60b9c077c080405c609500659087a05b10033097e0583044e00fb030103e0029d024c006307e0053108d10af108ca0c3d037b054405f00a6b03360b960022056b0b4607b10c71075b0555098505aa00d2047c04f702f20b7204ee058108590b130ba00629085105ff0ce308570cea0b4c079d067e03d7096d030608480992045c00a50b970ce600ac01b20922008d06ac06fb0254074605c50b0607a20901040805180be508b1092b08e606fd0a6501af02d809f80b6700d502aa0a56098a015e08920c960497053e0077074b0418031b0b9c068e067300f402a90c570923030d00680c9c084000c3083706b402d20a0d0366006b;

reg [4095 : 0] mp2 = 4096'h07d904460cb000420a2c05f608dc0a7200db079b0b7e0c9003230b4406fa0305042d067404a2084e026f0c1809e10a0f0056068204e80bfa069c082c040d088c028b019e0923060e060a0bc90c8d09a0081200a20a27094f0af6016e02d301a70bb2063903dc0ac60aeb061901f40206081a05c205000b7e09e7072003ec08f30121096301a70c5602ae056903af06eb0a0d02fa059c03ff06a007f2083a0afb005a057e0496022501c804ec0706025b051b030e0661087501500103025a05a1024a00dd025c0b7d0a3101a3007b003d07180b0d012c0a3f026d0b6d073d0a770ce502710c6107c80120069103400be000f502e906570950024b062502e800d707d707310c790b9109ae04db01410b270bb500a40a120cdc049507740cd00a7d071307f60b6a09fb023f099d04220cf705a3014104e802e20a9b076202780082008209480abe083f0ca300e908950c2107ee0beb004803da066c0c1d07dc0765093a017f081a080c0b1202c8082c002003d7003a05e70a93008e083e0458059902380a390a7703c609ab01ca0c5b07480ce70c0d0b3d0af40bfb061a05ff0ab400000140011d0489043809bf026a07c0037c03ce04120c5a09100ae60385098e00da05200a320999033e0b6103b9063d01f0081d06310c3002c20996015a0c3d0745055503a507880af703c8058b00d304be065904ed069402f108f90384066f;

// 0e4d12fc0fd70fe313140aa70e7a0bde14fd0edc124c0b2213a9120416100db20b7f0a1611320f5c0d6b0ae813ee13910f7a0a300a9a0b3f0f8814af121f14ca13c40f0113c00ffc0a26116210ad0d7b0e2515e21225135012430eec13760def0a9b0a3f1294129f0c620ff80e40148a0e84117c0ad20be00c26162f0c8c14fd16150d930df20af513b90a7a12a4104f12d0130a0a490c4c16690ee10f3f11e21043116c12ba0dc0152f112016a70d590a7113cc0a27143c0ec50fd40dd909df0df215840ed711df0b8a143509e70fb80ee80ac10f600cee0dfe123b153c122810bc13ab0aff161f0f3b100b12c00a5f0f2413a60fdf0d54153816620ca81603154a15be164a0aed0d4a1167155d113d11c50f871311101a123b0f7209f4133f0f440e0f0abc0cc20da10c5e0c0d0a2411a10ef2129214b2128b15fe0d3c0f050fb1142c0cf7155709e30f2c150711721632111c0f1613460f6b0a930e3d0eb80cb315330eaf0f42121a14d415610fea12120fc016a4121816ab150d115e103f0d98132e0cc7120913530e1d0a66155816a70a6d0b7312e30a4e106d10bc0c1511070f8614c7116312c20dc90ed915a6127212ec12a710be14260b700c9913b915280a960c6b1417134b0b1f125316570e580eff0a38110c0dd90cdc155d104f10340ab50c6a161812e40cce0a29165d12010a8411f810750c9313ce0d270a2c

// 0e4d0fd70fe313140aa70e7a0bde14fd0edc124c0b2213a

// 014c 05fb 02d6 02e2 0613 0aa7 0179 0bde 07fc 01db 054b 0b22 06a8 0503 090f 00b1 0b7f 0a16 0431 025b 006a 0ae8 06ed069002790a300a9a0b3f028707ae051e07c906c3020006bf02fb0a26046103ac007a012408e10524064f054201eb067500ee0a9b0a3f0593059e0c6202f7013f07890183047b0ad20be00c26092e0c8c07fc0914009200f10af506b80a7a05a3034e05cf06090a490c4c096801e0023e04e10342046b05b900bf082e041f09a600580a7106cb0a27073b01c402d300d809df00f1088301d604de0b8a073409e702b701e70ac1025f0cee00fd053a083b052703bb06aa0aff091e023a030a05bf0a5f022306a502de0053083709610ca80902084908bd09490aed00490466085c043c04c4028606100319053a027109f4063e0243010e0abc0cc200a00c5e0c0d0a2404a001f1059107b1058a08fd003b020402b0072b0cf7085609e3022b080604710931041b02150645026a0a93013c01b70cb3083201ae0241051907d3086002e9051102bf09a3051709aa080c045d033e0097062d0cc705080652011c0a66085709a60a6d0b7305e20a4e036c03bb0c150406028507c6046205c100c801d808a5057105eb05a603bd07250b700c9906b808270a960c6b0716064a0b1f05520956015701fe0a38040b00d80cdc085c034e03330ab50c6a091705e30cce0a29095c05000a8404f703740c9306cd00260a2c

State_Polytomsg__masked_decode DUT (
.clk(clk),
.ce(enable),
.c1(c1),
.c2(c2),
.PRNG_data(w_PRNG_out),
.data_valid(function_done),
.m1(m1),
.m2(m2) 
);

// Instantiation of PRNG core
PRNG #(.PRNG_OUT_WIDTH(16)) PRNG_0 (
  .clk(clk),
  .rst_n(arstn),
  .enable(r_PRNG_enable),
  .load(r_PRNG_load),
  .seed(r_PRNG_seed),
  .out(w_PRNG_out)
);

// Clock cycle counter
always @(posedge clk) begin
  if (enable_counter) clocks <= clocks + 1;
  else                clocks <= clocks;
end

initial begin
  // Reset IP Core
  #(`P);  arstn = 0;
  #(`P);  arstn = 1;
  #(`P);  r_PRNG_load = 1'b1;
  #(`P);  r_PRNG_load = 1'b0;
  #(`P);  r_PRNG_enable = 1'b1;
          enable_counter = 1'b1;

  for (i=0; i<256; i=i+1) begin
    enable   <= 1'b1;
    c1       <= mp1[4095-(16*i) -: 16];
    c2       <= mp2[4095-(16*i) -: 16];
    #(`P*2);
  end

  enable <= 1'b0;

  while (function_done == 1'b1) #(`P);

  $finish;

end

integer m;

always @(posedge clk or negedge arstn) begin
  if (arstn == 1'b0) begin
    m <= 0;
  end else begin
    if (function_done) begin
      shared_secret[255-((m/8)*8) -: 8] <= shared_secret[255-((m/8)*8) -: 8] | ((m1 ^ m2) << m%8);
      m <= m + 1;
    end
  end
end

always #(`P) clk <= ~clk;

endmodule

`undef P