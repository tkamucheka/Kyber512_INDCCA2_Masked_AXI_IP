`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AvZ1PdAwW/ccANlc11J901QBTuVYl8Ao/4ZJVckvhTAlknj4aYL5gGsRltbT2iBV4vnt4RFbwQW7
1h7inJUsZA==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
PKZRAUQbH48LQwOvC4ffWn8rzps5t3vFD9bQELmuNezMlTvEQ7sVXsuUaQS0L09qKXxIoA4O79hn
JRzJa1HWOKAQlDqCGuifKay4Ok4hHZ67rsY8x2KHzB0VW9VENYFfRR/if5Cdm9XTlYELayJAa2UY
0xOqjCUXp0tA9IL2apc=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pdmj1lc49zjOMJkOAEytaK3IxLkiX3w3XQjV0jMbHDHIHHqEyecSsfK4TSzBbvsoPd3lq7+MDmdj
+IFge89RJOJxrWaKh/reSJSQNDI41bDC4pO9cZqExOtyCGtis5+qoOi7Smwb6/20a2Ty2C2vE3hl
0rii4EWi6qtkgs3Q7EvzDPLgY/pSyqDg7RVC5oefMIT9P90FHhWFfoJQLNIhB3c4HZq4XyoyJYxL
p3Nhi9D9r3MK7cZoHxbmFSzfSnFd1DsCi6Ot0Z5+XoIEs+oaaNCYvZMD8qvmqDnCVhanGRXR+G0t
GUui8qaMMsxvjPOS7gozXr0uJjy4H16lhzMhTQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AdXmEp+99olhcgYMbJSpozTLGw41PWch6bNb/6uFlWegW8XQCmvagv1E0qtwBSXE8GCiQMGS1U97
j0M8whENh7C5MChS6E+6bJcQFEwnpXXEB9TUsH5mh0auMHkFw0tO+PHBMHIDhDl/n9/TVnz0TnFx
NsQ6TodSR8pS6MBvUfufGtHQStRBfC74q9Vdn1DOKhTQ+ovyBqIUC+Y54v6+wW5so4f39KF/zS9a
lD4yxGMEdHUPZj12ZvfFTEMxKgUn219+dfwZpCYd5OdYrZmsHLsd2/Hn5CRRJBaEH6UnULD25sgb
YlQUrZNS5Pq58W4oQkUR4zapxS0pWZvTv5CUQw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
J8fMKMN9+GinXD2Nc5HYe8EoPZTLbvgje/DcjeH8Odp6mXo1gb8Cq5iDp140bfyvGA+Cj2ow0VwQ
/UTROMyaNM3QMtLbM4KHq8hNBAwxRupwEIk1vdI167L2LN9r+Km7uxcvj+7C6iSyvpr2mUCuDP3q
77/3TNWAOiYbmsk5DHRJt2VcZK4dxKvZymsABtbiPBg5/JUDuO080QknXWkLEcSQvOqysy+hQlIn
fHi+3dk+0x6iWwmOJ0bjJZrKhgvi2hE8BORtmFY52qypdTEX9C2L8zBDKiPFmP7vYHOeyaUHbRsY
ENKBVKyN7KjdgXp489GbYD9e1vAztxPTOMBmiQ==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BUSbCwuoEQ1xcQ7gxCKUMkeibZqy+5d09pLHfAXEUHLsO9aPdNW4gIySZmx/P5t4e2YOeAQYAzeZ
YjJnRlZnaxU289aOf44nkHTNLRvyrIPM8llrOUjzI01w9SIYKRrM6Gavvk65yncB/dBVTvZRk7MO
WsybsklRK/ZBCFRFxLU=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mlPc8GHem63DqZczGsjXGZslztVjlO4daS3aYGpXpO/4QA7Hm8Jrvlvevj9Vd8fHlDcun31xAxMO
nmrWYAkNMSuZ5obQ4yid+0/77F17VzY5JWAEilU4y+fqSwCEakrhWj0Ueae1YReLTYlLLaeHXLka
v6sg5MfsnRGIomBIs/0dln0X/p27ijiI4B7w8zUT9ckpVFFMhlXURGkgGkIM747gG6eaXs5MNfIU
DJzpBesfc6YXNlMloLIWVKPXwlWnwQxx1NrDi+XIA6io3RtF5HJaA9ig7ZeWiJxOszdlWp9qATc7
ugWHLFlG250QuNiaOZeZFenKpW20pC9b14dwJg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 132688)
`protect data_block
k0/wjaqYf7tMSgOjwPlRvBRm8KWo839DxVun5bFlhGgyICROqHBpHVB7Gqaw9Gm+jgrgm0dFqOKc
vTp2lqi5B5WQ0W//udKhFsoPc3OOisHVHzokkkNXsAfKqxNkuOA7CXZR4wH6nn9GeJaw1JMC5SlA
cqCuSaLo3fTpRVdwQf6f4ZWEXuVoDtzs9VDeSxDmbb0vZgq5gipdRJt3QGv521re1gkx6RCzGaU5
HGBfStTLrvkXDqRbrMZAm3Sl0mnlm7xcUzUdnzzOS1b2xmewI6ALJ0dqNRTLeBuZUnDhznRbkuO9
r8O95b3VVygDyxqIVDeZ26rXmwa8RdySbNVOdUQ85AvEvV+T8oXW9nRaqmeLxrtJz/5jpMaS0caS
RmaAkXn+rw/Z7+Ko6wV0lqbOYbryDqe2Z/mwscfLaDfB4pkIfUiVnt2LbwyIKH2wBVlABN1v+8bA
SGMtUe6JdWnVr+/iUMH+iw0p483KuN0XzlVHbvSH5na6GDD0CHPdmyRnGO7OnWex9hUVZSXYNaH2
rDv1qzQEE16y9ON8uG5wJF+64++JZpvRcnMZV/bas2VuZTl0I+erUI2ml0AUgv8Nm1DwMPv7M1IV
6ZtBTwDEKtn1Rj3e4E4r72yRpRDa/K+DztpXUrBGXTgMD6eFRag3RrznIhuh32V/tNjUJ/GWpEw6
XwsiL2dt0J0SRo/OHW0Q36mgAZdk3877d9YWWbux0MW1Mu2Nox1B7axcmquOvEgNTLA8giSuPZ4U
gX9v0NWWZxXArPdPBRQR5RuTFO6k5iJ4YXbknrQNHBKAYtoCyf/9lxc4stoJdsOVG0mKmXWIqoap
DjOnITe2zf0ty9BUY1aMiSWbRLi0lA0EuYhVwBIvcCEdjGsZL68Cmt96kCtUPcjCs7oY7D8yRHnk
0bEUli6n0CkDP2ULKlND5t3QwnhYQbh0GPb8QWWMo4oRURG+yWNX9XOpZI35TarHnHc3HfWsJbFs
iwevOs9YhSZuWyr1M09JPbwbSXIGbOX2cTjYdtKZcFoRFItHAFWs/FIE11crEuUMUYhYHa8Rj99R
h0WcWvKinVaT/78ZZurtIOZET2V1CueadXbaIXzwBJf3U3gcSZNaj2xtaf9+DovRgPTKlTNM7fBj
MoBbwhii/eMmTk6w9RSaoqW4y0PetiKWwgnMYFPCOw7uLSdKM9aUxx5rOptZPKxDfPCBZaQ302L9
p8EtjKPDhXUtv3Cqq6nw7uMd/SIWS96rS2F0DCbwPBexWSFbftCrSgZ5JhRmqX6awUi6EluMCCfm
OS2o8NGMJQuvikPAb+QkcLaqGMHQQhZBcebZYU3I12hwbxEdrO0qqLZIQB6W0nPDQARNr6udeKuA
hR773gHUN8SdDJPMgzrty7F/zn048V206WiXKSrFnTxWmEiAz7xuBn8ZxCW/kcEzpAxVB6jy79QN
LOC4vsN1Jzc9GeYLSbhRwJqzF4FQahP87wcjZxcBCUJNHc0JJTiO9i2EHy+uOLxb7q4VPtWXSJLJ
//yMeZnQ6edkbgENvkKaRzTHD2bkDVMg9mQLcOqZYlbWYGt3ihSqH9iUCemnpUCIk6KOqclmQWcl
hRdHjqBC7J+zU5wLmmuz24dTxR32xgvv+3JKB6jiwginGLEMql5Mxc3sbHVppeqjtlj1IrJ9w5/+
WHw9DvhqeOPIgf4pnqqlQC0/1B6PwPM1Fd/96FQd1FIKmqlLbLpqt7GYKMTDISLFp/f1LnqjTxTU
ga6Lsf37sgjB+HI5ssOEJsoFT2vGCK6PXYvREyuLtMZVdrFpXq/8/BU6PtPnrzhw3I1MdZuM/S8S
FwaaRu0UB/Q1DBXXwixGaakK4QyaS54DCh8ifO34pmYgkSw1I8JTC4xqbxPbw/XfQbePloLqQNtf
nxCmjOg/7yjlR+nXaUu4LlwCbDerX8VCASp2rxTFpKk/X+Ha+irzoBIjMoj6KxUDSh8KZYaTJoYi
awRcqZuSGqpRpxAAetJ2vEYUifVdbTfTUfrNv12lhEUgG03bIoHYYRZGTdXW+azusqUa/EDgrtVs
11dLAJpjnNjujbeVb1SNdAhNSi5BrZkUMdgBDgLuEhwI8kskyOE2678MB7IghhESuwxJSgxZhTn9
DEHVhgqLq35UBhs5uL0HgGzH1tZnuI22i/58o4hM1a7Q83FSgiw4CUPdPQHwb2Ddtka0xrxrZWPS
ENslScEcEDPuvG58ScVrH7lzAF9FJ5dBbuZJrLe2W02HnM9+Q45Z8RVS1uwi1N9YNFlAilYQEx9d
31LgCSfEH2Rvlop+H5o7C6VudgiSKyrhEKFodHY1IuZ4XeQnxP+COHeSBFC0wPDjF2yUnNR9ESqt
xTN/wfv3OU9rXfVeYW6Rv5xNQZZ67yEqRtDUhbHkJmb2JAAd/Bi78Ko6hojaHwKpd7afUjq2ZfI4
Sw2eIyFPFoXJQvE889FVWb3BYk4cSlGSnlRAgBe7hvhOdLj2xbI7CVEVmWbpPUZXr2iK4++NVv6H
d0h8JV5emEOZTw4mBleFlsdqvj44u4z6b8BpQXCi2GrTF61p4Xk6VCQUEk0t5FzxoGRMP8bVTJlS
dpNqEtEcNQRmyqJgO3psNcFW7RMlV5RnA/zQ5NkEvRyHDt+/m3jiRTvM3WJm2+Csw+FBJNvFV36I
QqjE7wtAFsZA6ueNPItDIjjJbZQXvqAZC+81KPMqyRUJteDYdDnww6/LpMZeX33AobezDX5EOmum
j1HxH1NZ9v0FOsLJxkanIhTp99kb+hh3fxqUgUY3ktPTHH/y7+gD83+B2DvaESNZXHrmqrbm/0aN
KZE1ah9j/JMT5rLFZzwIY0dBg1j8lvx2WKXg5TESRZt2dwB0ScUixNvwZjjkueCdm+BFaUNpQy8K
A4BqHUD6qyb050ErcvivPHjTaDyTDXiCwzIk3stVsW5MH0YBuaccRN2azwZc3WrxU8BS+g8QGz+/
PxFFq3IhvrkfMDf/jZ2n35jL4iYEVhsjnMGmJQyVvovZHlcHkf78sh0pCXYriJGI2uu+znwFEblQ
nlwOK8iL1Y2zEJV2O3lYtNbt64BQFypZalBQswqdvdxcNEqwI6WI4bGdAPRjcAF6Wt5XXhVnh7ch
hGfOCSaKPuSIgB8/ohxIxA2/OiaMg8LcclwzgGZVHT1mRyid3Md3udZ2Q4FmTL5Go1Chpf4Vaq6/
NeqW4C4g3VfZhGuXNGNtpRQLvQKvmVE0KU60Fqz2tz9a6YbU/Cl0rLWzd++uNqFMw9AcDFlq8wkq
5LBnR872XG5jq7lZCqj7XfFu8YODjO1u1gQ+nhwZQezwi/QAqjVZ9t/S9ZAYMiTjF/O1uwyJ2mGK
k+QxE6mAvljQrRzwSMFA3bBJbbBLMK7OLOcD9zZTIHLYmptvFXuLbYLCtUZXby6Ygyi6pt1nkK2X
Z3q9Q1RGXGD5I5I59/N8eUoycfZuk9h1n1vh7UQIE+4qc89EyFjHd0fwYdWEHYTfrz4gRbeWcJu+
bQXbD/WEK17zkMEIsnC44VN4X0Amtax8+9fZs2/Ivk0BwMUs3yHdST6ZiHkP2jd/a56Tu74XfejP
F7KqLbsRKoQ7eDK6A3lzi2ceSd4IFZJzQcdnV2nW9MivC0UcCeBvT82hYc38uEBlS0bV87ERclrE
AaRbaCGHFGaY/8cXk2/OhQjcZHO9/hfLJpNnkmKvjnCkIeO65xb5AlUohEE2M7ruR5mQklDTrdLI
Ws6DFDlePvV/HsOrUg9vuzQjNUnFwAcUK+mSCcCPeczPDEc3sk4QBrfoWC7m9as7truDq+MsE7wO
0zNpX1KErmnwBJppKJ6D0Nz4qlaiZUGtDjqR6umT0YbbI94P1KSxW3M6r2E+a1PQTMXMEhz9bCa+
SkzrAUBZUDXGMybUSAYl0Y9xovcr7PEr0gfOEBH6Tp7fBcmStmRxEG22yXMU/SudPiDrdWnoaUyt
CBmsG502WKE9orvMEd3Ywmm8ETqS2dNJwS+ZS5xp+vf0o7Jag/2Ky7zC526DIU0nDScHIPhW/pws
l3I0Uqptd6F5F/aKfDMAYUZnlPo133BCtlfLzn5PhycQvbN9asA4ACM3hyWcuYrU2u+109+kqW9L
tC/rp6v9M+hm37C39/4keonzoqs8ssPPzISVv1nXMO29gUIIiEo83XJaodImHLRBHhSXT8pUdLdi
GpFwR2hhTDhB5+0+j65McVs/WkuRSWurUCrzQW0SfSZB39MVD/HZYYAyvC8CYQmZp1OB5Kjk6pVM
JHxAUNg+E4A424nSAZE/ACCI5q+AX6kwAFlQhc6nzSJG92HGCXAxZPf8eH4XqHX118T4JjXLCJpB
ZX/c4mHcUvkz7WsS88KDmrqI0iMBvVC4160HXivHySyqpzyGJVIELYhC+vcNyL2imJCQ3HLXV8K1
FqseR+9/u+9M4Bjh3czwsxSpHCBp/aUZv8mzSEZC29a0yOXhCFdAWrTtsSrwupG6OW0PETG+oEox
iBCH6YvpbyfVzZxP38czUe/QrrE/Kt8Ofs8d0vYT7GXSejbnFmxrXxwVssmMZaCQM5B4YIjYcrsW
LedyMqQDSW+Lj7k1xV8NOaNE0LLqBBLW3xMzQMBoK3uRrCM2EqoVZhAHUj4TGDMqi8nw4KpT814f
QZlmxNWM2EcYKNkT0Ltd6//bgT1RrY7pioeMWFF2cHu/JwEIMYiuIP1+rb9XDCubX5lBdNhQXBmF
sDOKXEJ9ksr7CyEGdP5gsq4vJlEx5xOiwU+lesXxvelG7KKGKV0GgYzo5bkrfQukQifQ9ZwMdCx7
ckP/lNCFxvxErUl1vlH0r9smKiYvYToAZUrhdCrvcegJmIr45kY2saYbWJZ6xyKcotX+xT7rS65D
Z88V0HkZfBk3qtWpS0J0RGXW+UEUmufDbt2J0QVOWCkRByKewYrFZZuXhkuJEVss531AqEmyAye9
3fmC6PGSrOZIwVwSwJ8bp9Gp+ubMzDrfoPMx+CaUDRpAux083iU0BB5znHOT0ugPHgNVW8AV8kUm
5plHOSk2/C0jEF9Ak/o/aB3DgD1/LPyRoXJW60A/6e784n9UWstFTGjsH88NQkUxKpX/5VYzFUwI
9KQUEPOF6zfMaZ2LcLMTUD5mOCH+dy8pwADHNmlxkqJFJ7ylrv7HMtHT4hlFCkAG+lKhACeqn/cG
ZJV/DcgyqCdirMqNyqB+woQLNrMo/GYkk51VJjokjpgB+zFx+cv1i6qkPrELwUgbs1Wjdl7YV5xP
379Sxl1hrmxg5c88VsxmlEZ4alRzBpEmIiyXBLMflYI6bkGl+jbZLghabBxHi3Xs1Aa7MIrjnFuI
Ro87hrIOS2Pwi3ydpNd76q91P3QHcu/Y6SamAl8rYIaXy0g8z8QJ57DVkRp4qxvorkveIkFRGD9H
nQV5/CT9xOyR103q0op/ZJT6aJq9j/WF/JigfR6DoraVcIOU3vbShGMrFwGH+FWEP6ULQi9jYVd+
vQsLwroIPXd/+F+yeU21yp4/MQ3UQcFtuy0TFFE/w2wtU5wdtFfB/SIy/y1leqqZsKp/5OV6vrL0
0QdCHqqStHvLMy/+446XNN/Tbk3pOZOk5+pYFTVb9NIuM+quePKvYQnEBt2wApIOuG628/IVrJJ3
LbFuDOM3oFrRe4TL8qAfQyj2Tyk28h4FNrQk0vnIS8kJggDbd5EEX04JexzDIg0WDtXSQd95HiuC
zt0M/7FKzEIsMmDwXHIYbAIasN7uHDFqr1l5ikn+lGH2z+Nmy9lzuthu6VmWVJoOO3A9LkDnX/Bp
WBQ2on9WSd5TqHF6rkRhmFIvMtuikkc7b0gfEkdAlm7a4la5Bt2GmpSU6Sa6wHGrWhfkAwW7UMft
KrNaSPwMH/DhQUXggDnjgxBCF5b7Z0TxxjePObHf3iD5MBuNnRGLXbZD8YJZTRBzUdy+sI4B0LxQ
utb8+mcdQUEkYirmlldSfJelTv+3kd+mOSsQv708Ysn05+OcO4VtQipO6EAkkXq8hQVrnomzWS94
RcSebKNbVryU325FSN1eC4YgBD8i/MTuKxMGmH/binjbbGcnTGjrjloNx8t5dxLVI5efBvF0XFh5
OR94m2Rt5oIAbFablluDiVVm5Xrb8jAB4T55isEY7lHZlNHaEPxq9RbyXIe36/g8AFgt7dnwiz1G
MUPtC/0Nd2wsTm1+czMKTsGxlN9E9vQHNsj46a162TLGmOnx5IPLGBLjHuOSc4Pb0+ygryfgwIrf
Sw1aW9zdmV9q2FTsM73+WoVzWosPggUQLrU9qTdt9vxFhaTibUNcuSUkVRotIZ2u7BgJBS7M9QpD
Zw38Ibx0LaJXLiLHISOjjRs08gDL/lHM/NDqbgP01sXJ5ZqU+Ks5poFSDb/l13EIdzw33Kxh+aBY
vpdY4LkpgfrSHAg+Qui7rANfH8wY0fsAjalUU5HLM0tRD9XPPJGwcGyH+1MrtKC3C7Z1e60atzhv
QRTmeTEwQ+p1Atdynkql+eEYLts1kQbpP+KLshj8lUJIZ3x1/+M/+Y8HvGnAeQFciFbWOMRdEF3I
mlbG9P3gyxStqrqCh5fwRQT8nv5wKn+r+JA3V1pcKYG1ywmEcFMoXhQyCTwnfN+pBUPd3mkveChx
G3TJMhs1Ioc0Ry/46kReIUtMoXclcTYNKPbselO1PTYz3yrCj+B2Fgf6CwAN5bNKLSRHK8DOYak+
pC4BxTKjuAIKuxz4rCy1gab1Y0UWjmnaB+JN+96NVt/IzkyD7g6330wyR9d0SjgEgPgqW/lS9Q6I
f1qK8wagERuPXIG0+rxBadHAbDh9ZOnnEA2iFAyKlYwbZ5BZFwZAx46kWh5+MU5PbQtf0vpYzDf9
v4DbUNB6wo/UXNXD6f1fv4oqGFd+NQjvGJ+bigAl+fD4M2WJIUvLKGmNbnj5jCT7GwFZm/Vph/+T
HcdZP6L58ygyIU04DdPnCKV31h//jnB8I05nMaxe3uYXbVmDOzidD6mZddc2iSXPKP5g7zMK9Lma
6M75Y8eyWnn7Ojbd12PPxBLTSA5CYhwyhTDFbvYPFnXGZrdB1BrlFRI1ImmLu5rIEoJr2DZWa53B
DG3SSGhnyz3puYSV0jg5HnIlE7FNUhxyjm/yGUbkPjWyGNd+eSmSbEn4wS9jXkZFHBQDdJ1J2v4N
fepjUtCnAAL/lmuhidBXfaKV4BB5O1ih/5OkeiBaOEJAjGI4DgX+8Q+JXQTTa8WV43rQ32MlqDKg
idDHJUDZ9/m/bEJcxoG2N0BBTY4qJrCt25yGsfwT/UMNmlShBWZW9tUJdaNFaT2QhYJBKWlCFm7a
+AxuBX6cG0NM/s9v2f7ey8O4iv4DzOCNCXHc0n30fdcskl6NUXRQZMD0QloJo6bKUPMyQb2s8uYB
xlOvT79wVcRnsh83RlVaNtMV7LzqB5+XmhRcS3JB16kWnaVuQD1S2WCj3V87A3N66SGDgy5N/G82
6ZTh373P9RHTeRfdveEAXOH1/fgzVJXK4+hxz8dMqo7iLIV9ekjQFO4COGGGPfHc7ErQGERmhA6C
GnFgETt82LnPOwx5lWFxZJ5AjGAbcGQT00EJbw1hzpJVqSqiMzUJKrhp97erhGgejdZmdaXZpsHy
T3WIgjJE4tAWkYEQQv8QK0h6pHxC9cIaqjpHQXJVPfjSVkKJAKKBrqYgf/Q4f0FaTVHGPTJZ9SzK
nR2f6w88BUYjZyGj0/58cUyvCx6YZolDNUxYngJbZbraswCypXR5Ic1LK5F30zEw6BStMPsNDLa2
oVaPbbFgFHQw5Y/oJ+zVmPGtG5alWEOGcgPGCCqstFWbcWbELoeIKY2hQGk1hZMbWmdMWcRvsNOG
3x2xGbbX8n/IZgOvHwC0JZx4OGwhEy2o8vw06RyQN3mNxkVgRl5IYG5ULce5WZN34niVEySSvX88
OmDUoCON/7BnsJnoIF3GVHQoO5g/pyVwtRXRbDyPP65Ai0x4HGV4M0AkbaW/QyYHPvlnGc7cD8oK
mtfFsBioNGrs0KQlVngNqc/DsJmVkUwvXrOBqbE9P1FuQLlcbZiWNMu5yzxP6HeSjahFJP6g/Sq/
7VL1CdgbX5D/wqiCqnt4dqx/2mOd64zSd09/BiAjCPY7v5iSg9/D6niOvnHELSb7hXKMiTcAUAAU
jq3GKlWOnbA0dCp2WtAmbvI1zdDDVtFVeNEq+iwxKCqoxuM1dTyzI8lUZ0LpeTy6R/iHPF1fi9oT
C8ExP+Al4GvxHsXNYOMiolu7c+KHK6/EIz8xi7zlUQGRX1YP4IoA6ysY/6+CymK7Ng33tmJE6oio
aKO6rT0BFE9vIY/IOUpd603rwWl/V8wieTyi/1dZaZXlw6hu6DDuTypQ6ueY1kj8HXMjRI/rFfIe
8DlpgEXrxS4A7oRCVl+pBduaikxC6fuN9oyyILTk+LAMAP+WtcjybRi4abuKLizz9eUZptu6R6eE
A1CpNApr+qdxBEDNdfbkJKughVQlf+5Cgx9C6NfNh1pr3wStgvAWv4XAVbSOqGsAv9gp3kcLNttF
3Dp+UqiX5MBw6hxftB0978wmLmxz6izK5YuLIaA3YYUu+y6OWyj1VtgS3iodoQmtQpF67RzmcRVQ
9WdbmQjAm9CadMOqCx9WLsXfiq+HHJVTo8Cq84rl71hxw+CT3lZuJ62eTTtSZC/FSKUIHvYoyF92
9FO0L7h8OWzV2Iw4vksCNcVjPxU+/q0oAr1Iafk1QrryxZ4rSJXDcpjEDPqXcFEyPWW6sHdUf1wg
/rHnvh2crARCH5DynwIvGOpcLsg+l7oPSOAoYJGE3ovlX7xRSN7NMjsQah8l+rnWDfZNYCqLQVms
ZBsAM7HkaIlpyu8PVqyQ9ouUWMwrsSFxpn/jyVBcElcMursLJt62fCSwdZQXCKQOFQR1dC+XengQ
SF5o0u9hJSb4ffBbJqE76hGSpYcZW7xlq9T+Eo/PqpB6mYCdh1ZMKHZt3RUSY3qUi4uOSth2t9Md
+m7x47+BFo+D3NXwEZdT29YWG2KpVXl4bHTlSoDGYafdhQKJam2rmwlCm97UNU4zlBkb1KxJ0t1E
e+k4Y8R09ft2JicbAE+ZsAeOSHEpdBr1ZS6vuApy+H6lzISTa0nghxiAJnqagudV9DDE/CFub24Z
9QzHUM4/AeAv3YahwgqbDsyUyOiqkfZpAnSnM334cnIK0mDxX6BEak8sRmfXCWfe54njfUO9jKGc
5DpU/20FfzFrBn91KsmdgvSCzwyqwHyalWoYpOk91+4vC80vVKocam/ka5NjvSOa/VjARKE9qEQZ
/ANnqAV0Fhh6loCmW5Vfv097uW+DvgZ/gcpNFGP7OYffzyNvipefRI2mjWYxSaE76qRhBmd8vOMw
dzFklPrXzx8DA77zmfDmJdSyCrHh2Ea6OqmUYKiFJxgMUM0v6BoUsiLagnYPr7fiHFk/KE+PRo0n
hYA38pvskc2/YLMCy8Rc/CMXmMYWGEqdFXMJg2AC+ihBELYsYQwcgE3HFK6vrBrU503Eq6LjQJNC
2B8QeYkg0aaWRWHovs6N8r5ZN/QOckogEOT78i6N1mLNXwT3eqyvb43mca5c/Aq/5mmmjDu0dUqz
HYynVzv4hB1zUuG0fhpnNkSqmnBwfmMXiBdIZJxoUE39E/DKa1R6IFpN+11UUDODDAE6ZLQhWSCo
nEyfojazMqPO2fl9FshmkptbQNLqOX+YGBGkoCU4i4stJwwlMgWSdWnUSPSlgH6ZexO/OQCYZHJa
LVqtYQ7bxIqqUNFTxmvXgzgEMSc42qBDgZ6UgoY0Rr7Ji0AuadQ2STrLyAp1YGCjl55ksMCeV/ry
iEDQPS7DpI0QfG8h3gBVLtVeroM2rvao9K2/wsOOZCYcHYgWmXU2j8BeFaEKN9SsPNz3v23BJ8Pk
FJk5y0sqLbXxJ3iqMbSlulpGaO3UwHULC24VNrIg0tV0xOS338jpfCgLrhpgyzv6z0wBroaS28VB
4IFG6dqSfw5W1wxgxKDqA7LNyriNKMm4y+HfxvQUPS39y1VOB6EUcJUs6JuWn7x5xHTxYOnykerL
/khgv6cdp5deUTQU+kFQwhhidIaJAlhxPFpCY9PDNG9qhL5l5ag8rF0OZv+CdoNYcN6V31XIx4WV
iVkOCLKck0VCMHO+Mm2s4usCyBHWsiuvSOdfSp9hn7heSIAPU+jm/u8Luhs5tC0DoZsKHa5MZYvg
SU0fYbKk4EbBj5iTB46qlnEfNGa9oYbt1ANwfA3cdPiL2qBJ9TSnmMqtbeBRsjbtPckHklm6utch
nrg+9o3j6NeysTbp2inY+qc+87wVOorptAS+BEbfnQY64pk5oj3iPh9sjMYl50aIIOn10KYBBIXz
pDjxllXWuGzZaWDpkdaIJwFGJBTJfH8Iw7EhEuwr/cqocRwpJbIxk1p8N5HahcxnVg42XgzPrbUV
kjYqHEZLq7a/RouC25BgZcPThS7SABJ6Z257vR2Phzd0fQrcECb1koCji53aq2xu4RBFyCCZL4xQ
fPIF081k4qa13twMmRrPpkb96Ub2DxBm8x7haq/DWx8bB0KwBx07CiVdK8lb4Ha08Tgou0YXk9Nz
qj+4bOr0xV81G95QSpv7WVNV1d1V2yOv5lxcXs9YGvr27tiwc6ffsGkGO9rgCgDX50ED44CNnUYW
MXeZOZGMfFDGxEUJ3tTwLNEhtJ/jFpu+PqdrKhYK/zqHxWUP3ENh62OS8ipPiv8a5h9I53RwkelK
IJw0LEyeBrpNQoqcONxoZsOrTmG9FcggX5lxz/x7OEEeky/4ffzNa/ENO5Zu+5f2eHUZ1ymMnmgG
MFXVabUjAgf783+n1+KQBg4Tq3XW6M5pcnZotcpEn28ZOhvpPOt9bKoc8dn5vTD7raPK7ittw6xi
Okbc4idCiOeDOwanLxoPmq43fDx1emNl7cDleIgZCYidOiVRLOH9eykBAgaTtC7vxUpKLXE3qvhJ
qHl8NeQtX9W7fDxPr8PES05MrK0pHlupPEs/vxH01Y0qzIPlf8CfV67PDngqv7SyqPtG7tNh9XtG
RZYKwTqqHnIlId8zSMF5Gz9P3LhnMP3oPm8iIc1jS9c6X/dVXdWXoe9t/1QvN9lc8b9Zkm04dDpG
SiIvoGLvEmu6DsjjI8/fweFByKBfgct2OtY8/y1c8PvtG32VBrXDVSacgi4BP+n9sz6EfXqoslIR
aA6uY1RvTrN5k7P1NETwbvN2zC3AvxBAeDAMgfF91VNRb/rZKCaf1BwWBhfeKpAIaPYQLV/fuxAL
1ROrUR6ThJxTekAwRWMImGFwmvAC2Uo+E4igFFsOSF+7PuMZRPK1FvtuuwANuX4vs4H1y48TK7Fp
2PVdZRJjXB4cwqfu/wl0Lp9oKZojaqOfYFodrzXoex65Sq0OyaaGWrWkUAxBGaJQ8ntQpUT+JP6L
qq7Iw9s4UOqgV64TO61+igQaQUkLrrd4eU6JUB3yk2HnjFBrUUs+SK0QGOEV4ZHc8uvtUpt9NBCa
M4PZbWeQINwzMpNONwxfdqVxX+7vVGnLJ+srG7oolkvm+LrP6abfdS6rs+cd8zh0xeA/Pjd1Pn4o
QBwkj8Cp5R5N7frIYMP1LBJi77l4vsHqJkR6bgu+BYt5+K4DOLmYx1cOXhQXdIPrafs6kk82tRDu
HjsIGKW1HjX48+kBCqL0SRCVxqVpYYKRW0KkojztWwNlLROGK/vvJ6kBYd6c/Yt83SSeTakMO/zA
8O6OIJJ0ULmKo2NPT0obndQxHAj1Pppm947m257cPguspHy5C8+jBvgOWLMvcYtPIh3xbMncCbY0
gnxMqRWQDa3ZiGvNiuh+LwmWqayS9toawbVRr7IZAPB3RSKyzpnEA/2iBYP/D+LVFU0d+xTPEL9+
PMz7gUdt4UXoZ86DGnJ/nlnfI+4qZER2EQ1EeQ/AYxtV1i31lVfe/KkB1nRHOeSMMc0Z4lKTUA3G
dcFSTbfd9yqa6j8BV8KUoff9w8VIjDDyzFEse5I5HBPwDwb0oNK/v2B2pm0VM13vlXBq34x1unlW
ctFbvCfkwjBF/MkkeZwRUh85yS4SPF9CM2aU83pOtrKU7pVTjfo3MVDU6Oils+FHIzs9zx8YOvZR
rXq8EsFIjrBHDEBv3nChgEbRE8bR+nlFjcAFiWuHeRiHjYulpP1PXNrYbdNeo1T7mNy0qoWj5h1D
ybeXYo6cy8vcXLktsLrXSCXVJhY/rhFVYUnPfOX2FQM8GnkFBZ5qloRgpc7aBd0aZY8mPgSi+iGB
kyKFnYIVnidHeAPQzyshInOGXAY73+22xs3gETivEIoaSf2zfRjHNwYdGp5Qs6dhuubsjKhSxzUQ
08QYlquS9W3cviywA7yg9A8/l3nr8oJk7+Mnjfbc5v/U5JYHfepR97EQ4KIltxqjIhFsjlgX7x5n
BowyzCF9Lqqcx8xyD/drqRgnReQ5jg1jziudeXqwub0opXyL3d05LoeOrYUVJsYzASJdVwrBo1K8
V5kCYrh2Nkqv1oLhbKVxowfr2KzKp4F2DNMsaVMWi8qo++OlP6qEj4+JVHWWRzDrT1A3apnmoqdk
Ti+0+1FEluHCVSoQ1zKRSWuiAk6UhtBwl0X3p4j7twkA7yxPGiujrFfBB45qJ2o3QDtT9w8f64+Q
rZ4staIa1juFVm/YI0373TXqRHC3i83svUynZ4UjpcKlVqGu+bcqM6boQ1U5mBitKvyZYPGdiT0Y
sTX6LtDHw4sLM0YWmG0fy4UcRL7ReaspPnhftBK13rV9uAgOPsPKu/O83naHOj47hfoSvWniIBfu
3/Nbr5/cJ1rhWSDT5AePZyuAdXqZy9O7anQHESj/yagyj4GG6ZNeJwKdQYMLaTePYckZ6Vh+UjHH
aR1YfJbjDX6q6uXqFuMvSPhuoVVYfkiAyjF9+ecDEyeBNDjH6PNFslOuk6li2jhBPoT2GQTmHie0
WynwVUEfMCPPZmlvYS9JlLoMa032lAcM9pxFPQ4UIdURsjDA7ds/L4rGKpJcjJ6ScffR+UIbirXZ
54FyVyRyINTBgfKl15CSvySzJyEN1nE/1fXbgBPe40xcrchir3pBVCCVMbe9ZwUkAQdbhXR5U33V
OvSECeBLU3ag0Hd4orj6sWdJHI7mb2/qJvwT4RXMEycUkaqgGVe7OZGnQlF5ljwhMqKvKY0+cLrw
Oss25A1GbTITBwkoqxywCgY7ZwoIArbLRBCLGodYsk25+kiUMq02J8bI1ZJaJPpugKz/lhvxhqId
OKkdZae6U17PuSmcXhk5LAn1zOqaA7S9i2Ve+TXLAn2MREFulZ4XI6t9aAt13QlBwlVZpMNhmWGc
cFF78Qruzvarsk/qlm5Z7WTCUS3AFtC4ViwIZOvqDlD6eg4p7hKdIDWsyEgS1tt6fkucPF4QZSbR
5wcpuxYJVF8Ped6ErTg/TjvsLteSvq0whc/KkSLIKlltN2k06zx28R+aiB3gsOQaBinrO+zn5ask
1zBOC71hAXehAykO2zTnKlIVX1uTaFoERHmoltwzYnNPA11PhEVh8SK6CXy9J2WPQnLAto1O0K7l
AtpgZgVul7WN0Q+onV6+p8nk8InQVA4rSfdfPbShcFjruEDjN/X06JtGc6JzF6GzAP4PoYVAEvZ4
Pmh5ge7ST+Lg/VK0D1xGH8f6tvAWC4SkGZfYbw0/AlhsjoSxvkHbQx/Ydw7Dwn5qsj9hY33OC5AM
s1RJTkGGkLdquBTQtzpjXL3TImvfG+yziFKuQe8QZyu0DYnW6/SnzUlWPR8670ft8AzmiP1LoLNw
8J2viKVxeMD2PQvixJCQUvV3yTvu9Q/Z4mjapPXQrGyxESZ95YtUxqvTB84NHx8ebHcDduCslstW
pgNjSy+5OwerZDQFZ74ybRH3aPv7dNkALQ/kp0jrZfN9Zmywa64v6GdYDYWpZRBWLyneWk5dZhbS
uu3f2zvKY/L1TIkUFqD2oe9XA+Xh44xyDiA9fj4tTIMzaJiRaAaJLoJ65Ps4ZnFaui+Juxv1YiWZ
dsRZoH9WrXbBiFbpJ4RNk+sM7O8bU75ZRxy290BJ34FSm151PqeWDSOKJhgPAaRI3a8icavWOx4m
v40RavyOoc7dbO4PYq2Y7O5MpGWPXoeHlelK0iPkMjyuCSDPO5BtVgEGBEX+oRLpCiN2L85AxHXu
U/1zta2kolkmqwIJSQfIRIoXWsWsz0QL5QGRh/zUdtoZFn2qbTfmer0lU5tmLTILS/gSUbSEZXCT
OkDvUvVsIR0qsaLvO6peqPRD3qre3/TJ6/hPUFy6f9xEsIbDNe01vTWJK2a01DhhMtZoX2GIoJHv
Ioq9JexKKpSzQ7eX4zAWNtaPxklSKrSgZt8thYLkU81xurJp/c6uRDxtQwFLRtQVg7aa/v3G/7um
PhJv5WHfQO9cJBNAz/GYaa02DuMV7K8QeleRU6UrY0aztV+xO5CeFVvMR5wqH/soSQBNelj9oiNY
/Ry3yAGNz8PZ3nut0uq6nQ0XDnsuu7A5JXig4BMmJ8otQ4Xp/8J7BGSVjhR4dLg2xWbWl0ao2PTB
x0eAXlhRNnxEOofdkYWOTMAkOG/AY/nyObl4qWdErBTPQ2YbCd4KUe5oiWZDh4GtESSmiBoy1yiw
jwN4B+vGp0HljPpXVQShC7DBusYQqJCr0DKrEsXSdiJ+EDQt5YOtj/iXVyhCG8lGxAoYDFL70pt0
oPFDhVD8jukjZgpgjF/SLWGUC/SR4i0JuUMWSsjkH1wCtMEa0ncb/bgREqaistUpIyl6PLYC7DU8
Qvrxg4Bm87a5f35ANwsuSvxaGosqKBiYMNt3lL02HJziuwwf4NpedvzAFF6u0Sz4DNM94BXjKMh2
cRBL+QFRPV9RzLNZrojKnNP0GhGDuNY3TKaEzFNR1dL1HJV96PUlNPF0fHAuOwdbvIrHy2YtGAuT
CzoKYmiqOIlIGFSZTG1JHuNHwB/x9VzZQ4rNvTcB/tGxu9LtvaIrKh/wFRmYeQyqtgGI/pMwroNg
PgowdrZl2FUdH6wsUh8hkJpcQ6o3fuMymui2Xu1OpTpKitpXI2nih0FITNopLAxKH7jzuWW1x7Wv
Mi/v0FLDVuJFxYAHkzXGcGhdhJO6f98pN26PtvWrXKr81r/JJuR+p54ik6S9PC+5PSIYxgLloTC0
tNr8solEfH0BBNxjtK0dSE8ZakdubFNLaORw1mGMI9lrYBg1429vtWSQ9wRrKSGqRiSeF6rDR+ug
LxxPjF4+Cjzo22r8yuOoBAlG/YIJq0JnZQsazrFiprj/PhAWDWzsYW351J2v7nvFztlPwOOp5Bti
um8olYeIos+T1ZxFIYTQbyBMrr0O8bojohMJzH3H0mRQpgBZBwgvgrKKwo8/qMrM5p/9FXEvhEjm
+Tr2z6BlliFJ+IC31Fx68eLMmKnwiHZM3cDNEoyL1tA8TcAQXlgmTFr8ph3sIrZepzJdRJh9kx/y
3SybuLXpAHMbtCziJhk55NfRyeWbghOVkxEQXq0w2POtizULPlGp/JjF4xQZLSbgXhfVCuZleRzA
+1EDxC0Qu9GjySi/kYyEO8+QQfX3ideR4zE+U4BPyDWpT0oT1lLcMNzxPHNDeOJTAt35dNR7rn9p
v1QQQz1h6rSExoFRFSJqJeSdRgUq7Br2zAysPYyJDZlrr4rW0jSCMAvHHG3H2wBePMPJl1ILaHNT
8YCwl142XjGu89YoF4D8OTZQfKarHV7oqCyK3iY4xRmYETJK6Cum5oxNvle99WYUKcb4oW+mz3Ax
cZVRaOEWj8n9gaUdqK+pu3ZJ1VDzRClepHsvddKA1J0rwmDetQJOrTZT722bUQXVnZh+h0mu60HY
K5q7oVxQpnupqvhecT3VPt7wnFtNlfHNMJMkKOT2iZXX16/RXD5TB3uCC7/c4ZM9o1vRrGvcEiik
SGKzKD9ZWOeb+MOMWpxcvziaamJeqLY6dlL2oNSpT+toYByawW3sEAKNx109fGki1C9rNb9bF0Pq
+fW+QmNk+5j+vfX26skYBnGiU1wHuEMo7FdKGp5ftY3hnya9DVGGvhkMkSaUbeQKcu1oFqqhCtZy
ylyKYebjUuMwhz4tVCSiKptf2sLEWhq+Pmhfdbt2RL+gz+Hdh3YHj7i4NeIh6Kx075Wo2/3sVxVN
ePT78i6gW4g1WgodeswsszDrbwwFK9W5S/H+iIF6lmtk+zJulLr+Z9tKgEctd8H72NecS0cSaueB
nhQ3XoY/DnRLQseoBIIgXqqyz6u4bEgaFmqobEhUPVbM8H7D9SBXfPat0hBdRPt9V5CSpsQBNviB
a4/D8WEzIZ9cPKXUzfbA9kg49L90a5SH8CeFrJFtG9heOOQq67pgzyzyvMMhf462fQ0Asewfcq8z
F1dhPbvRDoFkK5sfUx1wZdFYrhS+otNMMc48PIxf/sDSUUMX9kiGwR+6STUnuAZFOoMP7r2hDWCr
QgejjttC9Cmjh0PSOKU44eI3FpeTXGCnGu6oWtxYJathyqm6cH7cwWCtFx4NjelLJYlxfrd+lye6
thqZyhEFirnGT984I8b/ZctYDuDg/zle44kyJzq58txBryYSTgA0OkdHpqTR7Bpvn7p2bRIDHUed
slFGjSF1+kgdNXbFSIhfycL4NwD21MfFTBlDhn1x6HbdGBob4oHDOrsbKq7Jx6oS+C+96kpuSq/L
i5bAIp/IEEfUAU9xIew+zhV3yBbwLQYqk7F00jiE0fcZo2djN01lax0lkU08dU73uqogYbimZBXE
wtdZ+BNH3vlIC/Hsyf6ytqCq3GtBq3+1L04M+5sX67LylL4a5QkgH7kxs3DsSns+DOolpk0RExxP
IU9zloloCjLiW5vOQJLZ9nvXlzaYfaIpcHooL9HjEfGDDQytmnzbOjlbsZICKIFVZO64i6nYyLcK
XjKCqK9rls/olkshyuX5r8qW/l7m9PCygAeU/3QBkj8xD1gKkCX59cC6OD55AEgtEgUEtVQt1Hy8
YHnB8NMoRnRppjw98XgrBr8iGiYcBHbn+7t47kxqzRCeS+DijTWYfp+xUlz1kdxJ13nQmrw5QWWD
K6mOvUSX4sjqfSHJ6Q5Wfvmlp3LiKlKnzyjwnh4MU9iHt0Xl1BEAkm2Yxe9FhayOCsivTTL3ifLH
vteuNcnsr5CGk1vIMNumOd22ZoGoSHVEOgndmtrzbqc1WftvOkZMG3j7HDMOdDw/DWfOJACUKe8X
5IgccUI8MgpwJxTiCy+Ykcjjr6CxI2yzfPE9jq75zZnnnPcpqNnBh7ZJfRIXUsce3HF7Fk7hV5fW
8JYY/2Ndg/fif+m4qW5D5gvyGDi6uO5IUNtVKem6YVEedopxuuaym8mzizJIvlnbolU7wOyXj6R9
h97xHdmUYzbA1tAy8AhTiS0STJtZEWDJA1MjdDKDRc1ia2ZxWXhVLgTwkShvuAXCOUqJll34AEjp
gSWCwq6rk389OuCvN0SF7epEqlXBBWr0DobG0WbWZoaMlSE+ChYggIxVZgpHJE6tXroSjzAK/Mig
+PyyHLSpRPBsOolPaUFTiGg+CioVMMuvjXXXDapQoEsh7VldvLZCSvGFuD5SDBmURY/Xi0+pPJ5V
UpL3K2Uhvmxk5f6IUHbtwjp2iV4pfqW25JkP+Uz5P7adlfSBnw9us40hwLKFdCn1QtIzbTquncdG
6FvHRiAwrIeqVgSaWETy6N2o+kzMtt7Bs7t8HoI6CPfcAbkYR5D9VgyiZ77lRdsWEAYGXMLEe3sp
bVbjhysegWqdEnIi3WCgslPYuhJXDcUVpFjRcVQSJw4tIKoPLfWAVOQ9qhQeZtSkn5QCwv0KS028
HKRYoo1XwrP0hjhG8TYFZRxgeEWGIcKyi6uJKl13BHWpoXB1+83KKosivEBX4ivK5CW1+36dpDWJ
u2xduREAwnDH1cwdEIBu0GkE3Ejm3nyuEIxsnayhWPkTL46YdvHJkoYgJmTPZUd8HVHe6KEg+Tbt
ew66w3GPtKWdxyXJ/IgtaAyAzA/08CG+1NHtoqZs9ni+wHrj8I386cMXMryncUDXei33KFtNyvPs
CTxsU7CoN2EbZLIFUX3DeAXSFBQKn2cx4ipd6exJi9aevy0q7YPN8Xuy6i6uTHoqxr8Cl4DoCvAo
Jit1Xi6hsT/D37Xn0MHIjZhzq2R92i6AfLZyZRR3FFJ25kwvMaIMS/al2D78NTZTF1yUAVLc8PRC
ieTS9mpTe5NEXHIsEvHWAst1Ng+C8vOUEH+0s7962PrQBkZFjZqARDNU9VSKiJLBxS+0u/QlykeK
EeK2j57XhM+Wqc3SitRTp1SD0rJo1gkaoMtiylP3lQCpcYQvMnlsKV6JVnylUGy2vOI+cyMqrLlG
BH4ZnDMiwniY/UZZ+9Qw5+Fra4mnCHifnQeeqms+SW+LraWHoeRgFBlwMB9OLLjmMts1ze2cvwdu
sxuJSKZC81DEPXQi3X1Yo7QnzirhxLzxeeL9Q4qzerMkIDLG5me0augn4baNNi5XyvVj75DYU8IJ
MZYp0LJ3SUEQiPNaO7j+SeHtpqIrUfItbykWOCs8H/O5XsPhn6XaGiPzqTZP4zHYBr5FLGPwZxUB
71+hlsSkNOgUCXauzigcn+nynXtGgUULZJGRUrEz0XisW6HMNBvKrQk+7useb4Jgboix/Lg9/YNy
N7Actsb3W29Qqvj+HU75K1lg2nQH4QUzRBwQml2WXn/NeTHeasVmoK3rAaolDkah4fjeCFkQHXo4
1TlsZx23vKKjFT4T1NJvaO0/oGPNNkgWNq687/5s5p28aUZPA9EkoWobkYdKCPepic8dqQwu01XT
XxApJoCjFetKOQHE2lGfXqOuqy/EK5z64QMocaxt7pdIuVvU9oC6H1/bYnh5fLeZzzEut9OuTRpB
0Cm4WJSX9ovNZq28nqn0MApvZluWaMUpWuU0oFV/CRNytdJKop9ibJKmeIf5/jYezs7zfqjOFbRx
MWW6FlqAaMJPakQI4/wVxIXUlU4+it6GIGXm8wgm1w16VsfYkdVcYJ3E1OFkDHf0UI+7025f1QgS
1TxhEzeud0xv+vqVb/gzTct6ZUOv6xi/PspSUU4TciAWio25umJZS7BPC8/Mwg7GSE79ox3uttDT
g0/l/fP97S2ipVeOAQEAbneiOqU3PLWwmPZCFku92wrwXQvPUE6FDz05DfF8O/AHHNj5Bahztigt
f+tucgIac9KyhL9PtejXmIYc16RUDFRg8RSGfzBBKjTVh1Z+N0KVQqz+VEYGqdEapjiPuBvFn0XJ
uP2HwnzVm8zbowY442OtXrJYOj0QNOyt43i5/+RCqFPCerdSPrTdiyBaIKCWteAvk8SlwpZaDkWS
vmHNxbab0sfOfKE9KWlPQAv5stzfgFQhnbdG87vftQsCh7/YKyUhH+VKIdbsfVvxzdlGU9cXrB6I
MmV+/g0TOYtkwLU277rj5UogDzYcclWqjLDfomnVtifcqhILBPEHYRnBsXuDp311vT/108bY7uP1
2auB5KaOslsYnS4Ly+RCeFAkxa7HGZy60B2j1tG1GMh2tBDnJasMu8Sk8mxMTB37igTj2eaD/oZN
6K9Ktzob6ZnFf0nMxwjIBdHAG8LindB0GTtC9LiL/9IHDUN984spgW+Jnx+p8FmaJmuarjaelFzw
W4nz/sqb5aAVnwA2WpxZvO0W9g907gxWSYSr9TblS69xPqEr0ahasMvHP9wXqq+LssbPUdfqDMsH
9j1c+Wi0VJUSQfUnSSYC6mRfAPU4E6JcJvgHDN9lIHeSM4QC6K6pCeoaL6bbUG3g1EGYn/L4WdLq
jEVbyTSBczZHNVLTgy2fhraO7xRsfuoxiPTlA4E6qQmjQkSgNLHFbjK8FkI4N18Kg+TQx78zRWoO
jsEvY1TUC6G6MoY8GGM1FaV86gs0LUmRmPWLdWvxVrhvJ0u43Lek7Q57w7BeBZEx+W4kTRrPS97d
w650aR4U8ThaRyFacSJCKiMEgeLKyQZPB/KpZioUSBfkyRNSvlan7690sWEMOYtGozWbqJwFRbAM
OypVAG5ryVIvohLvz/+4XlhKk4xq9AbQE6Co7UIpvxjFfUImXU35bR3aPbsKMUGYgEUbDqlJmSTq
1ZnWtpv+nPFhk1MLZQcgNs67+KETAmjoWZ44pwl0959aKIE+p7h1yKbyNvCs1hKqDruKe76RLz/4
1JbSnWKXzRikT5pnsJ2pzhD/2X5h43p29tQkGenSRjpK2w06kxqVpIKnNjxtUJLCY9DoFgcFmLQg
N+f6H889PqRj3x9f96qlNEADMpCOR9q4Ah3Ud3tZcNwhWr661Ok3Z41L5tmenrzCn4ZVX4eJyGRb
ltUkzQcu2dMc08IsveHciwv2yhErw0cb2WcJH9k28qa1ucveG62vesN6Hm6tQdfhQkynYANGEKL4
s55g6/DD4g9ta6nj/+ZU3ZfNBOT3w0Uespm6XKHBzsfgIf3UEnhXwXXXWaLITmuYpDvyLi6spAxH
AKOA4j8jugmqBiQSN+yOvLmw9paTrad45RtDgJzeAzpy+oqkiA/w9JFAY/UmMdjm5Q/GA9xTlbsG
ueuM9Of9WtLy72nURK4l6NmRN3AE5BfLpnxN/zUQd8aJDWrsPovNpOh2oGrEhBOVn0jsE+o6kYBN
AjzEIksdiv0pbC86YngLyrXk9B/oujxO3/t+7r8mN3dXYdBlVCXJLhRzMS4rlxSmjDjX3w6Oy/62
SR4Ny5njUM8yvzSNT1R5+ZDuc4SPV+FZsqVQxh+vU+1KvROdr3PILWt9eX/c2p5Cmbt2z6wNGRCL
cJyIoBe+r1UBMp61sZN5HwFk4KwJczwWyQkx8Qd34EkSJNlU7jQ6VJ8O0B3CkXhr20Ehh9q+1BHW
fq7sDH42uZ8Qk7ZXgTEZpuRauUbY4zKBzXJVb9hMnRYfCodc8PQGMSPjh8sGuCkXIqaK3nhFVLlx
/JvoVXcrDhnjeBK8kPVCXicO338fL7o0+98uhPdrbmHzWN48Zj6QIteuO57lzH1NXrp2l5eba0wj
F9j+VjjEB6BYolMEg+ie4gO89SnwqXzl+rgEvrFMjKfn7LjBDXHxssBCFe+RgTlMu3dq1ZT9SFqu
HTx22Fh1gYx/2mfVurh+W7dd3hQ/NVEfqf0Y0eBy9AQFhnd/tStDNVQGayquQ9+EsZGoJwl+Vcrd
Cc5Ju+0qZZiWgF1LLygW4yez6oF35JLYOamLrXKgNorRv+m+AWhk3SQwZlD1+3dD7PHpCGd2Ci6K
mFl7uaGooMSD/m4PqMClK3Z6xBWSs0tdyEaAujBGXk2KMF5OtjCVIYFQ8oRW25MjTxEixBoXesOi
X5AGXq3uxyM4VpjvqnWqbwBPIdryc6GxIyaZDIYoh3vAmPMZk5HYIaBtTqrk3DO1KX6kRXZzrJMp
A79pLSQn+itTxm8IMXoZ7ecOxhik74ctzLD+Oa1Xu6iw6J+fOL16xDllhzGyhdv74JgpJ28aFJP+
bPQHH/Z53CDEKN0aHV/6RylUDESsrrorWPNaAQ1vMJkmbzlEnzCmtHFetXfys8bJ0ac/gXd+4iyz
2WIYGjFpPWIyjvcXjJVk1Cv+kaAayOddgtf6N99w+iyYP9s79YEMs1OYizbEwIv8TwTp4D5MTaTM
JRj6mnlI8/RLLjR/Ym+GSs/1f35KSRFt39HgksWlnjCC+tytNKMfWuZSH7wtnxETNYy7h7UhqNlB
2h2RFddzzhG1efs4r1eteD0qEWRxsBUd/5Ooh+07SLOwLBQVxMIQhWxkb2+sBHWAy8hMOOOmsm4v
2e57RQCE35Q35uaxFyFYeGTVaSyFLS6pdy6UolxXsr5KsD/QMaR2w+iOdXf5N09Z19qx68cOM067
8PPBVQqI1nMgvYiorGrhi5rUC5y50DktfJTvwgdHCad7JPaadOjOFGtR1xXEe19p96hCpD3cN0K+
93A/hiPxc5b9LDiZ9DASKWuuPtzngeUir/dNrmIq7rvTwevo1EFjAlEZlN+BXfUvQ+nYE5k8qKMd
4q81saIIuheS17MSHPXD8Ye3a/o1FtM0Sw5jeLfrEiPDGgjEINtKe9axZBUynctOB5y8/hOiXXIt
8udDh7hNfQRVf/AUa7JeQgDMgFuoIT9aVXSEV93TYU0GtCr4fb+Afhm3ZdiVIVyjqEvap1IKXRXW
dzxtI18WYP/pqgsau06YCsjJx/3ymCE93gm70989BNW91CspjBE5tSDEuh/d+KTWFyBFRZoEG+eq
39ZTOX1+MScbd8R0SFWQLravO+RQLqEy808nxKL7Bq37LRb5ccm+y+rpiy0H0Q0+gwSx5126ktW1
46MTYQhICF2iGjaXr2gUPb0Cl1kJ5mtOCgTbtBB3+lfkjJmh+uvhC6ApLefeDRx/+G9+bZDlmvJo
1/OeXVo2Jnt5C1m4EkPU9Lc0+BrJfStqmYNrej+FRTAImG/curmfowuAZ6A+gCHoAFlpknTD0Syt
QFruROpP/fjdacCLBePb4xCXJmCBaPfQ4u+O/wjKV5x8YMRKBflxJgpKft+NNN6p4v7UCAuaLnCs
1Eq2sGo3iVjiDSh7DnME4uFSQxujDgGqSSyWsMR1gFeIm9hTRgxql0cKpFOatx6YC8QVxCYn46XW
ewrDY0+z5ufS3VqzqQtAsdbMcpmkz1zUrC9D6wmPkEvBZh2RRw6O1cXcdDjpuZVTfpuKcC2tNkHz
2U/qNge8TYjl8LAMG0YbmxI1FTfwgRlLeNinGKz4fU5+WlH+EcwvJd9pOvocTrKmIB36nvLAQIfb
SBYjsU0jzh/36ZvakyCswi5IM2/V/iuCCry15rKY88yXeIuWZDnNb9ar4EP67qFzwxKWQ9Z5IbrM
iEOGd/808SVYx3IosD68txeIE0fkw4O0fURiKaBuaIAqFUXzcI8dg2f7CTu7dA97RaH2XGBtkVMB
jBycbRbNgjosqLTrm4lC3jSfeUkXOITSXKE2yVkOW7W0Dm+zlRwvmZhR36DZH8SL1tALsEaGP21A
mW91BqpCftDjZqRxHqmKFgsDbGywDOuycclDEQripSRjHhiLehpUDkwIV9xvC6SI4l/nG4sMUFXC
oLNC0Lrgpi9BC7t04LaVMkaw7bGMRc7Lha8pepfvBtgKPDDhZtUi6MdaEmumCcFRRBVJI0/cI5/B
Ll4+5XglydntYlfSZ3nrGWzum9avAAG+X45AmGKJED9w1VSc8KHIuLz4ixKHdLyxl/gAP6xANMip
sRnKRKIb/fdcxJSmrCOTjAn+xYXNTMK5cL4WnSkqDjlrey0wpiuM+kcwiA3x2NRA1hQ/cM++AhmM
XHCFyDAjajT+vUgIyLmOg7c87bxiVshscvUV+2ItVX9tSZAYZXezZMgWdQyNvtkPoZKJExce4SxI
qFJP555JfDt1OQwShsFD9gJgmEic0vTFFnZOAC2Gq7H1EZD/w48nbh4sMCXZ9YAGnhqnCjuUeCBG
ulzVG7u6vG9EWabynUGrteYa9ctTYEoNiszsTzhs2X69UeFAe2yCdKZfiUUYOMU6VYK7qsgqItyC
KcZWMMUbNm3br9YT+LJXW17e0lQ/nKWn0Dlo5ClojChreJe6W/CzbMPc9NdLL30ORovRqQWmtevL
N1zVvyGVkqy8nJCOZFWMQRwtcGUe6zo0b5G01zCvxjuebwD2+FmDFSTDO0Cj3iYiyYUEycSRZBBz
najYocek5MeVxwqovp6OsWePpFT8/tSv3VtzdhxBn6/oNHosAFmI82x4cMDvf6fOD02ltELnkOo3
YuIF72wDCbJUh0ncGsqt0MGezkN2yG+CWwvldquvLTDqOsdf7EmcetGJnvo4JA6+ZVJ9PKGMoBly
ctLhxQnvjS8Uy4/kd8PMuqyJSGiiju4We/QUbnSLJwPJlxTsGSSnujXq5NLFsmvwTo2xwcdKnDzD
ebuKjaQDnN1GY/QCJkaso+MbyDo28KEpzAWnSNNI05K/xHGLKEKXhMHrMufiNqAcVswVmoEqpGJi
4yAZ9mFvun4QEP2+NHvEmOml2JW0hnEoCx/mFE8GOyT7qODuMxD0XxTtMpek8RHH/gNyXQzftv0+
+cN8oD5kcHLS/d8hh9AUmZuxvj4ND/tgCCDUvcQlwwH8PzkQI1XVKFchcUfKGV+bqQ5QhV8mFRAI
+WVGACBye7q86+9sebR3axCVRZusLGWYmjGaVk/ngAKjYT+8btTdLrkx9VbiSz1V8Km3jCDgL6ME
Bf1523WMpLCRm1XIO4PtmhQYm+RrNOUaRsEU88+LSAewJ9SuIfZXjQmCZ4Ev0NCStxuThU8gqtJI
rRBIB6Bk/xWZXRRyxY5QJXZRKTEp7vcu4n9UBWZUNGdQ5IguFUtn6ufX0sBqet+xUAxCUZW5a5QN
FH804L6v+MbZYFroZ+WXcosdGmSyGr96g/LdI0PK+Wl/QErGOuK+avKtht6YlziUccOpOv/fzIYQ
CVGUzSlHFDzdy5EDU+X2bQiTP3s5EwzXO35CyhKgojvuSo7RCGkuGX7btd7gQBGJyNXwe8L9ndvg
NV2acxw0PqXPJgDF4icHXEf5IJGGvi91vx4+pMRgOo8mrrE72ZLWUFfzPHAO1hC+AEizeJ62UEr8
qSOQe0xMEDMeSMySYojp5foOX5o8Gd2oECwLxcNRyOBfzD4HbJhsJrwqhmVFfkI/oBTLuVNqZaUt
aZIyKRpH78vJvDRbomZtz36ellov2199VX+Ma4p5tsLIim13HUU6wUSWVL3MgZBENlDP3Cd1lDv2
i2xsnXJds1QCpwpvDEbOz5NwKv3OjK48kB9fxzVoHG3eLRT6q5vyGkpzm7Fk/gFvJJka8F9m/ZVf
dVhDxWQl28/Tz8svuTKbimVRxhupCuNrV9sedfpteeKAdnomdRct2pW5Msghca1wKVoI1GSWWg86
MJEdrlenxoXSgBz4bF14M2PglKPQlGjcLEkOip0KWwjxdH7cOUNjbQhYAI2SoKP0+u4i1eLF9rF1
KPDPUHaC5CoU+h8h4ESFPq/jxtsLK2FmtmjAUmKKaHc4pAYxwArClLyRILgwdhcMSoxH9mfVXFLY
Nq+rQyhYpQSizkaCZqwVISNsX2a5rg2zL/xOIE+l+Dd0ZJNdj//XNtysMjgyUra9h/SYaQ2t/JLK
O7qn6iEJ7lFBa0qLGMRXMERmhP9clcgvUv4NqU6vRDJHiyeL3Fqc+oGs7cnpcqsHzF+N298Ezw93
BJtHJMJx5AQKdFSO0Tt0YFJfSjY8fIjITqUf0FFVBnzeTismaH2PWzPYQGUtDeZ9aHixZfqjx3Co
9csEVdQdFi+SPG4wgxnrCei+5TOhUmtHpuiz6x7kQaKTnGLazVB5Mvzmfr6MtAjMRwxRrcBOxLXU
iG37QXO2Vqh7XcPO+qrzR1t32+OhAkOjEdlpgZIwIuXdFxERnEUsBaeRHcC/iwWZucfW5fH56v/t
Y4pAOQQwJgS3sq55+qNfuxr6010h/1T5UZSoVVPFReUOTeR65SdaFBWNG1PQuh/D2s3Jvu6Eh9F0
CQRSaTFXLAHvdl27psyagRbzEHXXbz63yalLe+DaCL6tKDB6WsCT/XottxoEnrJT5nJZmf1m+Qeq
gz3u/iCQ6q3cHCbZJTfz0kLfLdZfjzPCYNlwzO6N1WV8yWsvjM0WHJcUhd0CNAopfSntk0jBx2dV
3bY48bh3QKeF3pgUPV0drU0XFT2WaEzJ9+R+6yDEHZmAT/Pbdh1qQX3QZYMbD9MoQ9vUbp5MIeWB
5jZAIpDR4ph+IV3k+YAuWIoPDJviejnQwwqsa9HrrJJnWn7bqAMmo+aVz5r/cWnkJBcNlBqnfyow
cluGRmhm0ZJB25HKEYSz2GvqY1IWKB9XS90wTB1n0GjfYbZwu9yzJB4URXHV81hFBC9QEaSqVMfb
BhZTcKvy4xRH3cVGd8SUZ71GS/VuzuPGzUKWzWao859R+bPNHKDMp3a2mgv9B4WIXqY9xWNLgF6g
8oNj+eEjlH5i0zgHncHPVmJI0oytBMDOBSdHsSd678JlIWh8f1tmbLbvBDl5dZGu3mwklXd7WbDE
7wKZ8DZGz80UBVWyfxb2r0Jyx2ArsNXTSvbuwNiD5BmO5AJ5mSiO8A6/nXF38ioVsPQsWak7u0Lq
SGBM2EX/XqqVH8X2nvkSgsSGbVb4IsaqdmuQuL7dHvTtneH7a+cz/QOPiOSdXltM61N4hbWgDN1V
l9XRxUKKmBIWZpJ4CHDlDT2J73ArxykmWdM0Lvsz6aoeSM/k0pSl7WsTH4pVroyxJGE6lLJThuEm
MC5fPXfQB9Tlcs4YK4Sa/BQ/kMvN3jQzESk1cVphZkkSHBsvGQ74sYPWSdXKZ25TepOsdlHxNGy3
2fb159CMuPP1TWIdpwdeZfiWDsBkDuzk1pd3l3UJSnhK2ilVNT7cIqwUQ8cwRMPvafJ671djY1Es
2R6qLv/V5gJlxa92wT6ejdPpyBNWADgCYBijeMXyl9O0R7Dc3PZdORFPupdzVlc7VN2YPTHqvL8v
NHmSPKArO730lDM7IP91MSpAkpBgwxo0IX25NZcCh6BmFE4os+E0ZBsdYjPNDipz/4uh542czgnd
MYmE6djXEdIbV6cJCwAznk60mGIUUJWsbBhzfUh7vuybfxn3Q5zL35DxeTtzIB8RX8jID9M0WhVL
NdJd1SketCTUVPaAjqLKP+/qNxWazrQ9QjWnpn+AsQHJEA3kKTtPPiJvcdWzT561t5BSb13RRDp6
pXrDFBta6TXZHU37oGbvuuyIc5/9JN9/49tOmnFnOdRVOcIeeCeR0pRIEn4o9dDc2CsrfZNDBeVp
NOCpLR71+oTLqURUaIv9hfTMf6hSOon+3DiHtJcB/3h2Y2v3ZH5OR3LD3gSSr76rcHGRE/1xwB8g
a7MEk5L8nNDGHq2dM+SsER1Hv+XydV2R0Lb9Avo9RYlbc92aA8t9i6Zpv3/TEEgjDfpz0XCGOxsD
lJIIOKNNQ59HJCYqAoVKOnG0Z8iWh0uc4ipuVPeiOfOr+ZzobjhfMOV6TPlw305Rqz7Izmpy34k6
vEUkM2YEWq/QZKh4oVsE8SSRLf8z3vtw/Fq9aHy1IpyErOyh+SURJdh5umymgWskN5tC4vqQl7lD
Ee9VGyvH2WZK97Kvjci0eowOGcHHqaZz309w7Pbv1W0DTsWFGa+7rbRabYNLxuzk3U9uh/ncPLhB
wKYfKSdj9VmxPxIYqDuY4eDam9rbzBjecCB4bu8g/8wVmG6Ve2YM0XX5bOLaoOE8Fxk74e5Bd/iV
EErn73Op7qiI/nK7NWE1VJw4teTWWl3kFNyx6+FiXUQS6rIyM/nOMSkZf4lnL1hn8h2BoMHh6Ibt
FLVZ6g/r9m0ydGExuNPf6OoI51s1JCiI5VVxGtXvhXtpZLMba9xzYbtuBPVTrtzG+p/cFbvluYqS
c8+Yf58StqBgNwsP/wWzQLuohn31TDrpmG1o6gdg10RXd7TsBGjfqJ36SZWNqGOjgu64a41TCrtL
Av1JGT/eqRWOHovDwcan+TLVKcn4NAG8VIazNowqCABAdJG1WfiDGbgsQPlUzeXVjhvJzWMjKRk8
+UilCqKQCO1z7icc1qie0oJA7j2hAkdKBFv4L2l6dPYznL9GcKUO2AF8LNbs3I/agxtC16OyC5Ln
uDzAyRZw76m6VOlpIFCluPN5ClH/1oHWvKNCu/kpoqUqa6g96oVSm1hPXog2keV141wXLnUjpCD0
B0Ww71C/wmxg/COzLjsN5F3y0FPqLylDiTYklkzxQUBzZN4HXsDb+tE9AKwdfdMVctB5MnfRe4lF
CWwHFgwi7Xr0XHM9L6We0VzsRLXERrqXr1p2k0WoU4ngOh+SFz/aGSWxCwa9lYo2mnX26beX+TgQ
kah2meQx9yGO1zT8MIRm1MgMyZldR/NAajwlZCS6WLnfsXkcMgMT9DkMRS8H+RhhClF5FONg76j9
lT8cYPZXBD3dmCY4S4pSGiIR3WtkcGRrIVaL8B9+ObMi0k2akRsBGEgqP6lIO02RG2Zi5kkgWHye
Q0xwoqPcODzNyj68awr5Mjg7Iy8ZHOERI+bErvyLatPcDRuWcgtZsURoDPqMvBa/mrNSwQH1YZlY
Z9p7iXEV3ZdxKbGS+gHTxHUvv25lf0uAtA3Zbc8keCzSh5GPuCJZef+0JlyKtDbGquJDQ+ZIykMH
kyRjrcA72nWYEUgYOtuIu5lu1oEZZ8vZknlyZIMEsmuaD2r/D+BFiTuPBvDwLXYOii2yveWzChGn
RQKqjVC91IYw7meJxHV/SH9CsNBXJjvwXVZO6QTOtznBXA+vk4G6CoiFa16aoV+X57SVgGLot+++
DV3xBteydSN6CTxChACuwoIytIiCye1QAtvVKDNU2UwFaMTNz62iBDhHN6W2WAMAAFoIPbU1L+M9
xxFVM3xsLYb+c6DuFcAUTUiKMuCzNIzRANMySKw0jQS7jLGrk4Xo3YNQZZmqi6bZH710B16aB1xq
GZH8LBcOrK0Itguhh21d3Ye6HwyFF4VyxatGc9rorCq1kBX6X9y8YfHhfhz6WFKzJZOCyR6/YSLg
9VH1GiknvfjOmxL8pAPG6FzRvTUZ8T37I9YOYpuaYWYqg0xipSns/pAGhtKnfFNr1jc7ZLBaQOCf
GHixzAzbbDr8mjN7CfRQe8rY7A04YqwXtnbZeHv0FRr68X39PdTw2VtJRBPv+GMpbm0hnXcu/EQZ
I1xqpUaZAq3MDWNI4oSTRPRWT35nbAOjP68k0wIXzLgUn0tcmsf9gN1wJEvpkdHmsroRLcub/4yV
5bM7qVsdTDJSR7PWxuP+34EHVYEwsWvEtaUDFi0FZv6hfx9+UoWMd7cptV3opf1ZFbOrobs2ReaZ
SAFr9+ybQ4WMHi2uFQvWmr++6O9YB/WvTcpuimMa6GN/SDyMP0FWwfnl0jh3XCCXbCf6Ei9u0GU8
sUsuBTcDy2Bt1YpniiHTfyY3IZFOlYZU5MKagkggu3rKg9NlQCGJSzvuZpKvy4MuIKj5yyoyL5xj
6jh8PCQxbwvPNPkWucTcltwSCik46CwXPT74EbkrlhZX92w0U4upE4PT9lGKWsa25p9as3HK9bPN
pMrOzZxBE3vsHxG/uQDgLA3TsFdCY10C8JryiF+22aXsZlX0Kzae97G86k9hhhszvdMYnTMt84sh
u++EYXy1pzS417B8rrV0se7Q0D5wzaiskjox2TgVpBUlkKDjRk3uCPY9yjeAncDMULDwlB1imWYi
K7VdLByEnK8eV1La6wiLQro8+xrlho6jBP8SkYSWl86RBaOa23rLTUANuARPsSRhN7xwFpYx5CAi
u97ifugcKMmLQRRBo+E8DJMC6TBdkch6iQQg0mU6pupVAesaEaplsSOfTygwrbm+DRf2MMrqP0yk
xReMAze7EL0LDt3KXDE3CylbJxJpOOub5PdQudlyHxtaLpNTSj5jgOJBIT3TkWTFU7mbGXR7yrRp
rN8OEkmDTOgjWyIu1Rwd/8kyd+rhX/U8Hvm9IWmO47LWySB02ADzGCJtvpJcj/bFM/dYybzMJqB7
oguJC3LawMug1mjfktIFst1X0dGrTuz3WzpaIxhHiEOxDeaY4/C9D4mfMNS2sbrYOZFnqcQVQqJM
+W1IkuKP9F/b3CEszD8FHTSq/N/MFPS3p9Zo5zwxLFucMSBtKHEdKbePGO3HcG7UWmhg6XLQ6iYz
kzwRxy+Z2NRgFjcEJnxjnARw9JvVUzJdfTmFrdtK/cJCznKXqzvMuAnbwqdisoJYVpjr4AAPECUv
gZ7SZMVq3kZJCNS7qPuGuXBiJnNF5neI+2LVY1pv8qhCuTOr1rpuIQxfwOMh1uDM9ezNpkyjyfZt
crQIJfWW0w8/sYEvMN9cNEPSh29GHlciOqe/bjggPIKg18FBya77cH97v5NqVx05nQvS/ca7XYkG
IKkA4J22cH1xKIOtF+CatcvgCeqWO+I7WpbBq6CVzwZbaqYWYvWX6HwFfVs56bx14ItfmHYF7Aam
C/s4P2vr5AOTdr5BCwWofpoZJYksJ1N7ffWNcKpljFAcoz9jDsgpUxT+ebIm8BM5W/k+dNP0I1cn
PC7dnZRkKomT+A/uQLnhLsorL5wQ8jOPr89J8mMTjc4BIw33luyUDkVO+IWekHvSCHYHIWlYvfTs
658WHugc3krsPfOv4qZ0bbK+5ykS7f31r6OAeqIr9F5pJM/ulfb2cp3eZJV55zXn3frZkeUu0t2R
mtpAQpaskLjwvmjnOt7i7YndZ4qx66PEzsNrfsNmJkDtmm/uDtdBOZALbvpea8he0rla2CDct+xU
t9LUzSgrElgD5Z9+EX6CRGKEbCPLPwL4WJOpVDm8Ni5+DE3/JqlfmVgUjDzHXfFBnHtAbPFQQc00
g+ZbCZAWP6SJYwx0yAhKjeNoYtJPE1YAzbSNGCTZ9koekKN1mVeAxVbZiwCLcPVxpA5PHWYX5U5F
jajVAo8ZEiHekkTGomWesEVJWsGYShjclgmdfCsAhfoRIG1RF3ejIuiF/H7w0a8L92ChvQE0x1pU
McAWoSmiAiAwndsZZ8XGN2eXFE9cznpvX+lWjJFQB0lQRuRpLFrhR1BwpLLutSsqOWYEk/j+000W
nu1DKdw8NgdBPuuIKaZvNiGeaqnwhEwaL1JJS8jc4305E9NiHthcw6bSd+QhpOfsCkXfP8YLxMOP
zSIAgEpbFdemrXvVbnmDLsrtAtx8YiwOQyCde2vPCjfJz5VqAM5NTkzz/R5yjxEhuv95oTqbVjEd
sY24il9TBWMEWQZO3WUqf0RgPLam5nKkPRBU5sMpL/FW0r6vNcOdBEA7IPm0f+56Uk4s3U79SC/d
wihg3R0JGqUNypiy9bzoJMOIn5AxrJT1AXaNaKrooVtfQ4HkEuj3L1wEZuR5qSSZxkA3YyKJoNfG
eQaetxhjqm6LbYnx07QheEaDGT3pN6NOzR+mCa+n4yZVuft8BTQfQNfrHcM/qKpBwaRJiEj+TXFU
8wvzjICTg3M6tmYjeHhqq5ITHoBPL7U6xgr6rSgBw8vLODR6kUZDNfZdXM9HVTIJEXxjW5NwEK+S
4l+LjS6bGB12SNHByOtNbL0EI+6rJrMSfJ3hMTJap8rSn1RB+7rNVCLvW10WZoVBE94teKCDfUij
4AznlSGevZezF/mUYod4BIEljtHgr2vPLhJYucECd8CiEMGuY+y3cYlL99d/zrRRQmuFXX8Dw1he
Mp8amEzPyuJEkDjcNFpx5ilDHZLM3iesaiADyvvkvFPmupJgIuaSudH2NcG55qvjzTzmate10UwP
csSRFQeYs1lIuFzJnpNrVWq/oTwm6g96gR4gviRxfQYc0mhzbDeCqjeJFeiypCpQNRhndU9A3MPi
SK5oRZQrosPsn2/VlNCsud7d4MUCBcewLsrS5e02VmF58wMCDm43X5+7kCSpyQBTLoWM2ZjhF9eb
P5WU7eJkmrMXEsw8eNJF6BabYFPIO9XK9hMj1puPJPtvPqe+DDk7tdEX84vunoxDWv/ePEEFoWHT
PaHuHdn+pINVC58hOkZWDqANgfB0PmhEiTVKF84MX57rCBfFlnG/ISy9P0xCS0uTMOoWOOYVPj5n
uN62yVAckm0jOucRcuz+zhu5K46TVBIJCiKlbBoS/1+6rNhPdLO3xa7vRH3RNzY9aWHeCgEjfg5w
u6gehI5W8EAdhnxYklcPNVF5+OXbx52+pR7+gern0UfmJIV/2V6Dt7QFhPWBA+HveaEMQn3QEbtO
oNxrEDOxkvajZ1mSXdpyturkYpzQlB0uAG3UoPq50wVPbvuBAtJ8SYLgKcZZZ0U8HbyysnG1gRzU
tJXswt5Xu0/zQ6DJ1pmY3jK198pmky+iSBrIL9P1ImliHkx/hfBv00eegdjW53++qZ2RHBm5aMj4
5hXsVIluZPQU8hyQhtAW6Yjp6yn9tcfhg89k/+AJgUs9vUc+P/xrRMSxVjspAqGi/SSpHVb4FbIp
Gn6lEXwLUWl+9EIf/mTmULtWN8/gJXS3Bk5hqx7sLIaK4btYlQNwMOpySNJ7Ws/QzqA6ORUPN8L5
S7cQmLcS8aLnKG0DybsGWkFKSocJKyzIv7MLyriz6E9kQdmi3WpJ78yg6EP/A8g7Baxif+IBvtLi
qaHa2etXtQ8gTxaDvGzc7sYbZxSmgRPoUBtuIdErrI2W4Fz8eObXCN0DHsePi+R/2W6nH3Snmlzw
aY9O/1d2PA0ifMMwLnqV49CwVZmViLn28eTWzRXAUIJ2Eft9t756QErvyabe4vu3Y1LuHgj1nHAU
nh8PT/v13aNJUrTcwYXOEM/b5E4+mZsL0ATucvNwBhobJe/9W0EEUlXoHkjyXm66hacDdU2HWyCh
j5f+RWiAI9fPIkAo7CFyo0zZEV0NfAak9GrU2WuhLqqmFdEJeusFW1iBj9jCSuGsE91sud/vs6OJ
UphpYA9ujZ2UbNUv4oMsgiZhtm/rXospmeTxLlfHGlY24d7nBKPTHnfeo7924W7yZ9+4cVIsizjd
a1FeY0oUtKTsQFTERp69MtTtep/BOw/tuM69b5fNYRUigm0l4z+bnjNvRKf7kUW9x+dadrPoboPL
61SFyZkf8FkNLStSK3VlUeoOegPCp1f8FcNdXAUGlslcJQKxl9KiEO6dWhJv9gKdT5Yre4s3UTel
RPSox/er1Y+T0lwdmTXcHyzSUScheBR1g8b7K04K19VM1nxbnH7QRpQs2EQNxh+k2wMuU/hY6832
TWwbVDursMGOWT4paCWeNeiXIx94iUG9jq53PssSXuN2ueQWpWEZE6R9vudFAHCiIaGev73is5DC
/vYpAKgwOLl/cjlrJFTCrRVSs8rD/kDZpOdq3S+ROmHmRdGTV/cVJpoqNYPatvoYg6J4a9xbJEun
HcpwyNGv52kiFpG2ygyjof/6DiEyiAbFKQPNU8ejvOhB5RfUD/B9RBhr1dSFUGraj62DOSdX5jIX
Kvef+Mj9467oUNH8t/zZ21JBV/afAxu4Y0oF1AQ0N1IV0Swy4F2VJGNIFbhApE2byYZfYjQuHDG3
2bvSHWlGNfVs6Vb1YvXAbMpunkxNLf5B3yAMRgDqrXcB5oI0E+ojJtSVckqpLtWobEZQP6EFAVHu
5EBFgkjBmQ7EYk7Ir9+mV8Kup6asrG0DMgs1uRtLc4uBKWrwLmMJfX8O5Y1XM9FkuUFM7cV6QONR
L8cbqecWZUl/14d6VOAFV+PmRuN7yzq/1WTxEwcJsQSU5e6DZwoD8dvLtWRuWXqJnAJOMf5Qh944
5aEW+wWgquCrhBhmcji/uj0TgcZzJT38Oj9gPgN39M4xXk7rRAXi5BghwIigtq8Vdo+DU+mszJw6
PsZsklVHgQqbOpEfkHoeLKto//V1La+NsF7pFgEVfUtAfPxWH7I7U3HMvgrwFhmrwkEgzsEsZ3t2
wLPalpty51T9wW24OO9FEdOAsfLl0KA6Ki1oy+6LOwiVAOW2txDGaNFb7iCWYYY5v2FHG7jJu6mn
l4v2Six3UUP1vOLOXCGaYkL8+FbuES6YupEk60w0135mHkVgDCCrr08GxmqiJcmLluOWUVPipxXr
lq9hCF/3WzfxszAu/vadHk2eb0OBeS+y4QMP6d6ohc50YL1KnhOPHoZF8OTWZ9I8ahp1X/+hdDaE
NxemDPZqXDJF9iHDH54VorO8whLMlMYd5bSPtOhTD4luqiRK0caoU5KwSZFzXN6e3FXUhlgCK5hH
7+/3TspyQ93phLS9RffYpal0Cry4wNYP5y9v8mBUgJPC5ib1YXTFTQHT9HYVX2KY/NxDl19QJFtR
mhQgszsaCNc7O7w05Xqz4fuJFZOOw5jbvW++b9gXaI+E4IEHFSvEutPTrBULYB1llHogzHHvH2rh
bAqZKMID7Uin9smM0ENZAUMJQoxgRM8LmziYxIix6qG0rzXUh3QeLg3UuRK82EEFHGOe1UNbUqO5
hpprOS8mpWgTRgc5/ZtvaplqnswH+Kr5BolsHjGOuvs9O6osMI9423BrBQYAPDewM0Laf5XSwK60
Me9R+UFgzs+LP4hSuFiNOlGcchAOe3IY7kL0N/rmFCrcWwv1OvU+CrHPH8EFhme99hC+xGqrXO0+
2lcARbF2wk2d13oM/mKNHRND28iSRDY8VWmwsNubr9aFwY+qnL0xFttjOvpEH3TSxXN1bULUwDKU
geMWi7hGBiXcEkSLV1K/pwx9mdpaPMR3Gpi3FquhnLlMmJj+KlDntx7icmJscR6h/mV2kXwpLrIy
dTLSPZOgeiL/Pf0CS4IcXR41+D8mB1p9UJK5iH9q0qqs8QxAXuxAUJhkxxpzpADVqpBjpAftJYPB
dZkNcrLeyVnQZbTIX9UBBvk3mYFc5evvEhWMRTOpfD5q/9YwE7DMZ5AQ8ldJCWMuhvKpEcNFntLY
ZHfipEMr+AkjGSyMoyeMOkSFtgxbI9hjU/elS/2GZeodAI+nzNmC9F3tB4d1/PMKOiTj+lvgsER8
YAPBP1NXNEYnaim7NKPCTlaQdMPpdKr9PqUIrxYJBGpubZO997SoG0WiULzGXzIEQhDighnzsorS
F5fnWXWpZ/VIbx34L40v9KznCh55UrzzTGIL/z9ebm+2ygkRleAO28FiU9vJPHbv1RFB0ypBBL5Y
IuFAQyf5AbQGHjLCaSJP2xf/0fJOxheI9pfDwUKyYGX03lsxHA0dWfAREVQMx56gv1YqPWlWPdPI
z992j936vlyvtxToUt9bfdKY1/j8VGRJ80sZ9u6mlpXd/DSK5Ok4qgUqeu6YoYqQfutKVB/OAy+X
Gdj9bDPuIlgw3v+dOtdxJ5BsVa9s4Ra62K5RPJ7z3N1TNsAzgP5XP6yfhgs47CsRDUphafcx9bgX
nUG9IhteSfWBnl1LYPirvpK3BqDEpkCzVhdFeV3nVCxlrYlgZUNfoNNVYOW7dwS7SH8AzDgkCz0j
uxihsWCGNDPfke4JM4leV/jpJBFSITjmRJASj4RMJjfVZ+H/oXoR06teyNe5cyB+wNkbXYK6mSee
8k1OWywKoZRlehLUH4blQYNM65CzY8PH4noLSSUG7Z/AycU57WFMzFNQBBBw0T47URUzY5YArBkJ
b69QeEZ1PogBMWZAxbur1agQPAn4Eqig7rBc/w2kgUQyaaCMYHngyX11ulcQ0SckiNHMaV5OZj45
twGlMNuY9c5pEz6BNsa0tG/mWrLwABc2DDPgvEol/Ko+czgDQ8+K8R4tyXwzf6CUxL0hBnMtS7pL
FB/plNn59OiK8HjJgsjaBpyT3c72lz34xArKjFjYtHNToCj9KywD5yj/JijxdcCu7BGS9sYpwmJQ
0eR/oQ7NPJFn5ci5yRy2yDbmz3hlXZsAeVJhJVX8k9Cy6la1i6OXrg740/T3QUdK0Km3Axbk/gLY
zWlxWT8XjV8rD7mLBbGJ3sTzw0fAflNwkXlp0Mpe00238TZRQ57SmPK5zmjXyyAeWrn6a3jbIEij
d1yUX9renFxmWcxCL7Xa8bidkKLvReMXPNwTqjirjUft6q2ZjT1Z8MoGBt8V3C0r484SX6Jmswk3
aNE/XfmUut5QoRVyM2qGu0bAsQkAQzMV/UduBXVqLvEIbBjMEOw9RLfu89xqD86/qegN8sdIGQgj
LXAQ8Rw5g/SXSSLj2rbIeQnEuAHa8dhpeEOk1TcC5oIr2yAxKy13nsui+jdYDQzM1YFGte6a/2uW
rzaSRZ2Q8YCLbvoCQfHmyhImKoxhwH6YyNupWQgVBag7YbODd+dQPXpr3h8hpc+kf6VFYkwYSYNH
2cFOthN0IDDJqJfcdskp3909BhLneHKACGv8acTfk/8oobp8xbx76ekvz9lp3cr+T1DNMHEgHl4g
HhYqlGoFXJUQv6vtCR4WEc+JdRYQjda8T3SxxwZU7wC/5xwkNl+hUGUsLe9WyYBWUSPLQ4gHjxN8
S+U1Q9IvxVvyek7yPlelD1svzlxy6Cxa1399WWRsV1HiyyNfCXkXbSzsPlrNtip0psDZcLysqnTx
bpB5Un7+ov3Ywv5SRdeb1UjNkWLrsmfrVsZwx+VVjBSWVlM8YgImaslYVXqRPVNgjXwB8ktxaaR9
w955+tgu92dm4ztLUDCZBGp15u71NJWkfdIyYfgPEd83Ixy61bQ+UxqNra3SJER5PMZdUh9emcUJ
JkRefV6OpQFCyk/QoT/5WqF6NkgkDvqQonAlNtzFIr/X6AE9UTiH7KalAwfD2EAg21uwH77Wxn+G
3sDHX/kLIo54UdGRaCdXk/tBFpo6KrQkuacNNvHqwT9yNR9PSRnLHC6m6XOK3a/THrXcLnCC5vkx
gjftkgeeTpEI16kuueiX2lJkaj5Ek6Bmdxop8IUCWb4YxR9GE0yBA9uib5hLiZtrPP2HhMUzQKeX
1rmowqoz47TgYhD2IzZAjFYoBGXkPQRO9/hC0BpRZEwIIftsDNQMYQQFC5KyRXSkmXx3V3dlQLeM
GWqg5jwaILQezpdt5aurrSxz80LN2WVJv85Ggd4qGu2tH0NPG6KQ3JOOOgmZvmzp5dBnLyJ+6zja
jVecPGHMFBoylLILmAzEAWNp8n+T/NXZkDwOa7q/9XN4Dp4x/c2aUth2Cu2twTSryhzXHm1up+vG
F8uBYBtBl0NfRajfBZigFk225R0rL/dWq7TMNb96haDk3BcmokniU5LXDDRCQhbG2GfkqugLvmmG
5fivO/lQ9j+zSpUo6xssM/ailX8bF+xjVRn5IljwAyJ/fytSPuu49LDS/t7VctM2gdw/0jku18WS
BTlNAMqRD12iRr3QQb2d9KoZXwhrzxoWEx+X2rwEIH6mBa5zU53MYjF0qEriQdrsIeEKFff/wNvT
qVQLPkQ7/nfk4LYO4vdHpTwMc5vXkmxENMuoHJuxvbv/IgQ7fBp5X9ije3jJcryf3JPkTA+uY0Vz
abECfGQqotnRhAL0SHehtmZT3x1Bhm0wKXzUzYzDjoPw5/fSt9esDfKWt993qyMCbM6ohOyS3KqR
DjS7n9DLH/AIIT6AyIDgSqfCp/bsge6CVIVPtZPXduXWuK3YmBujHr7RQiKWIesApRIE0OJq0EQA
ZDpIMucfF0B0QCNbS5HwGRbrp77NAREZtD1jOvsX0nJqjAWNXRXcC3sE1ZDYCEDK9xEU9hPbwBIt
ycUXSEN7GTUBiWT693al/iRUvZasWbE//LkfECOY9dVk5Ksfsd5TT/wF0/y4gsN3+23XXgncQmvp
nFXJTuC4bwYXph5VcQJlgQIaQ9k/cqFDdkiCBOv0BGPBOQnVNEeABkUZcHRukD0L7Evfh9aTLTb9
syi96lnQU2WqA1bQS/9PZMETxMHxmThi5zz735A/K3jnhIG1X7R7O3sBRjCKHXXyQ9/mEbYqyhc8
Oqwc6QzuuEzraM+4lkGR/zFyACrpOaBNygksD21iPm4icESOtWwn0G9PrAcKHCpK1GVZiKyP5dTi
gyjiweadLCTmxYBA9XDgI05EFiyoRggnPAciVy9JDO/kHMAYPalX36TWiLf8pmW1UxKnd9h1HoEk
pHo84LjTWIjjAc1v26eQLkIuE81M83cJESJy2P22JT+hzog9IB/J1f1unLm7ImJR3qXWWw9IcvXH
++YVM27EWNisVdcHQgsrmadn2wTEd57AXAj68kYcoXLfMaiaBakZu4pmQV3FItsN1p7pHcTNQx2j
Wbbe88rZS47h1fCVuagcfa6YRNIKS1ys+HUcT5J+3v4vxTiYZoTWPPxClMJ9x0IFsngYi+SwjQd9
3nR8w8jFjKzRJXD6biE14br958TUdvmRBolsFnMcsNbENRIAbGEipfRiPnIl2S3tjq8T5p/zTo6V
yWgNqM7SyMs78c2LlXgZp3oCVrpF4HdHNamZ4BPAMsgdWNzsLaDegNP77xZTN9+fuJWxVNnx/qj3
WIkYLwW42d/0kKs1XLwd/mnySDeeSRWujMETDJWV2FOuCqIEvLqa1htFFyNUhsIfBrLQuGyiRPi0
qu9LYh2KZePnWPZx6YnDfp3l/z6R/x1hTGa64QxpBht17tSKltVlTKY4SDE0VuQu6D4RTA052Qlq
fy5AGUzvfjhcuhvvYHM+pUMCDPld8BYieuBtz9XbDlQU+Tqd2hCcrhe7FsIJFy06mnh1qh+oxX17
SouguTL/0DSXVb4Hd2cKvP49uLnp10U3gt4pgok8jmGzj64l4Kawe6zYmSaKxaSk6VNhuS6OfPuD
3vQHYddrDty2x+FpetfZNOItUyRBgpIS599d0kDZX2EG7PtN0hFa0jyuZApmDWRSUnHDdvm9eWab
PnzFxZ1DvqCp0F0i64iEDVOP7qoSCOCd52X5IcwEMgtWQphQtrIUs+v7ofF58XAqSILuu9ndfYMs
4zUj7W6carB9hA3FBrHpkbF6wHCg1qQOKI8RShPAoCGnUKNIY+Q1aNoDKLwGvaN0wrphxyP4aK59
2nqA5bfa6CXyiTiv8pgLA7UrydCLY7EeSuLYFv2d8htMtIlZ3zk8lwMOCvATqmIesqyNGH+aOi+W
95wsCEN5IczQZTfWRSNINnQBL9xrRcOnPyWdhNDEMSSddpm/n40h67BVA5kaAcJg4hjeOpqQwwti
dMHPXBoLUIq8Fo3LPwk1mIGTqK7ZEPl9UVRaj10eqO1vHordSqB4rtTpDc2wPRhW+1Ks2EstpZwm
KXQmI8VW10PSSbcIY6YkSu1wVX55dn2xkhNWFY0HOUQn3MoGuykczzYNVZNDd3gYFWrfR67/rr+1
Innj+H69Ibl4WUt4y4hNSZCHY10yC6TbW4ZGtW3L4KMVNC4Q7FWX87OA3rvxpMjcY61bMPpvk6Wt
CbRgJdUsOmrKOE5pSSh/jJJiBN3jijPKTE9BRI0+xtd5Oo8VX93P8BKgjchTtk9Ukn5ahooowO0p
oaZpYAb87Dz5J7Kmv/eW9dv7FbIZkcDfwuGsOjuBto3zUNuDQ/+Oa6pFLmAr0BSiGppfFhKDSSjo
LDSpOXXccIQm5prRVPiv5g/cTjCKU9kKG8ns5zQgGYLy0XoG6Y2tLkuU24NgIyD2xbu8u5ThxRNS
OCpJE8p5H3nf9WDcqE4m/z+gVzRAi85YLEP8ReXODp76itiGBtlh+8B71lgTO3g1VZqUoLM7CPQV
EHvjxfplPRzwsN8OF9sNV1fNFl+l5/eP8QzgydWU/xDVZXjALjz2/f1+MRdXvUqqZ3Niqtsw84xI
guyHrUZCch8MJ0LvtYyH9tSUA3Gz1exabx2TpFUKTJ1U0995zYX7A6uXyYsfzZHryGiINwhjEcvq
wIQAXt8kPosJ8oeDnj/+rNEknQoIv8nf7ta1JwFw1ALWmm04myrbDidVv31iNCC4kJA2pA+/ZsPQ
S6DJsRUkydsFBTtuKJrw59I9nxLPUSXK6r7ozdEohoSDr0SwEP8AbFFEZyyHU7ypA3wW/T/FssJX
Q+QgHICobyjFFtZzwQ3nbTBZkhYAqvkYRYHD0w9PJdvcb4Z6Iqr1CVNUrsd9i052T0T91HBFkFhV
hjJlw1/Esi62qwczW2lAG8ggIJIuzFSbjn0feUBCMFVEpaQLJnYXWj4UtQdTwCLhcJRJ5f89EKFo
vM3SgJzNJULBDCr+fvOTjZ1Oen/Iow9APkj2komXtZL+9yMtasfciImX6Ci+REMgr0kK+KiVlESx
oOv3mo3D1iTh6I8UcCwYtnrKYdLAXR1Az9Zqn35AX24GqwhzlNRzX8YjJj/6VGIyRXTVqj9jnfGq
MnsX68seAzyMdrTj9sc45laZnUi1dwIydFGtHLs5R6D1j/5Bs+ZPGrza9vZhwVxn/l/5I2r4dIhE
n3iktUyY1EyJpNYlhckpg24nTn66RXeNgcFRfbwakxRK6h7ASAlJdaRvuPGx5PXid5U+gqb4yuAN
2ySLHvzs7gvAGsCGrfbHU0VsDcxEZJ5LUiTyyO/R8MNWQvnfBTBl+3jFUBzFtnkboRZerM2f57Z8
lsLkdFKAVBijDWsBNw702UFm99jE/ibwAX731H5oUB/rO6QDCQsHwWGkpbsmZ791RZtFJ97xPa/R
Q1nQUHGfx+MX9AowJLdiHcCKjyRjvBMY28xbIXZDtRjZt7aYhDfBjQ8gL2/6KuBaDgVifKndcb8C
zuLB3nX7tjBy0QLxE5f/M2SE1q5bhR6g2QsY582Q6n1YvpVlVnwoxpPftdqkbLH6FCrQ6+VxaIa+
JJQUtWM8vW6Q5OchZhqpy4nHLhR0i+bkp581TCQj2WFlV+pjuv/NA2eO7ViCEBuxez12zmYaJljt
PjXVxU5U8+DrLn7egbJkxGv490xgXACQ9y2BiC+FthxxM+KUTk3rHqZjg7CU4xXx2hgSTUz6ky+2
B9f8qgL99/DNG12tnvrhiUlfK1qy7PJVm0ZkndQxaB4nXJbHwWq9dUoPAr+u4FvdFaDYGwspgv8O
6viJJykgVIpuSSZcPb96zw+s5/wbLxmyGw461EZek7QVZ4J/1SifrNQCId+JO7lSagZxJGhu1WoG
QtkQpNDcDYPV8UjeF22u3xNs7T2CwCW3YUtCQ7iDEA3C2VGLCIOFY2AXfdaqD4wflE6FqYD+SatM
RmsxueuLaQFBdDueFZ+tiGb1ysK+vNjYOcLCR1X7NuHJ/9uEgWYRN8MsBgRrc9WNjSKhsgV045fD
7HF8RAGme2MS/HwBvZpeI9BIPLa7M2C7EqfxsYMMZZpvbBUP5DSJChoxnhVH8eVXHULCPjxTJRln
+QIlQ3tDbax5iHl5OanI2+fGeGBdKQsefKSxkxmB1DQGRCK5SaBMup69LHEUVs6nMDkSJ65nKBzQ
puH/GjLS6AaeJqujFaFjRV5dQnFTQOpSgaTtvccbAixiZKZY5YXDeDCHBwgyY4wPdMxh5HCOfl/x
PQdCPY8IYTMOfcCWHAvxNMUkwgEK7i3zlZ3NqyHnOzxOrfk0rx79gxpSSKblIwZ1H/XWYI3mJOvM
13REKta7F9Q9b3GBTemmP+2Mg9XB1YLHX6pJDJOvtxbS7Qm0xvMz8yjC2kMM/OmUx+RdAJ8/PtF6
x0yzCTUNtnS6ody5R0UNjNbQW734n8wBYpSckIBUQZCSdXHr7pyip+Wv1r8Kpy8TRtwOD28TlUVf
YkM664KjlLyr3Sus1heIVBmTvP2eMfUAYBkj9vUHve8XGCrgp1H2DUiv8aROHKaPD0Wf33/Wq0R5
IadXPSG6MGdplfJCO4uGTbtT2NOsF7Zu4ry62c1loLGUitFss2GmgHDb7vo9VINSXowRMt5ZDMMF
T0d62NvffT+AYQf8p6r7YNsL29/jI3eCe8ixdHPZKvi0Mgld51hxGjCICmrv2ZrCg5DnuJHmCmpq
GSmgbiLke0IX2FkE16vcrGHhMxhCItZ+7/dTnwi/PIYhp0RoC7G+5gAJhHqyEiFTrKO4TF6iDDTA
NBRr1fDCya0VBL+lp1Cmx/mDWvo19xTNZ4EXld7fUiBOUDYfcVTGhVMPK3SXj7vk8820axu9aE8M
6gEGPB6qLP1uoG7gW/86iBOWkUGGLLRxLhZd760EAfBYi7YUi7Sc1yp88JcycCbCV4Bw6E5qEhHY
5ydn6veTQcd9L22Ya6HmeptNg5bw/If3/LVIrZ9Wi9H8ku2QfQj9rwykjHL+yZ9LDWvZY/XlsBfN
yIM2vrgJPME9q0D2V0XhgmJIHjEt0O2H8I/rfhDKu/OltNEKlmQH8kwYcJ2AlEAh7/8+a2zCPYCJ
TinhkSWxrPQvU4+a3BkjLaO4KaX0SFt5RuHvG/ENl6OalyPGVYRIzmDpB27FWmIRrIOq5198gQEY
AOj6FvKvi8LT817sxu/BleJ4Fh19sjddq8WmSCe7+SE5XfmNJeUiXZcwEnJjzHLw6GSN3MzsxO+T
r4i/RqIMBYity2IRzJ6tdSuYDpbyCssD7t0yD2Kb96D8YBlDMfsf4bZPhYyyT5NoM8/r6uJ5MUFi
GQQnukyGCvb8mc3nabW4kIP7RIg0xnfFA2Uj/k9lk8qVRGZ/oaZJi/NFOBqM6x5aTpa50nI9U1Jy
Fo0OUCO/RSnTVXvL9NANlKG7jUdbn2au+Qd7x0nCfBxaY5DIJ/hjQNx4Xbh1AklLn+Ffob0CokQB
tTrKNgc8/fJNm6vGQm3r/twolJSd6Z2F8yuLCmNbYzHUOF5Cs2aZeol5/UzwffzgwgULpwzscfHF
LWdT0DcMNmCWPehzGd2ZG0Oobls7N5SJsbHQliPtMrdK+f35H+poIU+7J5/xxWQJsf4gDiLuCUrj
HmLBHRL6e+PVfcv2EpYXrFX3SrKBXH8eWeoGAzSbOxpKRmP7uHB5DQQDNvo5MJAig5rZEt9Tdiph
L/ZQxifMuGplY1QhSffhjaVd2MD09DYo8mQaZQa++8YFZaBakvxxQcBYfJqk8NrVXKg2oJtYaQ/V
3lWFqS/Yb+8jhwiVXcDloyZyiEvACh9OQ6txfwjqaov7f8kcoCrrxM58khorqL+9i9XkKAJPM7y8
hR9lK7/XHcsh0nb4/QliBbA5DqNdcDj5/7hXqFRX2FDg77rd1m5FtN7DcX97MdztG0CH7/3hfHqm
EcGcnOfNlKWCgYRFSDTKrp0r2o9QJ7JfLAG1TWeS6OZsCg5C0g+w0sWy640mH4vec/vI1XVVvuWw
UnYGd0KXtbdR06gxHfRyrcF8LK6rm5fhtqmJ/WyQfr8+4pBMSOMQnc8T0d24h6TNiTMIlZmqpqFU
IbrWls3aE/PGRat2ywEkm9wSBa79pgYFHU7hFaREjDk+ybYvO02yoGCy4L8h8b9raimckh32I3L2
bCt6Jwh9O+5r0WvzxY5Rpugd3cS9ZrLMXjphWt+KMv1oVjb7lJ6Fa3PhAivuSCrC2Hk6QxDBwq1+
edCZEPMYmTtQ0Ae0/Z4QSkY+diX/xT8pP8oPKdPM3xXLSzTJM8vDswqAnKVqz/7zIfM9PwsjMetl
KRlJqKD66NEeSKZQKsBFK6CI5FmK+sVF9NPXULzNbb2LDXx4SBGubPJ9pRcv/r8veepQQ0RYrzlG
eMV3w8QCzUx6lDSyTfe3hxWAMFXVKsgSVaPsfQK/787DJo5mcKE4wXVXi1B9QP/8ezyCtkNTOFkf
zhov7qUV4XqIwMj2fmCFMyN4e1LBNqLx81+6qzrCzifMD9tkdU7CENXFhguWwgEV77csy+l18pJN
xwRWvQFLP1WFGFNKNUmRwceZBq9ME7930+sWQu/BE808NBUASem9iHEuDKSet4wipU2ENOpg5fak
jmrS442Y5h5U5h+lZ+CgkJrbfBeS+X30p9U+IJgdjpHGuAtHZo4VN26xH7ZnKOLbSVX7T+Q+Iifs
omTI+r/M5qTnIByWjxzmPOLWnx8MrdKNaAGDuJ2bIRx9+h968qreJmeBdGdb5LVu74wEUNutXJ72
/nLCznQW4vPz56ykadLpb5PWMJD3j5vsyAEW4FpGwL/fNHdQTCQrL9P1TEAO3JpsEs0Tvlmz0FrI
UFp9Ae39m39KW8XDrw/lN4cQj5pVHzrdoPlkU4RPskFZfDiNmVHjcH24b+1GxxPHYCwsXdBDvqUu
SDsFy0qCY5qUu3M/3bD7pWJv/6DlC1BOM/h+MXU6mavg2BILlrWwsXE00E0Zhk68xOTdVfLTBol+
gr41GOdrLIEY946GiO4FxLemQInIiOmhT6mSZPVsxkoBkXDr9ablprvWJKEOwOEg4x+mUVLNqUgK
MsLn3xz0dkHTxOuJKKHdI+mSZc1tsRxWBPkN9xyS44xwrMbUib9WFg4PSMxOereSVWVs2a4Q+tFu
deosTzKew8fSh365EP4eur8PeeK5IXJQEoAWmk1SJiMWSAOo3C2kpAnJIP29laYl5EIchaoVq0/7
cnd+nYnKjTeLbjF2xuXUquU1wUxwT3nG7MsZZr1NC6s79jRASmc6elQJetc2FN792IVypt84z4Vp
Dzc8GDnED4ZY7uRma86Ax5/uvfz+jZ1Jcy0PQ4832hg6ZxtqEcBgRtGpszeKTMj8AJXFyCznbHhU
4lq7SVs12SUGhpp+Yio6yswf+AnuGw/DknRZ7AdvrMaDvoVwAy/Q5XSlS8VbcRzJqgd6DFX/kXN+
4NpFFsVO/mjOoDgf7O3+7AtFegFHXUTYahfa0hybDNqgGwR8xj10LQyW0FaEC4gU/FVGojNS+VVI
QLIpZCiod1QvOWPqccdF4sa3zsEI9IHQ+XJ9X++NlssMsRyg5eCF+BwglsAYNKGXUSAtZQtAaj3J
Cscv7XNTzyjSK5sQ1qXI01xgxkUUpFjWgh6h/H8rWo7yu54wzERXXvfWbgA/idgKQhtwSUrm01sl
T/+EAGDLsBOareiZL8BblZNf2Vro+W3/EgTmOPEwCTuc1kZWJK7BfDZTmwnx5w9KN5q29bV8eT6V
wKdj9UCQ3QdCYb9kn6z5xplA327DomhxMghPghjsGRXY9afsHq/hoQSinqH7ybMYUTurTxqvfrgH
k3O0oC2dS2racAqMu2lAHhbV8VYNqxPeEunjUKM+pzloEURSEqvSnNgRdmIb6usrKLSisj6w9dLA
tmHo+t8Zl0sJHj+sITk2pzw6xwxhc5kVdmvpKVLt3gX7EPMk6sOG2xUODY3gBzhEGV9xN4atKUGQ
TsHG/T9m7M+zg8CNm+HA0ZSR6MQpPKUrKJHklltnnnrLUR6HvIpEw6tEAKh1Az/1PXNi+iNOIoua
A0gfoq/Y74cJRWA0viqNuacAD9j9Tb6FK76IWox5Wgr9EpCfOl0KHGhsvFTv2LfQWnB2fcla3w1G
J1jY8xBgSzCewwbI9H6nZP1Njshtql377q8lD8IGEDXvGs9H+V4V9KdhOEvvtP9NBwUDVqzjleJ1
MFLCa9n+SSzjYRZv5LVvI3QnZ2MeyLcc1TF5S0kicJDGOWjsMo/tknlsksyFFALTZmXnZyViM6nj
/Gye3NykkEe+oW5w8NnvpvuasjC8DC5kjpdi/FFbCY60LqIhqx8p0oPfLTH5UpxuMvaei+7XSuvw
Vh7p+7Pkx3haULbVjf3sng/dr0ut+RT6lovy3TXylBDcu6eS9Kna+GLVrefXa1cj2dzyzh8Tyr0s
IXn6AmnmiQBg13ObwxwZzcZIkNwi6VNGx9oTU/8FSqRzzXdZ1FWl4/Bklg9k94DhjSFWyK4252wb
aw23bBz05QRhYS7W3xkfK5pPODS73B5NZVgZI9Am2BKDSs+q+TTRqiKX3naK+9xtUYL+YDP6KpoA
24x8gLUCvNc5xsrZNc28ENX/vbc4/NcXb5ru8Alo9gjBWPzXOrEEOQ+/bF62+Cz0L16hLM2AGTZg
qOVn010VPBQqKO0OBV0XX7+M/xk6t9i7XqVEzMfa/vIncznyFdMQF+hY3DN82XDGpPTYSvNau/Gi
2hicdadj7LuuRTvd8HeBTIOi+NG4pEZO7lE2tViVwbOQXdOW01USl+IL7muo4Tye2+9h14jRxt6N
LkmRNQW9KsqF0DWkKOwvOnN0jFqSeGll+/fGUGZKiRo2HZt0xGtkfAe0fLq7tyokCZQ9AfH3CdJ1
WXSFny9y8eNGnMCS2U2joQZya/UqhjRGK7f+EisQHsF2o5LUOU7HxWOCize2AjuZphLJV6vO7ieH
+yqixOqjmmJtwXZPAhMjqNKHtMnDeSGUiMtaarmHVfVvTJwFKi53L//KoeAYxAvn7nvdDiwxArFr
g0QwoaaNPuMxeaPuL/DnMO3cdWI4QGMLUSIAo2gWbbqauRRYbYAVWOvBErWcN/7oBe9S6xfQkrf+
0tevqBQoWPneq8hbo+pF4bdHw6qHnqk91ZfCjjw6jqNJSOb2akEcDlJ1wvTnoRJzkmjh4nenJFu5
MyZtRr8qyT5s3yeC6POg1+vIowHj7VVEEXoYJgEzowupd9ulS3OCHPS7wEQbq0g9RKg6Fd0Ghphu
G9x6ko+qKi2sQBDAsxpUvmClFGAL4e5tomVNHdM55go6f2B9c6qmK5mvXPXamlWCY3S0jQUhrCwQ
P9ZqO34H/AAm9iCBhUH73BdmgE+hSboQe2QbqxMO+7tbUIMAIayVGWD/U9DqqTpLHv8lscAiPE3q
aaiiD0IaKgqmXe4yfLLcdR5ZyTGa/ZoazOrfFBNFdIp0P2RSImSIPyHqSLuEcZW62ZXpvXe3D0R5
BbVgHbYL3GkRMtj9RMNPvU5n+bIOFwv9H859un6huW7JH094AUM6hnnOpNrVrekTJnwkF2cNh3yS
RelrEqA1e0UdlrSzQ4fkzlgamaR6zonI3qfjizmJsSnl2BijPjaYXDNNI1nUE2cmoFeuYE9IBVJO
O4u7aQzlfYzXsBqhTbh4Vu9eYi3xsoOxeiv9eVapLtfSAiNBWIvd5CN1avKyJuJ2873/KxahASw0
65O0/PpWMV9GtoSdPz4J9jxs0dsNALwYuEZ2V+lElHSp3AeX87iwoX0nEPxISLwfKWWva17B7VNl
3nnC9WUqKGlYKs2I96OGdziNB+HLxEa3B+i6HTLMKQZJw8syGlbm3XjZfAB33aPGYuVhQby/BU91
q5jrpqiH2ALcT1vXes/oaumI5l/SHUFr4MnyQ+kBCRnx+268agiOHuJ81E/EALeIwxCL5qKHiimf
aU6jweIbEm6cdNzyWah6kYNFUUnqxtfTLgRl3l81/ESM2kyIiMeowu4tNDSzbQGs68/ZXrC1h2VH
FtXT4LxYSJuXDRvmsK3VU8o7Y4N2H7n654TeZNZJ7iaLj3cYF17C/YEwN7eGVm+ny7oqRYnbxuzY
0zZ918AUt4eBm+m6Bpsk+Pev9rrwPwkHc0RC8mvn/HRgwMez1IhTNXC5LukLxYgTEs+qquXwG10i
CjsGXa4Pfose5CQMJe4Oem6rP9oGVT00YRzbHjJEEOP2uzUKUI3Krxl1YYJszPB9vG8F3vxBk3Wm
Ja9vlJIetZ33d+tro1m9yU8qNM59J6Tr0DJZKSVfa4v9Dyb8Hfl8oUPNbUnojokGtJUi52Lqu+mf
zz3JL9sYVf5ooe2IHnyGrMMWF4eV7Z4rFefkFPixIOwGIVRgSVtnNEfni9RTKBd7arOLm/1i7fOp
38UnR6x5rRKrBFxO8AI6kKzfWq3iQgbqMpfj+pO2irStDiQWeXDdSUwfhUi1uhDjigwRPqnsy7vN
Quc5ddJO4bLgMOZO4tLyK5FG/WcS/IWkHZ7rLdLvJYxvtldGguc2PVZEDhOTv3kG9JUq6X8i8vxa
q9Tvai6e7ZLVkgu2YjnXF5m4jiJzz6NPmobFkWiRjYPCZAPJQs97Io7geQQJdHw115EzReePa1bV
RCn7dVcFzhnIHdoR7bBhRoyWd0TFc1gX8yWPnOhpikNMQPYIi0ws6A3mGKrjqj9whl+UtZiMfwIy
x2mzgmLVFasOSWHHAsFqH3q9aVtMMVW2A1LEtlmDIUmE/C8VfcezRCX0d16HsXW+dl7CgRhx/lAM
oiVgdwIBzCbF64pvv72ZtfQuS58CAAw0gg8y8+j8ZY9NG8pMsgBYp0UNkIgKt4zFd+qyTXvCwHn5
phzLeJLp9uQXhSmE8tAI3SEtiP+S3canwmLEw6iyCQu0KSHlDw9kIxdBOwXImE3aldKJOtnN85zx
+IfNZV6q7m6AQuBnPDDLObw3RMHcs1d3VDOKfMAmBG0E70Ck4CLN07pDEsLYS0vn/5KrFr3KuPGb
EfDh3M9rfMJhlC0uKNsw8mMAlki11FItjNmK7WNBlVKNXHkJrYe/D+avGeTOjKXSF2+Jmulq+hbV
rgdYmns9kvAwPxUd7m9ed2HQ622lVNHDUrfpZI0lboS6THslalju3vGUJI7BlM0MgJhyHkhHBDMD
F1xBRJQJ2qQ7Rre9Xd2QgEGfZmL1xRSnpb1GX01U/6kFOKLDiUkPmyubLkYBA3MV/WWLqAKjskzJ
CFDIur7hssGTpA6ak7aRHw1wb/jXi812KObZhvW0uHizbs4SIUqXbq3Q7IlZaj6lSyhZHatqckpG
/R6P01RBzPzIaA1rpDsTrjtZH57dtxLnLOLJL1GeqgdBXrm54TcdxYkPG/9ySkmPRAPfw6c/oSbo
0I2zzQDRyaibyH/vW1lyO1yZIw8zjwzQ7+c3pHfpVWXZyr6jUdsjvNlgUIsO5zNDawINgquiP3L/
up2/ri+aGDKD3s59tgVpgQ7t/nsbFWRYWwtVvxxpQhtF0jZ2ErUHl1aYQTH3wQifz5y+5waG90Iv
a/fvN2jV2RQjm612xEKyZQazvCpaZMaHs9PeUWsksOar4j7Ztl8B2ijPHECBErNHQ2ivhYyScOqU
KWhg2JsS5IGMSWh8HUkeZ8tryZN2SvJ+S0RmQwFhMyvJGOO6rLu2wYylnQQhGzn0jZunbqQMQbf/
0O2OSS2/Cq2cgmLt5Czo7g9bkInmp01f3V956ORJ0l+VCs1EzSgKT3rmpPyV7t82Ea5ZTgyjbYR4
sufiOA9bkNr8LUs9HaDLC1pHBC0kMnDStOmZD8tJmfPK6kYXlSM4r/tLg3Sgwu3efyK8VFpT0/Jx
PhA44xKYwyGvCVE1vDnF81840zGUtIrHQ+MY/daCXahU8xwtaO9/JXg80HeDIYzauuslxq4GceEL
02grUoYsGt7r/3RPQ3qR5p1kjnroLuSXVfNxtTIqUMqBAKQK6Rl7vVk1/QI+6R5fMB/S17arBojf
P91Fmw65ULbkxxVnvrT8h3KLxNCOOrg1oOo4aBaoTtnzYLoJV4Ohx9S8/ZjK2DZyOZ84ES11mKEU
aCkvxwCe1KKvoUuclVwoUXMXMwOxmBAjEKH9aj2vMEtTbGHFIDnXWMQOT7yjNhbJ8vLjSWghb0GG
qKcKV1ZzQqKYvasnEgEDLcI+TUEGbQ/nv+SPyEGaZnPCnPxDFpQ4ZGk3pqxahmzQKt6wAO/BEzyW
bOZ/lFMubPKrsZM0QN9LDw6oIRBXjldXR+NVLiTVfxEXI+X93TuSHxW3vwzNT7uQpuoGdPuph+s7
ub4QV9vUePP5MeRh8427EKOs0M9NNiNqNVots7OK/aXH4m5+7fF7Pv/Lwb86zf4I0Tiq1j9TZKcL
jPlzcDrVCrnzs2IJdvGsJMudIRY2DFWWd0Cnj3QZwfWzXFMu8JdIGWnF1XEqiP71H+9Gk28hHhXB
j9mRlFTQZPfib0VYrZD1lNER7FR9rZ9ZKzuOPc9m6P9XFuuVBUDV7EfoO5K5GXMQVfCP9/OCYLQp
Y1KTxVEsn0dqqw+7MEmmlYy+hRDoKfurypX9b9UZEfW4le5SDmRglfpCNhhAgqE4UbhhuJZeuc6p
hFZmoZkSzFmKltu+Dwo0jEdvL2Rb35uH5aWHGes2dhKaQPlgMl87GeLqkGsafZjnkvThRHFxu8Sd
mocysUYvWPW7gdvb0EWDeU5lCbcq1DyzBvaUIMJmK0Ob/Ue2toFrMkXG2osej82QnR/i3ezQ0grb
9qu2iP/fULIbvwZtLQLqTRCX6pR10Ra6M0PdBf3xFwL/S+i3hbgDlG30M59ZL61dvRr3vigNijMo
SGd5Lgvq6TdCrlyVdOXqx2rYbjyAOY9qjs6ucxPVeZF9uaOfc7DE/rojD4k0sG3AYc87EpbxoXR3
tRoIbiEhiyWDpwihfmr16/LoyPn+TWySj2aUUE69xiOrVzuJWzIoXYGSqf707MgD6Ifzh7oRwzap
D3M5Fa6MkZ4Qa3kU0EG7wtSOYt5MdwjRwylx1IFeja/knvEHs24EV6H7J80ZdsqA13wCSFGcjRIG
PU8dSpaTPB1EI0hirkRVKVGKstiqUQlO8JDXJD+hCH1mAW3J86fgSmknbmUSbnhV3KEOxSKTdeun
mmw9bB7UdiEwpzrtKHB2igEpwv2y2RsB3Li6OniFVRgVvPNjp4q6WQfpf0+RIMXyB9iPwGxF7XOk
RUDS2pmCMFXYM5DbCQAcMmcG4SpxFldG5mvHq9bnky3vVGiP0dYhbacCl7OZr4P9o9JgGP1mkmsj
mCmRf367k7B2fpss/utgfvzkacC2Qtaek0nGXCcfvCK8ZpC0k543dsE2Mnx2qNaQ8bRuQvwwBNsn
Ur9Ewx1OI/AzhXt6vXH0v86iMSvCOS0MPfz59mraWzvZ02r2BhnN/Td1lC6XWiC2f1/Ag01/4dsf
2T+LZtwPHMfWzXtP9O7sNFM5RpZLe0t8h0kEead6N8CoD+JKAjN3UWAJJqsjsDTKrLv8KZgDIlhm
t/F1naRpLmsWIF4DZthGFBlwoNWgxX/Q5J1nn0IiN2BFI6K1NSW9GzOMlN2K36GyuyDOYcsERmlm
ybYYbYjNGkGnvrFgOiJk1vpYrK+IOWjCm8u82JIs/AIgkfQqOYwbBZzBloAmHI3SCTrdL0hJgEV+
5XCxz0jc1Fs5ccuqUxKSKFlwOQ5M5sfOcpdFxBFg7vOo1tsNTynWGz+OQel7MOW7q6zdDfmmbbtx
cxpBMFgBXyyl+/knFY8/AAIX3ZVNLqtDphL9V1xGgpnolYhbvITnwHFbyNj1hjBniUz3qpKl9ZHL
AVa/etxG5inWBs/oCbrsndNkNRWg0UWJJ7noxkO+VahDqQ/2cueLU3jaQirBAQWEVgRKE3C0vg6m
Zhhuke8/N3Mus3ww7U2ac+a0oDr6JfKM2B/EgEclGfNJmnINdO2Cj1pU5ohxb1oO89glAbH6XSGa
COzVx5UxzMLi2jsIYlRPqbV1cOlibRWwAsySdlyONVz4q+dNuxGDR+/JaHxzz75vj1WDPDrlGsK+
Qjg8ny/YapzvIHierHg8iOQ+VVqAiR35n4A8PdRhaLOt00FSwLMOjv1UMV0+LJmJPqz+6m6wgb+E
S5e/16pDL1Mx0fLgJCidfs2Usi0mxYvWi4P1E+WqgMOQbPU1fsZAk/NbvltrqPOn501b0abi50Ce
8b87J+i/vtSY6+bGTxCZWZXrzsl6eeImoTYTCrw97IoCrxkiN92Fb6fGvEsGVFWHnLkUH1jd7hy7
zssOS7r3KdRniXSsaIzjgDglJG+cS57O4wzfbjjTNKY7rmfKmsMYY+58CXIFDQfrEMscFR2u6c4J
AjRe4WVHXW06665i8kjZYkCCpOwnmn87W/CNE/TKJPVP+xm5SnmWik88YcOCJ27zHd83/gMRYceX
YA5gx2cRPewGoSUyUnlheUFzbN6aJa6N7MfGWF5C7xJTX8448bMmanhl9Jkq4vJiU+blqvEhLY2D
T9s9Sjz4hEfcJIZworf3arzU9v8jVE4h177hY72gSkRGYTectii423LnVOVF6F6c+ShW/qMj/7VT
hfIxtsSWT26ZH4k1XN2+bso3hAOHAw4awc8lX/3AYK5AfCi0jrLJEj2plcsasLSvv5EUPAdQFc55
QVmt38LMnpj4Oe5Pr+JRdG4HuBEMMWxnJ7dIYz9cXKfHPLwFhfJs7v308dnRNmdFiOqJdrQ/uShr
iKiQzv8wVlIpbPB8FUTXjTxbPu1RaJxsEu/8G8VEI9f6+VSiaF8dt19KUS76eQw7QrEQIHHGN4q8
y50N+PCdsAK4sStSUSMFKE4DwHLQ6PTc/GilQ2CSbFd8+YcC6fnTGTdJEpOaJGMOu0PCf77IUDjY
fFK3PDs7RCTYkrqNKYDBUujs4StxFwZTiKeom+EfCuKy+rnqtqYhVSTvVgwLTT1hoeccNEjy+XoR
rcMGHfIlh6pKNp4fJ8me3QGsq9q5dIHvjvChYhlcEt4Z7uefG53tXO+DpoFaY0dsc7UEVMhrnu69
D8pIa7Loo9H50XjoDVUrF7cZ07k6v8IN8P8H+CbV2s60o3epmOWkEvmniE/PO2y4Qt6GeeLDmfs3
5AiItTL4504WfQawI3mRCEn2tWNhD/wwTGHafnW3OPPlIFLmov3Lm8CXMnShYpmO/lWG2TOpuaf7
gm/w3uk2pCGnuywCQ5ZLw9wCSc4nZ8fHXirMXLnH9lkE5X85ZdtlqgssKWl3Rkk8NrOJfh5VpP8h
ibH6QzUramaT5pSJe3W7wkOgMCw+bi1p7cMHzALJA4Fi34mXqmJQcI+QmIWfI7GVDR57PiH3IPzB
IFxa1RoRUF6fLgkTQ8J18D/IA84E6pucGK/iKkkat0N86CNS7AtYM1b1M0y229auRZ80DUzhskgJ
euCApHuTWYraxyaTusjJDSRQPXzgaSdwvO5F8B4qei3P/WYeWAj3wePaLaj0eKp7VMWoeJDPCHqC
nXXv87gz47YCtTvC849m5j0CBq7pLmo4quQkGm5bgLttJhS+7H1h90bLR0G7BZ6tfZcYnQEHXLNY
FYPvGJ4gWjl+FEWJ54b0Hi3P81sG+hMEcKYnp4U0MdQetzBoQO5OQVkvJ1r/qPiK5XdjDae752PW
oQ1YjaA4eB/LgcMFNvaXWHAGPAazR9pwOMplzwbz/arZffZFwhc2plG19rUTrbNNMlRougCtSoyf
KtevR3DLMn0LBGCvsuIEPVvjs2rTE5Jw9Y5HBRVoDcR5fRZCOHV85AJGDI+Jf7byS7L/7BheDhOi
zQjoiOiRAHmR8JLMR7yKGIb+d5mZwtcqmFoPyv7cOBTKq/n2KQH6MZALwM6WgnJTFdHmnWDRnkhg
Dz1AH//Qj2z4k1s5usDG3Yk2ReEs03T12BYSc3YzpxfWI43kbcrFbB2TNTEUSEWo7F3+liLtD5Xf
I/CMeDweczb/XUY7nHc/JfUHHteGWTjikr1+AaRdPnlw+uIoUreoSf7DUSLKmrznuQbtRWkPpL2L
zeP4HuCCIpHd0KbanZexsbpKZxQyU0pwP/4XavtBjQc0QJ9zh2dkDTEbJphleqoD3O6WmvrscO1A
voWuZIguZURM783O0dZZTnzvwlMiZlQZtRTOotCBpBlgjlM5uVCGuYpYTwyfM7QLn/wnojYztan1
SwYmviuKr7GXZLpfupL3Uf9sgoh3c8zai+2l6nu1mvSnrDhibIa+hu3c9ENVLepWPxUyJ77tfK51
f6kCOY92MWh7lEUrDurIuHD8UfA6kWml9X2lVIgJsYcYlbev6EhZB94bYBLZ9VERzSGlzb+QKB0k
1P4Y3tU0H7PgAkQX9m8XIj/0Qal8/Jn+QbPPXWNWUvRjIujV+e44PWNHHCLWQImGHCctx/qI6P+K
l3MMci5LrPJp7B5Fp3tiBdRkA8OJWV/ITcyP+A0VEAUeBbp0M5QT7dOs0XJG4PyjF49emoR75OTJ
EelrbCRbeFWYr8w2AllnbD2f+l/8JvJfJdz58ps0nHOEL1UiFeorqLD/XBTgffGzmO9EVcDMsw0+
sYPFYXlpan1ThCfOSfvnQCtF/NRNuqvs0Sa7Jhko9RnCDWCJORdv/hpUqLYqQCenmJ9KZSYOO1R7
w70gz2A1rbPHgwllrFiPLt0+ZaWkZ5NptmCnVcixRNcxJFAw+V4gKP9I7sIrD7WE4zUU1PEHb90R
9ARp0Az6slqSn727rs8VKjCSlYFO3/AkAUUvc8e04920TACzcXw+weJHhB8lUegAeFqcBRJXhDB/
sG6B0LtGTtImJdvvBpb9dCLrFq5bkmpXvZhdKjUqXxUCinHIDr6KPINCgFHQyWbxnRejIEGqvl5c
2Wgkzv694i0dNjYlCskHlQmUzo/np6XnUqXUFIBpjGTMJr1Zy/g8IXsJPtRNPr0cJSKak9ypPos7
8nFu4zSlk1EBftn39uTgGBbgo1Zo462CEPa2QSWc6Nsr9a8PYYJkVilv4geitL7OoeZ2LNY20sWu
1Nh+KTHQHmx1IDkQ7hqa6yMKfCqTYaUSkQrNIGSyrl6rduN3+BM5a2m3E9FtCHFEab7CPzd0Mtmk
By2+a+QGFvZhFyZTQ/kuz5UsfzOhZGbLKZ0oLPSvSJROck3utJ0KnfE0WwXwFExE0PXPwGhhoApo
42V/a07F9MiwXMzws0P04Ruz+4pzVLvXUzR4tEXZDPUsb2t9x5ctml7Y8gx1rW8EuMVNdJxnwpST
ONOBDe7iegKwanIFv08teS3B4yxaIGDF6RBA8HUn+tRUtrRCeaz/PsViQfiu96nZdi9oVHjLeTcH
40+T+et5EX9mQ+wb2W/IbXzmyj2+JidrNw7NG5tzCSrAdlfI2BWlqLn8bJmqPMRKJp0EzbXtDA3d
tRurIyoKJap4+LyqaNZToR9kfq6n3KN7Hf5euC55ooO0OsrVSNygbY4WCM3Ym8m0cJJNjVH8588v
Sd5dpSDv7jcvSffEDt7RFGTYzoLp3x0vICbLVKiXUz/nCPc330m/ivSCQrfRbMbgpclZD1IYRjhL
rlVFquRx/ISjChQxXeX18Za27TMdA4enR87pu1P2AvkKDb/69L6z3ChHF9zT68leYwFbCIdOse37
1IjcL7WPhixP1+zv6+ZBJTDk7dYSn4757xUtZLRyaLh+Ygr2GoKAm9wBMRF3Po31bkdMuY47G5BD
l39mb4AeQiuKYITaXUaM4X6RkhAg2v1PPsj6YpM7p+gzX3SH+WE1Sd4LNH8gtZ78iROJ8LC81fdt
rp/g2VeO0p8QNsUWrzNzMavhBq6UnYc84KKJ82IQe1SlGeSSgvjuC7R1BgSQ2OzHkb792LZ03HDb
EEvZ/wzgOC8KkD3sEUECyAGjMHZJh321w9eARKgt/eIZ+Wbqkq45QC6m4c4Y3K/4bKWzNbJqDenz
nCkQaZBwBzMRaMpCJiqsbynu/2WCe/9T+Wi9VySK59g8A89mZMf+j9xWQOJB3gmbsRystNmFkaAb
co+bVXLABVG8RrLdvGF5N1+MChvTB4N9ovhPEqO9uMpbm4Q0IXHUfXFlHPDXOdDUDI69PrPCB8uZ
FBuofoZcLL/H7mq+I7lDPS2QptAAN3HLXIU/o4kyMnbvDDTOeOCbxalY8Nm3yqgfhfLnklvr/hlH
0tJ8UK82fzJf9JoRyRra9XcY3DrWYSk6Ppezdd6iI7aDVexCrMgHHFe8KFh1bFD6TAB+SWVOZUP3
EF2n7oLxm9mwOg00WhWbWtW4uUOk3cSaKYXbSV+1orc8ghy5bcT+gpTdCZjVG8QmjytgFxa+LamX
MTKUygH2Ru1s1g8We5uNzx4u2S8Vmzj+00ui4We+Z1P5DgsRYG8PY8QXRUoV7shWI4lVWuzpHDnb
N8sdXEYQz2RRTixN7Ao7xkl9aJFsOc0RivpkyXMTOJucQE8mVzXZjT9IfixsvSHOlJltKiBNmVw9
gn2CUXLHJzkJes43sh1WaNNelLyciWasfdYcktw7TsNvdAlJDozlP0bj4z2vEifqm7XFKURLEfjm
Ho2TRN5JoenSRGPvsIHeqTK0mRYrnUwACt93qd1DOFWvjFb0+Vt39xxhFDeuv1O/yGrxzFRt8D2V
C2uRcxu5uzhNx4QLhea0fLXcyaR8yplF/gYqpOJa7W37UeUccBWEWUEo5KZVBJyXjkzbtCbk1lBW
oQ8WNQ0FXxx4nDILSpV8wpN8qi7hz1OZlVKOB8PmJ00vdhg3mLzg2SGbV5b1ezT5wv6ImeqjjXyZ
9ZeC9NsRGdGvKhfwnCGZDQPdbw7j73pAdMLph5PPoEga4jw9tGvytp1UQKWTIimPPRegv1zp+B39
Yq546o3N20E41YCT76vEhVosdHQdyJpnsYMrfuXp1N6tkOY1xm+TTXvHLnLl21C7MdbvqkMRYB+I
2rgsUiHxmlBCTNc/JjpJNTur5CRTOsV/OU70IcUGeuKsqLRzcHJlyvaRtJE2F5AUlBXbE/lH0BiU
rcHrG25WLG4mOmnun7hYllVHreIpTRvewJgt4wXE0Sv82wtoDIgemWoZifJLFPfLsV/afLuqniwS
u1i5C++SNWM07jWVFHkbnA1sSkuNCES7yePdTioznPuIxIPxdwz/DCSKgubKaO4xyg5AFMjNbDpN
JkAypzcLsSnPm1cw+8FBHOsPXiSv4ZNar2/LA9Fh0fSuMQKPTEdfTV/meWc3p9RSyoxNtaOAE0wo
xQaywf01pAl1XyyHRwVypOHJUeJHZ5aL0MNVjManMctikON0NVEbc7bAmVZK0jQki1lIIPPqnJ6z
Z+BrBhyTwkZnZlcg5m/lxuHEIcmnqxunxfE8uaiYV33dsJPszFJI31HYbV4PoqoGdOcwdO80tXn3
PcPLjkFYJfOe4MrGOROfCHX4Im/Yzges1qzc37py/FMw2m/KYC3KOtybYSfZ/mgdSvGtVjx2v/Ks
XGAa9Y/j9mFxEqJe1+T67IF9l4mEHd81UVtb/FLXVTxi0fPqXMWPu7VG+a/BruV6SlXVjOTNf0oK
cXlSFqGbl8jbiks2EIGjyGg7U60QGaCUbkjdDc70UjUCsGkaSz+Pp/z/PsBwFxNNMRJSnZSZqO3i
EZus+YsCuFEoHOdlBPyKPjHRwcC5V3keAQhLtsBMyj0bjHKniaduqPP8u12TYfg7x9P3w998urPf
XQBjGLolhqRGicJPAjYBBym0KJf2Qg+DI2pRHFogowwZpJ2YNFumCukWvrUJ2JvjvCAAb8kQlkOn
sqXl9KfHYvO/ec/2QoisxsTzO49UpzX1a9qrsoWYjoUshwVDySQvLDYS6SvTHlGoT95J6trDnWkf
3JtgJfBRbz1QP1J3V3+OpeyrStPdrW+zdQuVzEcTskKJrPoJBh/+I/25Mf0Tpsw3duB6CGMG5xsr
eqKxBa/p6Ke5kfqadF9zZx5s5rj8NaTORGljn8kwx53fe7ysVwgXY+ObLtLwUC6oiksd24rso+mK
gyGBkmMW3cILukMnRbx6Axztq2m5vc3j7ybCvufEzThTjNxx8JzlGY4aAkWbI18CyxVZ8KlPEckf
E33coYjwLp1TTdSNA7f34Lp1OyltEzIcGAYN2aLRkytiUo4Mjm0SWYZsGBDgRULlJihQ8TuGg5XG
GtAQAeozRT90u+iUnR5zGlDNxbFvcZBFJnVvNNHhf/gxc925jttg/4+KpHwBN4juFn+cdKN1epAj
8Ouk2eVY3e3oPAK31rXstrN0SGEVfUySyW2VpOB8+Iq1BMP8T+xVWH8KOcvwmnzAG0AWMLCFUmcz
DtbKzMFNBRP82RkwqRNTjk7JY9PguXVHhAIN5hOFM1NBVRh6Pz6/XpSYVYYAzArqRFPaYpAKJ7s1
xfkTvGNF7yMdSD2VUNL5YT6F7lEV6a+Z1zyXyJBKmc00yQAkt3dHcW3p9T18HDyj8m84By61kwmt
LWB7qWG6e0jlE+yeO1p4HkdYwo7r9JhaQ+3tIOccJeVAQS7RYJGYlZ4SXIEodbkcSmsRrb5lMf4n
njtL8ucPkfyUfvX+GECBt8o+eREnWVzee6BBrTcMawQMpSI7o2V+ML8GfmcZ8nECI3/B5QdV4Tx7
JvLS514xo4oHjEPzIlUOmGgWzPFM/Wd1hqZHQ07a+O1os+Oco7z/XoabjR0p5Ku+ihkMDMHZoPW6
5KlSq3Ip51GOzwKcBwfrNxQBosb/JXWZBZeeuGpJVBMBmw/EFDmMsYPF7+9Tj8Sy3ncDdCXmdz54
BxnVe7smQt+P5a6GyWzB/DSiNJdO1CQtGBjPIPv/hlDcnSIB1fhpGlXix61fGxfvw/amIbhBbMkb
1U/6BwVoODbAuhVQ/D6yX59ftAkf8suXzaR1PNP/SJlfumwhYxS7JQy4ey4oxfAoAq256a12muVR
Hn9dPFEsam6b4debsbGOvjIbiYXPdCiuv15jIdaz7GJJ1Lr84bqvBCK5OaQGUbqDGZr30MTG495Q
iVh9eiGFuMxrrz1ABJ0cMxR6LEyxG56KNjL7jAml7G1eCNH5P4LdaK5/2N+ZAWkduHW2XJbYrs9e
kz64rgDMxcXU/ksEb+Cc75dlhBacOv3Xx9n1sOIPnkRt3fGHT3o39b8vOyW0K5LFkMsYrdIJXdhv
ttHdN7itwIZpQeEiC1S+IbFkNrQUP26EANOHGy0bEPl1Ft2xfk2IajNr8fUAUSppBc8fVBJm3s46
EaMGRSvaw4dl8iipfCJYAuetuJM0tSwHuFPCtBdpWMS8M587sW6ScmI3KUaR3su/lP9ZBekWWy+c
Y9Po5BpG9GxHe684x9o5ItjBdMO9YI50HYPXnHeueArlqVIrh6jTYKLD07yPGzMMbDi6TFLYBuQe
U+/Ec6BD7V/p35dzrhpo9hj+070OdY9VbIm71NFoVL3cfHre7DHm17atQAp2haeHGeWCAH6liZEl
23eWuHyy1yk5vnFNSTtsHYZ172vPjlyuii6jBBGmsY4KCWf+2H45zkNzya+M/qho+Q401upzUNUl
mmefrYe97t/9F+kvZ38OzZE4XOKn9pysmBH+1tNMCxSmVQerdYgNYdQ3zsiiOVyjYAIExtXNZozL
tKCuStAlyg3OIPFiIrTBntCmdsfzEmnVXMiApNBnLsJeNUfX444wfUx7Oybeh1aHNmIM/nhQ9DEv
cxI/NjgD3AQdpxt5UsfDNNLMPMdlqFR9G4uJJ+rPymkUc0/QG4P3DAhTJqYAtFCJSqSv+2UfD+MG
auJJEOg2/+TLhuZCtErHrvDGUhR0lFqFQmJWswvhrLR1jyZW5uo1Y2hXVO6eM0Hkf9SQ9OU8q9pj
gOKH4yldfIVgIJyY1fbNhQm0UNCGcwW3PkwrMtpxy9FzvZYeKUXUBrOOOED3xyRrWMr9uwPWWcQS
R7NLUTjZUfsq6e5CcIeIcaxrf9iEuDdibH4fNMn5ZZ8FoQ9xLO5f03hvzQuACp6tGGg2n5PIiSBf
wp2qOarZWJzLDVIPBbXh+N6SJ6oe7NYvCs16nJ0FTH8CWbq8vyEDRSdEzZMJ48eLApM2oO+YeguV
5CwKC6ci+oSV+driA505uwHAuq0onyXIgFzwu84hjPZbumnsbStkPgJGEY9IRRFCehv4PtGNsBBN
NRhwgLlGUpwcIlFUIkxZLn8ESAELRJKngYopF6IeBdNn44dSlMPkikeRrIZo22qkbFh6Zf0keoKI
DlKWAe3zcOl1mQ8cqRNq/vSBX5U8y2AAWpJWxmKNGMSubMJJi4Ilp0wAAizmdioraS/O/1vfiCPi
s1zOKcUkyDkVF279dri8Rk1xLnrZ+ZHKG2oHQIOol6wkIFU9bIjEfFjIgUD0K0C8pXNRS2HNwmAU
fC7ZVvyG4nqYYhETueNE+HKP5yyW83/vd7qrkalNbpFJIJM8KmLG9h2Tahb9W+JiTuU5ug35G64W
0VpzOuGAl/NPAKhHTPxFnLWwU2gWFZGXEx1MMqIIllV0Eeg+RwTVWNtpZdYPjorBVjrfutI4gcwg
OpmPvIVWYIGkbdZRWJsP6KP8qdDOX+So7GafqApSnD4rjrV1jxVxmirrjtKwiriz38RteXbRLaQz
XEsaoblxKu6CdfxYstI3eEK3JkzLTCgKIYQrUnEkdOtllu1UKkVJ43xmBRvvSOzN/y73erQFfHpq
DniaC+jwb+j4jRVNOEONnzC9ATgcgVNNHas3EbRcJbuoADDa3dt9u2JefDHU2TY/SH6N95HPauNS
B6Uq0wYJsFS657SQ9HpB5mxBw5M/t/LAtMZ6yKF6/TPb+IEQJWvVKwg9ryv+E4dZa7QWAWmI3qbz
WwxHpsPAmFt5fMlQ7qhh2LdV9CvxFsHj9x4l2Ulfai/5Nc51SiTECOKv3oHe3xJB4YQwW290lqSZ
i7/0mtjQBYIqq1q47lMxrFYv45Dfu6u3I/HN5WJ252VUm40KqHcXt7vWe77yZBljILVgyAU1trIB
JKYYd8YvR8SjhMAUcXT7PKHHbs+b/jZfmIFFoRilaENXQ6Ftg2GISNEA8w0wrjpf20qDAGLOfyBh
mvJb2qi0JjTjfWNk9MiEh4Q3qFw+7Z4UQWLrkJ/ugY6mh0vXDhrT3Sfa1U1QUdmL+Cxa1CNyFnmo
On1ZpdyJ1rocTVdRDJ8GCvBxhGwpW6LXWjj34QMpusyM/ZIUtEL8yQXreL34rz+RTcsi5PsXFxfw
ChR5K1lvqeHkk/GJGvy6FbnnkqPKH+/ovPRRqq9FjKmAD2mHC7MVoYbuVcGDZf3D4qNVGUR5fD2S
yWFdZwD9biKiGY2Vkv9qw5/WXaUgq2h9OIhAAjOi6JMgIExnPdXQUOLSIrLllEL8OAuZGM0NW9Xy
PM1hC+PlLV/nXEskxMHraksTcdAiw1B+UVN39h47fo+S2zG5ASUy0AxIBCZRd7Q7hs+DZjsU+NXM
QPbOM/z+UZSIfIJIJHVWF+uqaMgTaA6a0Amn4H2ScMVUZvW2aJ8oHT0yU6Cv2NGwZTBIldOPYkjd
x7RDRKttFGTjoY4Soy7P+ooPQtIGFFRDzTItui5xPO7MSdcQUcq9VaR88KPMeLOUno7Ypoek32k2
ciEsOmQCgQWveuw/+zNAyc/RMVl+SqSoukF+7f9poKFi06MB0b24bwZPm4FuqpmZPwLosgtgpEx7
gMppDKn2MEKd+njXrS2ujXsvO4/G5P7DfHxnfcyLjh3Kb3SDfVZY6iBxW+NFs2k44IbX6D+6HR/F
XtOr/iSPRpierpfjB4/f5ddz5LVDdW3aUReLa+AZchZIq1thvQ0zMHGIXwWtycscLLEDHfQH6jgn
AUtKMVDj9rNVF5dcsxYCtQobfmcJdU+nO1WrH7VU/3j0OozsHXlLuayS+/v1fzeIQ2f70N+B9XKj
VLtI2q6gcWSyWh9oqkfZ7SBAHLQ9ngtndl33ddAWmRpnViMYKk4v/ydBBhDWugXoPrDYTMeBqMkp
ryRq8J9CQBJcoGPlCZYKBlzxagOa97gvFNCeSqm+yHk5MP3WYD4AmZ/t0dLwpqyEX9WQdSFGnjJR
whFgM/mm44cDXn/6Lvyl+fSXdXjEVbdobFjSya+OwO0j4C2YqwSV3bb/R+JYCdysmYTyvO/KEhSZ
lZnPqE+DFpkUzp6LKqhrZLQIiciA2cOPeuhWEdvIn5wCUfS/CsC+skOtam273Cy6RZ94kQBdc2Es
TEQiNkLeglFzLvfDI2objUU5GE2SNffcDKLKHV99xQQrxqgl4za3+RrnqmXSkKyTK5fM9eov4Ls7
MJapNrjUL2Qj8jeN+neIGA//yTHgeK6wH+yehf+eY4sU2ekeNnlIC+VPJRAQIuAKc8oxMlsciLKk
q2L7w83tmXow1NLYTNSnBhRTolTe6K98GORZOcKUhnKtloRQCQenCmWfKxijTHe9gh4plnGNCMXY
V045swqzMKT7OHgQ6/nlsea9HmPMUhBumn/wLhHng0no74JnxU+nEtRBLftaGNi7iwhuOQLFKqwi
WtZH4qmGr4fj0BKk/CqsKEYuE2r2N5LPvuOGEiqOmfvcnbYgc/U/RHGE5/hKhP1jRCk/CalyVny0
2Vlt+7dCBQzSnD9nsyF2AIY7JT40O1vPoHXGkbK8Of5LmR1Ilq4S14b3soaPJql/A8IiGssxDx+e
oCYI6Q+mKCXlRgqpbgtQuFZMnMi+lpHBwtbiqCIt3yoF/FymcBJhuORYG/Rxgz9MdrL//xn46u03
TYb5LVZiW5kB+OH+EFKXZKurrZD1Kynm5cRB2iTY9xKp8DH2E61BDjfjt6xYn8vmxvkl08yxErsM
T4KKmt7ZFC+lRdhs+FYOiNm57vTpq85T9pgwGBzqGhOvT7v7zeFz75qmE3B07W9fKaSxxAW6brJA
HVKwztohnOvYB7x3ghYj9exWDW1cMEuuYYSJY3OpUNzE4hhVyoDFdrvKQ+neRxeHp73X2gEpwxmj
FLLUmGG8+WT2lWJdMcmi+ILGB1+qo+PNNyBBl9hdLmy0lUsY2dmchYq74GR6r4HXuTM0m9c3eP0x
qDW9F2zCykAJA6/nNMDOiHavoFUIL7pB7tcATnTkU6CuafVyTKVOvXUmw6PZdHAzcohemgXZ6y5j
ijoYJqvSgCN4xYdZ1URB3K3uiZiyrTp/5FttCWlfduOAx1y7C30Sy0xFvAX+R9KZRQz56ntRKSoU
wKQaAPHUyPuEyW3oBVad7Us7BeJAbcLYwZnvfUMGZH/UI1amesKQNj9VdgHBLSR9NBDUxhoZbm6V
wH2+rztCxvD+fNJr4z9nCTTycy/CUPZSIknXGK8zpGP39hjWmvrkXnP4OjOLOSjkooibC7sOS+6p
vvBz7KgbqsK3UR3SRVVOIQLYBk/SIWBH6vSuE6RMC2zc/0O72B6rSP4UlmhWTNc0P198LQs2iHUY
uJnlvCdpuV32DO2D1s500/6CwEwFPb5nF74eguolnke2M641WH0U5Qh0CHaS4ZRwR113wG5sGQVC
EDLEMPK59fjHwRoeu4WM/4y0QP6zUhStmaPqC5Paud5ZF2KrJf8bJgcnre7JBrVarwQtQ574MLv2
CfNLFYCm86cNMhwXu9nToFwhlfbf98RTnr/HPOBEGDvFvj52qBLkEO6AtGkvmMzQrDGg4cVkUxgd
7U5YI/W8x6GOQGO0hhgt4e9pJ5/Ku1VUiAlPFsFoF7C9l19pHqnxQtJVzTNI+6usEzKQnIfVG7pF
lnfwjw4CcBgGqsrnf15d5WaMXmdAtKJALb9mxwAE3j8fyWMa2dmc5xsXRKJDBWdZUBqX33LBoHFL
ioQz+7ncV+ybpGY+zBSzU/KFphRMCYiWLfzF63VVfz2fOfDojRYTD7N++3FfY6Vi/yeCe/UXFWpA
8Ncdci3JsVySY3eAtxdST+/pWLDmQkXPyDTdsZL6Zr3ul0+zsKmhIfApnB3WT/TdNQRuyIjCyiMn
iIwv23QsWlKK5q4IjRY+kajlBcvf3cB9UJ+Etpczv7FwWo/ntwR9vGs9Gb++EKnEa0TBcetUN2Nx
8yCT0SgQIDkdVmS+MSrIL0qghYQV2wkP7GT3qr/roOvEaAPPe/coEsPKeCGkwf+uXhF9A7Tax/uu
H/eLrRXrp62ZXmycB0N6ZyZe1Dh+m2PXc2GpH2eejI3OJN0kPdBDywO27iBvFZIDmFmtEGH4pJ8O
/ucLp3ly0Iyc47e1HqfvU8bFp3X2oJ0bAHPUePAmhTFcvmHIytswk0pMwoU1F4hLXcsTMs6Uuj1w
P+cRzpWeZSxo5EHXOD7mcERnWhgovZvTRd8xPM1Q7gVxcxqbncybnySWMNerbG+QcPTg/MnwqdJi
A7/cRVncmkiBhqzm++RE0DSukRHOUV2sJnOcSBkz/mUDkNGQyzNnhDTXhEa1e0qTMMi2bztaSo74
ZG8Bvtz1tDe5Od8CMtXNHZT6w0FGkGWdVAWo79ZHvYzlJKwlSvpIajYKwhqhedyHTJHb406ZW0Al
SdkrY9G2NhLx86W8abs+UF6CCAEw9OzFpfHH1A0S3FkFouH+C+VaxYSImbYBEilaLemb5gU0tLMr
2Ve1jJHrkxUnZleagG/N4girfMJbqV7FOPFfdWYzjCNFhO007LrpYOi8mfn2F9zB+qncHuRc5wXE
FNs52IgNFCogUcjedjIUnuPoOqOlM3NgmEAt1ye0ec8J8yALW376UjB8u2ZLp8kDzs+76HosPcac
VZ/hk4jZZOf6i/SSSPObcfxVAP91eu0SwHWvRtMZNQFMir1bCp0/i2CL8VhwlKy2peYOeOFMcfDQ
6zQOPLSinovXBWFObKL0T+Hzqtk7195SgUk7o2MiropRPf4jZgphHBIFBWMFGAPTaa8aMugmFHze
Cy9K4JhE33Wi4BKaxlVutOBbnE9no4QjOitOlOnF1VNPBsk2KY648MaDWhstdMHvLlcKYizqohAk
qgTJUu1axjMyypshm+1i50Q6huFkQy43T4zlKiOE9s11/v86SU+OtOK9GjVLfXYnvkXND8GaB6LI
mI+3drjDntqGMWbGHEop0qeGb4P9yrWsdS+l4nxEaS+xiFln0JgYnQP8tByak+nQJ74mwLZpA6E5
KYmPQmRGoxlPElhVpcQKztzlZqzb1KQ6pZrrpVNcMSfTBLx6cjo+dQ91SxQYQ3egDkJ41b5IrjJU
sWgJ1PrA0rrv3Z+OiJmZ12IggUrPJ3o2KmFN8qySY0VOqf2RwrgQbLx+FpY4Ykeye5hgPCoH5W83
5Wr8h3MYPADTnzDHgnN/BjaYB6ZXSUyh35pApfLzxElzQFFNbTTZqYEwFYdVvvME2bB2xqYmHXLU
QH7VadxW1khQtruY/9kHiiq0FBzNbmxMeXyWLw01xzwbAb2Pavh73ZykHMfI6bJtOcufoaBwsN6j
RX9/tv3o1H6cbS1FlDgyHq1gmjxEc0KVQEBJSSBn75mI148tfi94xu97/n08gAkfLiUbA2+NASk4
nHI3LVA5UW72TK+FjNKBBTJopLQMIc1Qqqd7WS2ivF7qhl6T53XFFNLpNyh4ZPbJP2jqNlXeNtsM
yHHq65GMPMzVgrQFUZ643XfAoQ1xVDbzAH4lrVQvR3O2GlAkDLG+taz++dxShaAOb3sjDiSXG2hH
ymYg5atQnxOInJEsIamDkit47BK6D6q6+Ly0jd8y4ku4kkK72gj/2YatW5k9F6/1/cH98PfJ2mcc
SI6YX+yQqrOb9I1gxSioRhClK9oZNwBpCmYFNvCvqk9dPKXw4VQYx2fD6OZVKjYBaJm7Wfyn4+z4
jFf74IF1/TnIKqd23q5N6S+mxxROgqLqIhKpxf0Mf82qCfh8gRJ7Ynra5+MFfG15yqJTkECsXx7c
BT+4vQdHmjXEotBUNpBcUFR3rxKaCza71U8AbH7gdclTDqK13JxVETdp6R2ihmfrzeCPfPey87vq
aOUMu2Vf8Y4ojMGroeR6fIJFKkVWEBGrUoMWMWDYqv+z8jatQK+F0ziwZuDC1gtxr1RncNYkLKyh
SPqgH389fDLzmnsjh6GSoj4kxT71TfhGO/JM9CIt/WT6ZDaIp9SdhL477+zg4L4GNZkF2SOnejvu
IlbL19ttAKWokdNNKRKWNWUI2LljqSVAO2sTRvSmO816nbN1nwApHoJHrtxnvY+7Kn1xyGk+8NAd
KqtXdXBim12W36BdBwTIEndF5V95FvFx45YDnUkA/1fkvT/uEuTcfGXFqFRjRsz9u5b2E99yxmfz
+Bn8CzsEUNgvrSsl2bh3ZyhMA9n2ujNorzmQpJn5a5VEwC2W4RYf/cntZWCRxysODmBC1SHcfwb0
x7k/ICGVaareM9M7kApHPsoo0Y8Aua4fb3omDXhiYvu71Id1hlRpxxNfbdJg2wkVrb3qHdLXyd6v
dOxB7DoYJqZcZZWh34b9zaYRbw31vC7SNWcHYuJdgvOsHXZEWFIcvvvsNbaZ2X/t2Ax3A2IaqwRZ
lIichYwpnTrrRnEEQ6TqUY24IjNphYjF1FR5ZYU1VsAPxeigVK7KAXTsmYOHv7WUQmoWMGsTvb/q
ng8okS57TEOWl1SIjl866jV+EgOgekrRmE38GHPvuE22uDy20Cfg+Gt3MlVwoq03scjhIa48Rq3b
bBGtPQOsWgvJCgFtaK94e0TpKNe17mg+UeOidEdtafUdcBxNxmkkjqVEc6tek6SR77garpvvYcdy
zLtzS0mlNsXlVTDwNwvW7RU8Dz1hQ4QqmXPqxbMEg8vUp8F4d8JDTb7vBxFD1K9JFePCFB8WjV5G
JGVc9Z7INa5SYVoDCmmwNPha3O9CCUUDePjh7VeXkHk+za6S2r8f58p6nhImhj7qrnun2w1xBU8f
JSBiOLGM6wunlKtYLuzGOJWsQuL8YbEd3/BzFYFFia34Te6R3Yp4sVXG7llsbjeYkupZmdAdxFEy
5BeHFEnLW2XzemJYvhrHqrK0ZXSMz09WycDJ5jGKB1mRiY68q0wpAvGtIbmRccvsygz8JUaEwjVC
dI7bdhxOuJTpiFi+bV8So8oO6hOMjmZpw8D5kRhKWYyo6DafFlPJqkujqbUTvUo4T/bGMx1453HM
rfD8KyCNpGVQL3ik2Du5WGmsvZ4o3pbJJOW0PBYfqpsq7slzhslXn3US8zSFDl/99J/BfRN0pRAg
gUGyCN1APRc7sViYibsE4xL/XfF6clSCF10YeL5En/y38sxCu99ovQo2QtUBjHq7gJAFgQpMGBmP
Ut/E4KjSRl+UpFRS4tFZUQ/I7ICsDaaCRyK1Kblrhvj6shNvwhDCCgYmL1/qs+Be1XVLsbu8zNEG
SreMjplufy/+TLKArOBwqaVPLKNMrrjen3gUavHFtZtIPY1/4zS2rOKAmjydjSITZWGWiPwWRLVZ
vQcYWUTea+G/y+qSfqdgKh5f42soCqmgrF/8HmmId/RPaGu5cfehJ2buFxOTbUnf8szuP/0xtCxI
+9MbFYwC/qZXGQaWUdPnV7DN87klQKvmb/hoBCMOM0MgA0iKF/v+SGWtegb8tDou8rgzGjduuYIZ
5pNmCZiCQfi+YR1EWNuPiVT09ybVUCTHuj+4bNGBA6WrooSNpRdVfFVxxfYdMl+O6eOSxWGZN1xq
f8f5Zw7PgqxyhbJl3Ea5V/9GaZ6Rk7D6UChlx0CJk4Vbk+E6KIc+H4LBKSmfI/wbia2iCDV6f0zc
GkxOfSSnNYquy1BMN7AuygV+FetKOQMJ/m1cABv2cWmiQeFjkDINEH8qMqp9JZlloZNTj7lHCEiA
0xUhbAIe1Dlm98y/+GoRkh3kJ2Vk379u54WwDAYcxRDvU3xyn4oeVGfjPWQfQz2uywugi5H8+5Zc
EMnBeuODXD8z2WEDPHQrs1/phk3BTlD4MJ3LTojMJAetcrzQCDpS94YaXDQufu49Jdvk+SFPXjGT
Yz6+4+psoSZkf9fx5+zEgYK+Fn5Z8XIqBUUGpl+dKEt92YDoyh0EXFm6xPuTGKBqUE/jSSqw9RK6
IRsadMh1iyWJcyd466Usu3IkZqYA6bnIZg+2XktOSOIeof6Rocj+D0Q6sU1/g068HtVz7JdgHDOW
jeA/nJ7qq/zJYbRqtwmfGxxtkil8p2auakTwpJn75sId3WP6j0hQEuA+iPOe+e8pZ4Q61v7wWy+a
ZgafkMtff6ADkAHZIMQ1xpZwLOyYeRssRhFh5r5KexU5zGYer41ZTcL2I3iI2tMfIiT/1iK3PZpG
rfUxThl7loEvkxoKaftjoak30ihh6SarenYh9yFDJcNeGnuwpwwIwVgQRCxEUBdC6Dbg5KJSPM23
42vQ+w1AJ+Gv13qHJiRe3RFoUI3I6STGXgOFCrwMRwp/zdSrtp8s9gdr3rtQ0D+EayPFHeaggfBK
KUmmnVepRY1Q0HW8cLVojGBldViaDT3SC+cfG2L8kbYO4G2O1xD+pxY1AiZlO7Xtl3lfeLaYoxrc
LwjV+W4vunlvjlFaOtCMUjib28hsbSwjjJoHfGzHco6EplBBs95xrRgfqcEudZdDrul+BnBxPkoR
inzyhJ6GshwfUT6Ubp7r9t4A/2a83PezQ8Zcj4AG65V8jYgoWd9q4jglSSiwr8/wnZX/YbKlAM2+
BuAfo+iPW6O8cvKSYzZeromCrSUkufMgRaV6KvWNES1PwKGpZtzjBQUg3vFGcZBFdc6RvIlor4YJ
nR4HuFKxtrRD6yWVPOzHozVPAX+1xAVoF6I9qR6x5xl1OrYJvYqgm3WDrWyxO4vR85PozFL2gx2O
9ts5wIqyuY2KjOjzXL8246G9AQpppH+lrOVrHc7zta8bZs2Jor+Lo2OrU0nlKy0P8ozNgdftlejD
2DpALm92060dosjJcxirEzBflxKjSgdF2O+SMER8jDMFmQKA752a4UmFHOi8Yf7qR7rp22ghAJae
oZo218SsQnNZyBqe39g4YPLbAshpY5O5RUgJAL2UAIFkwdn7dVdUlR814N5f8HTVpoyp9/vyuloo
hO1okyZL2VUDeBcRrIS7+B4OrvX9QDVI2A/1Tor2d9H4f35k4KQADvQJtJ6kUXxFxQlChKmsAtGA
LJ10x1S+hTo/Oaeh5/m/u8ex8Z/D/bCSxkULDJplnTN5iSFcvGWfaTAC+/ItJI6CQhdyt5qglbat
0AqoHJyL0D8pfe39YePR9+C8q41oVIbmT13/RUo8amNtoDL5wmQn1+A3YZyqZDSCIV+9z41Is+SO
QrC55hTeONndpSQ6BHUV20jZTu6cM34aj59G+YsJ0SPKG1x+yjiU/1W02E5zQk9cLlEwd40+UBUY
hewSla6C9cTS8eBugYLy0OJsV+gQauZMIrqd3I4nvUU04PHNS9QRZFsmOBEE7CgBj4YzZNULhFp3
hHuD8m0x3AOHQYBcHsA01QTKJZAdeTxTJJjvtoT9WYhCr9hqXdvP8E/b2VgFwyyjxgY/1N4qXTEl
LB/XY18Md3leX3At1nbk/ykW+XwqGQUVOlrJ6RnM4zFOq7kS20hxLXouAdtIlvzQ63BiJ+c+Rk3I
WPUADZJYtuw1JidA6iu072x+pHQWQLkxbIt9vsho7iPyy0qJf9Dg2VK/wqAv+3XYn48R3wO3kqLo
bjRSPlgarE6PmG0DewIpL9lbL8dVes/aajlYXoMthjj0W0FD+qJy4TVzLpv87t+GXcq5XG4A+IH1
gTxQBpBD0YQSGcM750rTbjpfiRMvh/XR8XPAymx6UnDs9O2cjVoYDuUuNWcGi8+Ey97rNkWZC6kq
kvjWq+n3l61nNvFlqGBeruoibxxAfz4PNNu8rSvVYawBq1flNWsgycO+TGv98yVEfxC5QT5EX1xC
QVlAWU2X1KzzXmPrnQ/n4/6K1YAbfukxj69dFfJpwHuyy05wXaDQicd+IdUxeK3L8X9g1FTXYUEp
L1WU6LpUaIykERoHqusqK9ditF7h3n0G+jU7tMoZgO39cYEaVU+qpQERVswqxIbG9KZNKzCUg3IW
vBXcY2JYVGYDOs6dLXYg8SVxilP0IdWgLIjwX01bKiQWDQ8g6vBMc1WJOa0hNi+y+M1A54/MB373
yx/RB1CNqCeEaOVbLbzIqo+rKY4Yfht8j/pdGDDWAclKRDTyphHZhqfgNaJI+6NaRqG8k3C8hefJ
DT0qu3QUadng9eHQPFhTPOqTdU6ZBBY+8fCyTcv0cn44nWXrtIizF2ZV5mPAd7qJlBsU8PcxLMI3
432eJzzWZvZ3jt5CgPu1BDw17/XPzVrBs0X+t1EDNbNnj2lMaR+zHosOeGHjJ+MD4ORVVBmKVjge
9jvLuGhRnQeEE53eF3qyAHDZFtwz1dNRKls8PeFe4qBwAqNBBX8KlKC92rMNkRkWPzx1FnzQmxT7
Ic2IyukDFmmEuNY+eMsr6hrYbD9/2nXuZPT7tPW0txOceguCm/Vshy0ZmkGBPuu0JYTGl7wISena
13D1faWrxfxyg2KdRU9kYLiye8yDa02X7YA7a9oJOvPLSFE7LeaYMHuF7DiBiAGogxI1jvPyWZp7
pcQe8VGMO3/ZEC6fFN31/rCeeoF3mA0KWXrus6H45jcT/UZFwkXWFBLvbqX48UmjGNKmz5JGDrwP
FYPhgyYJLM7wUjBcBvPLmgbNYQaLqoSZiBt1IfInHtiydnnZtXCik1dTEu7FlXgPL3/5RMkpfPeD
y/OjBbwqW0s1D/AkGeSrKnbBgPF1gSHOWxaBiN9/94NxDEt9/iwQSKLmCgXCZbZjuIBaBOPz8Kmf
T6aR2EeMso6uoP0vG8KcEkaE/lFcS0JGOzD0L2RuzwTXlSv2iMj4gikuR4/rrp7m7r0AgjB6qrKw
Mk2SRldkl3s/3QoWVByOsBtiTNo454Ha5QAUgO6l46mC/1RSfDAhVJyzTEPcvJo0PxXag7FKqmbC
6cmnCmTm48Gl+lqKPcINhADoIlhz7G1pPfa4h38mDupJeVtkXo+O7R/oiyv2/yE4HRSp4Pd+9sfC
/VvoatOmLdDxLpRXPShqPYSIZd8KmS90m5th+OimgMbTib+1qPwZa50l41m49BNqPZqfs2qssYZT
amVGWneSUqKOSkXmPVwaNAkPBUyMm7phM3UW+soATwb0/aV9Qij1rR1faqf1Ay4eSGdYiQsoZBTI
kBKbw7OjVC1381PNnvCxuNvPZ3kRo9niaEDsfUI/YrutjfBy4U2kKyZBIz8Dng1EjoLLvi0BCkUW
LrFpiah8p89+zA6LK2pKO6rrgVsS2082S4QU9dJ3aOiqCnBCVSDC5Bjy7GJxdLpsQyY4oFv0H/eI
ov+ImxO6UxOkq4G4A5SS1VxU6xHS1rDbTE9jF18psbd8B6MgW1R7i9ieL7BA86JkyA2QUFQw8v6A
xbEPprP8gTDM994/y4ymnODvW21ftgfyfOlQ06kDjQ2et/rTMzLFQgNoSJgKiXXKezb6Vki0S+6Y
FHvrkXgL1j50EFexLexI3UKnljIjAhKdyadWAVIdRGH8gXAS7Y2vTSCuD/jen5X/7eg8h4rufOLU
vziXUi5Etfj9mnFkHNsDsVp0xiYHLV1VEe86v91R5SxPzHHESoA7KqamJETkre1akzjQ2JPmKFW1
x6ibfbQFyZdYNiS/3EVMsCPbiFR+mVuyqGiDz2v+YASdfFT9jrZKU4zLeOcYEq9KOIZlyw9Kc+7R
kc0N8R11diF/nwZuzDL1ZIC4xopOrIA5Y3hOLBLap/uqpcsYZySuNdzzCBQwFlikWbM6LHwoDnvE
nkatGPkLJmPZEtGjvEkX9EwoHI7XF3qaoYU9O2qD5frFsDzgukMUAXr8nhInlp1rdsKJ/EsScm+n
WiSwvNGBHsRrO7fuo7q0rTGtmFPuzBDgm0AiK2EO/sZHrdgYaIilF8nRKFU7A6ZsTVpJcGRc44on
oLNioeLjBsuo1zDQdv3ouWasjiJBHNli6/wtCgHUqdQDoXwVCNqWNxL3Tqa0VLvmAo/nNcMrjhzF
TnvJGvy3xXdTh36P57Nz633fhj+kI9Z4mmdwLmzlXu7l7/Q6Spp/j+HLiUn+eBEPTIg3fO/TuJtQ
8aF9zy7X5RvcyurTBBqhbZBqfDxQrU6QideSIMUKhs1Ru/NC030/55IrtLLhKduboAgJ+xofxXso
LN4HeJHokaBmUwmXzD7ieIG4EltmNSBnPMvxI41Hln8tgASR1tfxIVU7uUj4qeA8Ghrf7dJaHE3z
jbK7jDPWyLuGBzzrvwoLyYzpJauYAaJ3pZBnUhB+H1uGQ0hJmfaTvzWoEzXcsobTNgxrYiQlb3kN
72hEmhoHAo6Hzm1gknM3zYphQsfXh9+kARRq4Y0xhsg7P7QGUgl+awc2SElDngpgZE1ODybEtIKy
vRF4bS71n/DnMotQb/n7DV9X9hpJVAxWzXfsC+3mo0l1tBSz283ACRUGtnk3h/oymkVs4REJCdA+
XjSESIYDe20AG1GOacUI01r8mvLgxrN3lw+FJfWynGlRKvJwMCYTcjvF6AfpEkU5z5DEqFJGEYFf
p4GgkdhYs3tfnGrroe9vQOt/3lwjfeUf33MTZtAsJQn5ElXZPLnIJiyRO02oW8sS2mFnjpV4npau
VxKML7yd1qXlU92CiGn6s7J3d6H6qdjL4vX+w67ZmFBtuI/vqLCCVPRa9zQ7gRxlnueT3hn+ly+G
8V0lYj24fipVSXQZ0CtFEy/GvDy2NYaT0oDXB3Jr0hVHzLjewsZm/QDX9uyPqlAsmhJmVnxyQABX
hN7KEC3Hir5gvioHiB2k049kBBEUZgOnSErUw1HGWJxwHaHfRWW6cClQCsVEXqb6i+8Dm1KfH7ii
CRIUZpfm+qvUw/d1Pg0z2H20EjUKrXMcryuxqdAI098RHrn8OppC8HTho97rW63rmHhvrjnulP8v
4CLGfKqMuI67G7TzVBU2V7q9KYLVNTXoTKU2wVLbC2+0fWMIHrpi86Xus/rfEUFHk0WKoz4/boCp
xX+dFOQ4BC4fYIPuIM6TjlYMLp1iyZh01bze4v/zf9sdGl2pHP7TizaCRCUK8vizep8tU6rDn4GN
Vl18aVMU1oAZFhkd4Vj8TyIY80ViKjBiYStj7GFDyYub74NF+4buzwys3uOUbscFFExwAXxOPiqO
X0oSW+tVV0l+JiZZw/yJ5qezPeIcjoiTNO3i0xPzqwDkVfRi8DNL0LpJf90TMS8j06MU9Z71YuFc
SvTndFtrRyUr1zE1V6tyfkfhY+/WdcgoP8imDCneyVYDVXZFKdYnbMUQPyZ6yOozwdWH+8eZ7S2h
UItgX8mq2rfs+B8SYCJ3bmbwmSTPGpuGMsf3EA3kbyK9mM1jIEyACBxVIPbL4F1JFIbyz5SGafSd
AzonLZGxvLlkSiMDqLJu2N2inxiFWkEw1dnQjg7qw3eqw7XhdBe09v2y/s8stj1x97eBy2jNfVQv
SmFElaMvl0NpHQbAXxIMMmTnCYYfCg6aJVaNwNEijBIpVGHnPe7QSc/snYnx5JQR6JIdwOfjEkmV
B7R5zOxRV5RtTn47P12i0fadfy9Gus5sysIWMIFjwl89ZmqZaqUGNxLZ6ZqEZg2kR5MGAdzzko1P
O31LZ8b2gSqN6RLF/gJTbxXcNnM/2NUOvDMgGZZKwlXb5vMJUyZUfsGLDS4Ash0tYP6bu6l8SUGP
Z1SRydHF9h91P6lQ1cDAMaui93N3OE0je/OJiWMdlhLvMV6Fi60EvVvlQ0RwQHLdYdXU3Lns2wNW
0kjsLMuYIxFMqhJy4AAiCJ9ZsVhAVKAa3xovVm/ZTd8Ocs7TGG6SIC00th9ki89v1IEKcJvrws8+
7l0SqXl6Jq1F9kfp64wCgbnfF5M9VZZP21YE/TqVqtbsu8ko7j9YF5UB/s3i5Ayoos1fLrT8+UP+
mJqNY6zKgjDMxaEE5LGicc/7qei5zJ2uFHeDjR7ZRNxD9j494jU91jkvCeqq6UlVyjjvKutxPuuC
SyrChY+i2GiqJBRnwCN4X32Vv4ExG/XgekIhbmWXVw293kqj+FJIJCUpkppyVPwDrHC915gru2L+
7TkASOoYiAXR09Zso8kZeWRk97/XJM+r1I6rNiGt6O/hEXVYRgAWeNZHYD9g0fDQJPzrnH1KeOFP
a5D3D9myJxA9lIGQ9IEqP7kEkJ8GBQ+PbjqC4kn62pZy5CP0bGbGFghtILow2RoOaL2UW7FQ6QhR
s/VmQsMNW8fWkoqOQ0nHXYxNoA0HhBD6VTs8fad0NW/pxEc3z/S735rTH2Z0HZJ0EMo91Go9/W5t
pBbIH/VucdrxKBgbRRyYbO5pX0TfJbPRCD4NxlY/Y444pEdeTmbJ0tmACUgEcbO2VTmQXZySu6Vo
Amc8oGL1VCtdzLcD56SEn8x8onUP1JSLTBomL2Qty6yB2O+FqQFZvKFhsN+FnrflwRzDREqNpcN/
ElnHo0TsPvURBkzSB/y4bmlNnPpX3wd5W/e0LTIIZ+NV81MULvvFOXizdXEO1grSxaFSH90jzjYJ
NwvrZ76T5dHcmdtf1oOGxU77G912oLsRq3rpXGp+zdQXrRgRPi59I/U9W8O9/Af19JzYwKjT8IT8
rDKsGJ5Srkj/rIhNgsR2Na44Lr0muB/ZEA+XkJpduo4LqvW+cHgOeE4YkareUejedtzBtS870yBU
UVpYzBW71xSRoZIZIf37TxfgXvOHAtFe+qqqtNe77LZMng5komITUvds5Im0J+Fa5iKWiru/o5VR
cgd5kVkaMTHGbQ3EKhjz7AVUuzYR88XlrokYOOxLdiffJgON0udxO1/beOyyw/uBpqgTHREG52bH
3uuVi4PeBvv8B9h8z2FAppWMSEN7J6TYhMPWKqDz9x8iTZGad16dI+hEKVbGLN/DDz1LyJ2cKEkG
Zosu/IaCQy9ZVG7wsPNHz/X/RcJ8LOZ+/MquIsL9YzF6HWyfOrgDMkz5kZXr+EIDVCpnKSSTtVbb
qscwISmltkZDsQuRfbcjpntavJrxWksE5QyNEtWleLlo5v+UGD6huDV4HdMrnksccyr8S591gouh
VSWUr47BDy/H5C227XQ/vn4+8nZGQnED6ErAkFUEX6EbhvsII0L1Eh5i3/KNoV6u53nsqTMl+foV
rPWZAjdmhR1n9+NE7+tcuwjXxqTvk16vLOwm04zqICyWucasTZ5IJ04vjYaXCQC1MHowcK/8f5wU
AXi57s/6JrlmF3PvS1uH1DkXfmFsC8PIHlALC0BCc/Brsc21BberybF2nMy5sj9fwaRXQYU+Upq8
vnySLby64XLTQqhNaf/X43JWfPVyB8JqI5gqdibTMFLRN1MeIMfbhe5E41DigHGe26ovCJFxXwvo
qsL6xiaovBgy0KvzPjQ+cnTdOwFS/FnmYTGENE9eIiGQScZkltMcEt6jQ2kJEYJgLQ6KTnoAfoBw
dAFDr/WQ/11wryBHDbiwmV4g7mom96bwPEF21yzZgxok0WAtZSNFN5VJAgmI6OmLKVXPH0zccubO
l0MEKADIQgiKNTWdpjXHh20RtjH97tk1UztANwfKuwU/iAjUVlbanQT7qfAL8RClgOUF+G0PXIVn
NDp49y5WUDwMCLKaRZT/lPY41lUOTgdql9BimbOKgLuvN0+ZA3o1BpCJrSmOz56e8Mlghc2X7P9c
gll8G9ga8Ol5crPHctPYYWhyz46nGyiMUsT1uz9k0FEMRKZDGN4WgVdURONsf2SbdMkGbn47QQGw
I7WJK4ECENE8IgpTB376KAPyzZL7SYaDMDx83dMEYCaU1VacpgyXr3FhaDdXzQDng3Dgc7ud+OTh
XBB1/Et3BNjqbXzBQa1Hr8IaPLlTQ/oyKXj9tgvGeiSWwKhUJLpiWXUTeNEtQVcognewNVEpLNCr
5jj2D+FGo4EB0UqlHXq3mUKO+Jymc5BU3hWIyVcRYXOu36W6HmYr6pvoRDDFwzD7Ci37PCpERaGY
uxA59Rgo1RqV8RfWJ+i3xpsAnJMQFwOl8Pb/gZN1Dbv5m0T2XQwKvYPSP0A2oqYLYvjyrVtW4TwT
lXGgoZnQVcdug5lfwPch7BwR0N8kyOvSdUHldxo4Df3XzklNUp1CVG/Z6GJvg6g5sZZdZ0KZS+px
p/qT8Pz7khksxRi3YnI4V2urZ+EZT1sps1uc6zVECFkuDtNnhse/SfgiiqvdPgVWKntfaIcE8+yR
0y6K3HEFy9NnwAUVzCG643/4od7uKMcEbT2SkEkV3+2hfy5KFVaCwuj6m/JzBbgsDpv7tSTSjAvj
OajaTEUnWFGrAws/n7vh2Gjhjvs2fpSMxumXictOy0KBbNacif6CdG+ryTutzza8BMLMEa/yUZXI
NNl1x0RT2q/K/dATW/jvRwdXEY6tG50vopItZjFOPoON2dhw+oz0UvTSTh0FhP0D8o7l/d19onDc
A+sgxy0YvWhapFU8Bd961j82Guq1kNKfJlg/nlEshfeldhbV71F3ZgxgHV+61Pgp55AbmKEucpJZ
gZdjpeooH3Xal3d+LY2X8DZafikJHzn7rHfvjhaSRZfWQHIHSdWDFB4FZlDaII/INltOiEfkQgxh
hcM2c2WoDelCnTIaJyMySjhraNzJiXcRQD7pqCYIHKUKPvC10rkFxCGG7E4rl20Ka7ilMk2KDaWr
9692dtbGYlAyZGGhkJRufBSvqnIs7ttfBByWyB581qzAkYTtxRqKEqosjRfw5y0OrO95+odYJidT
i/9c/iVdbHcrp1UHXpYdSKskJp10S6iXqoJLYvL1at1aOu+5AMZXiiOldeXXyH5HS7fMwsbV5kb7
hMfkKSxer+g4hu3nN3TM5BN0aVNr6Aj4OScOPpIU4ZZQHHoUhJZHY3Nilv3B8UBl0w6urOC1iHov
+wbdnW6d9906tiAKt7Cayt+SYHPa3Na7caYGEgvsfcevtVqAH2DInGXg5Y3qYNRY+R0NqhEUzC4h
uCP80d5Ah6KuQdnFwNYeJDLisKvIGB+5DChm8yNB/XV/bCOnTqiC9kGQClTNnMhZmv+J0wOJwHFN
aXL5n7y4LPLYf2b4WCWuKVVjKGnxX+60Y/vqt5DR3KD4cPp3ue9sPeMQZT9IJLzTM83lDXNpIKh2
XQLdzbE8g09WPocpnaU26rWHo3ifRNhA5n0bhpw13LXHc6Hyyk0/L34Q5eSEfRsz6R2t1Jl8ONaS
grycV6VJb0T22r2Ah2Ee0vYYuBf1BUFvEAgeciDKEOV+0vovNwAk6ZNpH6duXN4/zjOwrKB0GZt1
MDrbUAuuRoIHvDa7qgaRnGIEWNiSHjZWCgrEkwZ98eOWD4VHZ8VqHz7F3zFyZ4G8pYCyrbqAAUKB
m7xq1uHTofyUkkdgAIDxd1wejnrSgjobBzxJ8WWQTXjXVbTZ3G1oauhiTzgqcWWUMYFCwUL6Prkn
mPhn1fW71YOeZOA56KEPXWWHNtP6g89wHcgj53y0zLBK/OCuYmioVOCUCOTwvwcWizkXPoOOmYAo
93kDunJFXgjLXVpP30Yvn8bP51/eLC8UnJugy7El9EwG8bjSO7Ot7mgGctH3Z9Xtsx3PwMBxDiHw
FX/pvYkuJq08/VOGzyTDYs6kWhoAQ8gzQsONQptOhCo4dbhuX8axn4d6MCBK2lolg4uMMmRs9RFA
YJ2KugFnB7qTSIpJ13pr4ihjOOjbdMLIm71fFqdOyGg6PdcuLRB7HRZgBRhY3A8BbXwCb0JAiLgd
dToRuB4sku9RfWlRJFG1rimWx0UcZsSVxXmEaUxmRf9/2P/UegA/tXMTNSJU74sLKqRtMIr3kx6n
gUgCimYI0A6fhFC3HSjYj1JpPSuQn2I5lZA+C1iQgOrWi0/O/UIRvnEyDf1JQmzFNa5X2y39mbQM
IvlCTjl1EAfZ8hGJ2ipAa3XqTUVfGe5EIic8qxDSme/g3jJdotYxe+kP1PT1tjt8+jq3YGbbabKz
WvexyPy46Dcx+AjWQvNKUfI/Noe17S1NuyaP02NTzpF+nwVOJUOD7r8caFohWe7z9aizr34lURT8
QaiUhWiK9H0FqI+wAMUWyKFO0PgB5KZwqs9KCEBXHa2x4Q3fyXBiwsCZVv8kELXsvWR3FMklx2K0
016tZoYMJ/hP+GWj8bLjg7EuQUZgeop7Vqa6nnz+pzdF6c8D58GEfwHu2o2JHvDDEtzA9EBwc+fS
hZ77KQBxOw/BRCQXBtsezYqc2GRVMUcv5H3Y0VBt27FN0h0dCT9Jq3xvxE5EiSdObzms81bOjJ+5
J9zFVrvypgLI4TNY/ynY3osv9GiBZhCftbPL1GKq2qU7an/iyW+73JOwoosJRdFBPPXGqSiMeYW6
BL5nRV6IVWMb8o/4WnbjYCEDbhLnGWX7dn+Ck+VVSKirFO21+fJoCNgd+32ILQ0aZS+amvgkjV4J
JHQSeKo0qvyvhizWTqXSbsOT6iZJlzfHo3tXcVN1cplXUjCiG+PaMRCWwdkYZb9N5vFut3FCU20Z
b0iIQ4i6qN6z/o/a5+0Qlbsoj8DoV5W+OGAIj5L5JbyNUrDEyUQYv0FjidTwG1PD6Tx4WISOZWc6
qoqI1nFklNEqNQ/UKtFYXPKGYfmfuar6Xb0TbL7QAn/9lh0sjX+U/l9lFXyLwX7Za3O8U2P2T3h3
zGJ53az9vvgMAiPpdcvxH+nM6JVJ9ZrNfaVXXVSbjuG1bB3y5RYf1107XXU+X48RBg27Ck2wuhOX
gtPk2mZOj+9vXcvvBUzLe8c1nagEqLBhedtN/DybCmMcKWTt6ArJeYgkZ5+4FuyC3oIDNmsJfNBC
GLqUMGlXMwGU523gmVCLmaOV/Erkq/y4HTRi6cS0RCd9sCGv+voTiwoD0GE2v7OD/bN/ghhJ7DvB
JnWRTTPScxMOOyO+UnETh9Ixgb/FRJ6+ZLlSmnf1mtc9skC3pNnI5sNCxp2nJl6VHjnU16b6w08o
fao+VQ/gaUA9JlNKPh4tZCOQ+usYTIGqirVzXnnf3yhSy4mvm1wYMU6/oj1/UkxIsdSKM8MC33mt
arxHFWfdstAG/jjfMEwsBwkj5SCxtOnyZNlYrNVtbn2trhAjifxhUj7WjxyhLGFGvnoxOS+fHf1/
8GjIyy9LbjDO1Nu4vmUD45Y1So5Wn+3lHJRUM6lUjdIETm4IhjPvzc6QpQItP6yex/2k+anNqT7l
tGb56HM+RfHHYDvK+qXtDHbz7kUy3hewexI3QyawxiOXaUXDNfk9Cfdlix7wlBLtb3GVedQOL/Qi
0QGAXN4GIg2tcBh3cJeEx8LPM9FllFjbBBIz/LkEcxA5AGLiVBt3xwwbrs6W9LogoUfeKLryBksd
QpCS5UuXduA+0zGV6vL7HW4x69xOf0kcTwIh8Ul9Qg3s2e6H15BXXmNBwnj82dYPkHQtPB527Nm+
Q8ckLbIDoUO/g2tCg8bzOsYbZD/IkwhR61P348zHkXqeq6O+GYdcta9KuSdSa4KJxAe+RDu0O7v+
MgYcAn5zI1RUaeg2l2TShPsDTIz1Y000PBt7tq3IUM9MnRphvzzP6aB/k539yo4xUrLbWijmFDG0
aIr8t1V7zGyzI8Ba3rzzp29hCVu/VbMZrD8sgir4ENH/uhgY/T4jV88MI2kaISxYcfnX/cZYuZx8
Q2eXxxU2Zzr9Fca7F+3wZ6DrQCpNov5Oq+3QMC1bgBBAcLOYQ/zjP2j4I29dJaqjNGuQPW92muR8
km3v6mQMqwXETYk2iNFcjHbkwUtAP7FcV3oFn/X2W/Ee5ohgkUWagX/u6NHfXiKPTxq7eOyGMnZG
Fsn9kEjfLCik/46XBUlghf3HKsu/BW9x39gN36HNTnF9FURvyALjilOV3DZiMfFYZtCUT4vm4DkG
rAnZsbgTmXEwcthhmHsab+2KL1rp0P8PoEJmaKv9ERs0WY42RKqUlC8YZ9H35db3wnLGOWTllcGJ
Gyp/GzQeNYQ1MpKG0HLCwOF0vnBfK0pah/bQUfWp9UBBratKc1LyLkSqUC9ph73kWFcppajJP79V
bsqKLw7vzMjG+PXwQA0Moh2VOR2RNcGi3Z2UZ5RfQCb8cRp56huINuZ47QyS+1Oe/jjd6xV428hD
QORc+7AzzH49La38i0WmaH5qoWb+Eki1eEKmYC9zrBylWJJQQXLxbzRqTS5Tg4YujdtgPBu45ctn
+TLj/iyPkRgJy8KmuCaDiKJUgWwm5rXUKq0XW0ATgbx+Il2QUgMXwtY/4LNwJlVzq66enYx6b/c9
FSxsKQTbzho/RzRDF1jK3SSu/hN09fP0u3eApPx48EBaMTjUzIA8PNfF7JI30t6cnaM6F6GAx1g9
5HbXbcgWFQC5umqk7XkW/DNvbubkpKM2iIQogmHBAD9crTp1Gp6kQxMBcIf9T8nWHvm1Nu3Tg2ol
aISB7vB5WEWXE6eBhVi/EAuO4vFGInOX6yj8uyu5cYDLNuPGEf6EfFjoppFB6ci3G36oAoIOW4N9
gc5lQjoe2YKlCgaT5QuSPdWO7HaINx4Z339ltVDjn2h0sw9twK0YfEZNV9SVmwd8GymLT9mwjzVC
bhngaU4z6xKKbsFg9uEsRq4UPtK+YKP/1ZzvUBwCFpkksssev+WcQfB5+SV3op6c1h/jkRPS3zKr
xTBoGEAN+JPZA9CvO9v2A286RgSdSG5b8+KtPq9MJsnvWB3FXkIKvPltIxvdhA6tjDr3aDicvboF
kIiWC5Wfo9i3TJReHUB4+7g9goidi4uJAp6kwlTwLlqo3q+Pwd9ISdxbbkcf9bJt16L5jfMJty1m
2fOXpSIR+LbRZR84yyzTE29WfJIBygf3Ge6U0W+sng2wRBRYTQf0wkT9E/1SMONpBbaN+aeI3eFY
fJvU2YmtCFe72rL3F9E4aXqRf8Rd/+n86xDfxFUVRtrAZ26agy+1MlfAkRHAFJEsrzsoyEKE4ftd
se0S2R3brGBF8kNvikxpXDCO7LdMshTumZyJek0FKHpysYNSh+66zTANdjWvQqCylWN5WgRTiZjv
BojBmH0iWez6Isg12J/ErYOjGB0q+YHCsG4E+oDz2gKU42GUjaMolyKCvf3ULovtMBZdRKrOipgd
dvPhgeH7Zaublu20pQK4u1C5iXtoZ4B836v6dCmQuyByJwaez+P05muGxOUJwPZR8rg4UYwfbBE9
5cnb2sFGYIBPqnFUfAZuNe5I9pe9CPAxJxpZH9VYaz2Wq3pNxsUHn+Cwc0maQU5/QTWnD0wJHy1j
2/F7eWOlNxxyt6usJKnFXXz5m7IofIwQTO2opWj0pbiZGjj9Ymj329R0zfCuPzRNKanlOAvmd7iT
Kpxum+CUepBU2MmiTJrLOpzMAyTgD4LfEEY36FPW8PyCRYvTALJojsgbAOr3dSvwBcfKI4ScRgz4
swBv5iQT7i/L33KdpAFaTT+2KKOKDar8br/sBWFMpLYsr6OgmZcFCzCkAkE7Jrwv1YgFtdw7G8/d
rhP2AN9bn6iNU1fzCOb1ASZ4tBZf8RKrkNFjoENq06BIFApdvajAcKqNuu+BjICwaVrXu0x0X8ZR
qGarj2s4gVF2QR6aYH3Slp5gvPoRqjuT5MmK50pSiNFYw5jVh7OKhDCq9zCgRUmG1pl91XizXYso
aYOlWpeFkY2LwFeihHzZOWbsKQ1MQ76pnJ7gSiKB1Ps/70H0w5bWHVMUlE+Qb7oQd6qJuoi1BPXn
e6+bZedAq6hGd8HCDu5MIOsZ5wrqsEMvoX3dhb6e+0n8Mibnk4SVXbY7Oq5FAtxvyrTHdMVpPjCw
wFcQTsLWSwlFQR576YhgHc+oAvGFXyesRVvmcC3xRwRzUEQ40WhjAE8jtV9UYGVfYri00Bh0v2vQ
52iVF2kyT8m2HPX0YKAJGiR0N7pfeza2FUN048c4KYkNwV0v9B0lQ+ipPRsy0c4kVu4V+fA1kKzl
FQJIBvY9zqVGhG2dzYfX1lTSSYAmzU4jgCSOTf9MCv29vztH75V/+5D3zEisy6ORoYAIqRxCoxQq
aNzRn+FEeJ5WpMCDTXgEjtkrscRRRKUgo08CvO1HC7GxXdAoimYj2niwU2NgZNhXM1LGD1EPK25T
iiAI5W1RojjzvJcfwxQCuMf2HXwpEywucIZhoWvYOkdTORcdh3z5jXlH5+pAgXK5rd3xYx8KZxAn
W0sF/YVjGN3HY++LxRnDynQ0i3bAw/j0avEr5ueCgAnZ51QPYmE5dFu/nMC3EQsb1ZAPc39fMXpZ
nCjBrTDd2ybxjx588qMKOPgsjzdpEf/SuEmet5m1xemS2kOw4U3eiehXGXR1r3wEgTaoPZlDTTI5
IIJcvVoULLz5xj24xr+71fHzIOFE/w9MJP2gp/rm6JmZJXUGqBNuyY8esNk4ehzWDlS/DZjHy98E
4vYSertizCakJWQmYy5C4B2Y4QayUZq+eoUS/MKd/h0fp8gX6A66WuZoWRSoPCzEDV+xvfU+cfDN
V58cqa9YhqiXJbGgfl9kjqvAMat4OUQnlGPI5aMyF2ARKiyBUorCAgDFP3M4G3d6lOKQp5wUKl8D
xjCmhAADlDOyvubot+TGM8EEQ+7fhIM7ADtSmGlCJ/iUrRJ1FB8XqsggoptQOYI70x7XT8mYPVoN
Zv/3m7hzuGxbMXQHWnf9Db3y7u1i/HBECougbLeuLl+/wJ+OSuxgL2/2ecdyNQtUIq09/ldWLkv0
8kX4RQvZH47yUKG24Bcog6aaSKE+Hs/QelcVivmA5esFk/v7UnSHLK+oKPnEKDRz4gyvk7RK7Upa
QbSPWJSywd+ZYtMtEg8Fcpm08eN8W0yFAIkjaEQVg2uh85GppB2dV+u5UGnHlr+NKIeo96BxFwWS
yF4xlYcluGOyMI7E4pC19NlIXwS18Ag3n30KgZp62MCh/ZBmDx8Jnk5E6OsF3XhkZi2mOIeIk5kI
HyaPJlP+vg9Q55BUrcyTthgodE3pVwHBQHdwA++YBZTMK8d2llzX9jpZixSIXBlQgAGds3dtRfAT
APf1L5OP2TBlQXvdHmwEZQANLYRDC1S4Pdcij9JcETtRs3twnrzGo7+OkLbg3m0VzpTM2wNfYNZK
3BxfIN5tH8G6KNBoxBnNU0/+vui6RyVK9pPAAb38KN4c0cI8wX+N9gpgnkqrxYC2M2phrT6BDx7t
NQcKKVBbbQoWsjxytC388mNdvADfJ2Wx4qkb11I+GXRQ2B9D22GAZFsxrv9Y/YxnljP/hrfb1vQV
KFd8wWiBVtpthHVVf5DnKCz5OUJRfCdo5yiwowM/XYgUG4tVj6t2Pe7P1/P0LCPUyO85rT9MkmbQ
WCb+1Gg3F221p5k3m0dteh9Q+etD1SAaW2qr9XZgpaEnFImdrUKhPRPU2Za6NTTcgOzXRBzL5LaP
WFVAE7f4nn1z9LrdubrfVV9e85blDI2mSCzOIctpW0IPsJFORKbaBOutSJ2X1OIRKBGvEjUgyn9U
TMmCGlXNXzTDjvpD/gi+fGEuvzYTkXSvBrTvmpvZyIQq+C0rALn2q5D72eRfBa3FQVNOiRZRmPwB
1B+5T3vmlOG8y8bS8s5wA0M47EhP149BiQfgkVEjp0xwEXNkmqRsnNv4vwFZD5hJGPIYOQZ5+aBk
YgF2TRX74jcWN+hJlIS5V6qQLOx346WPKGu55ygChZqqzcB9bQq/YQbGLWNAQQ3uJq2M5STlTnTT
QEpPd5daS1fyVTe7fnQOQ7WWsY0w3iLbtwrUzLMnUQF+H8BLncEbpHybrfIljOJHU0ZaqX+UuyEC
M1LXBntqLKMZjWqqyRlq3/5iKr9rvzy6nKU+ZU7mpW0lG01SPCxZF1fnTrsIQEavarM59KclxJ8P
Sjm+N5aLzK4xoLA8tKI5H3XWAApNu7I77+suthiVRg2pC2uGL6yKIzfGHtpJA3SB+h6Mgb1USgax
j1LiL/WYfDotzbWq/TO9FIVQoqCWplsYmHsXfZwKbtNIet7EJK3WhD9evxzvgRlWROyFWPtrfRFp
tEbv/Pf0rps7Uh8AL5BiZVX1r82h78ha/LDz1E0qRTipS8ZXexJjH2yaqyUHPtsGCLaFzVy43FgZ
IxD5CsBJlCFo5RtOaj/XFzWpJ8ffJVmYbXTJzxQXxZBW3lXWdoxc/VonXMZmeihyl85RfqiPaZPL
pRacJXDt2IerF1I6xXy5ypxvJ/d1H5FvhbbdY+vPWTpubxyA1EyDnHZvV9nB3o9ONmtnCvKkrsoz
s+NCy9r7GK0qKJj2o/P0YX65skC0TxO3aV1uv9kgepq8ShU30BnlexA/6yWaShmsYtfrXGe8Zvlj
5QgiLFhmFNxLrt+HaGC+wJCHeoLofVLynXgI72AkMyM7Olp3FCVdEKWoyOpAAyk6hW8TNAw3Tjjv
JcYTGNuK7HIfLi4uM6qhzXAKkROP2dYIb6uAmA1p03I3Fe3E4Lc/m3JEUI+g6gpGWEMaFI8MBHYU
HPJMNHYl+I6QjwO7UQT/Z05Bp0JtGnAd/HHYyeG6wQDPstHsnQY1hbhCoM2/0JXuKoNb5y16YAIB
RKIuJQxx+FWHWRefW76oligeNsyOTpw056BUiiOy/quw8qXuwiWr6ri2bW5WUmh/GP6Ple1b0eFR
1nEpA9fqgPkqIM6TzcwO/nrmVQQj5+A9/d2Q117bPOKg/AqteHrEuvxVpRV8iQbma+YX7We2kY1j
nvBF3qQmBxABksLsKV32UnnAwbaTKOF4Y53SpdXbxd3d+G55tN/P18Uln6mUMLT3iz9aI4qbeMQI
XtI09CliVqArZpI4JxVeXoDc+jtmF5Db86kpfaUvs9nnJYSfFkJ7uo7IWqOwfz0i9OMIBGM8/pef
J+lXPJR+zQjP7yT7CqmI6AKvzYgEyQx4AEAY2DV3GEpSWsZfYNznjeAzBCukOLBTJKOXwzI2z+PR
IyYUV3K4iRZWxG6fZZ2o7qHaVQg+DTj5UBI3lfYRY0CNasv8B097X49qlLIV8yQsqfdXXL1n8Nho
cNy7uW0y6512NChg2WMha2DBfPh+LuDLt8TdidihQ8SZAJZ3OoR5dRX6mVbcsVY+WLiE7bRxxjDA
dQmb/BVkiMxYg6rTM0CPkWEYUg93vYy+armmu+ErChlac4+F3CAMBnCSpPC43osoM6AZnSWHnsHy
Hw98LqKRAPRCGy9hi5wiMoW86/Upr3gMje9MmY0df9MAhDYIIpeLieWhTM4TCme9z7+4GAHDRPGl
uyqgi01PuvSEqkj4n4gL7LC7sH8S0qaXb0SU5JoHJ++Lr1XuCosVYNryITho7gpPxLGBf0CopRY7
F5zKC2YuwMqaA+JDEq5iVUh3YAL7BFbW/21+8ZopGhA6DeCrRvHiz6Z1pPERrOCMijed0FYOyaJs
HCLtTfLTWYF00l0tIAnWSFDy3LjHmvsZh+ltmZQZf2H+BzMCR4qZbRySL4cj8w8EtF4b5K5zviVR
5kdvyMYzQXJOSYk6MqRnYUJ94c1XytLNfsyFF2HkcKIt/Qa+s4K2Yed7+WSnKo4rYHt/QxyaEcq8
kJXqPUxOBSJJOh2LREecFOI17EeSO+k1luv8bRqwIKilpIeHxA4tS42DZTYGjTF+4xaM+Pvw7fuZ
YSUE7R0DjtajPZvSxzEwGQ33p9F5v1LVGsHjkdKBn55/JBHCIsP0dN8dEr7oO2gELjtT7hRcvvsp
56Y7nXJK4TiOf/6S63z8b4Xa6iMLsP0E+IGmoKUXdVI5gWMjuA669ube9UESZZy3o1QiGGegFl5v
ngvuAEHkgJKgBlxZRmh2BddgFWued8z2G4bw7cy533nX+RBKvYna9/hCiPcNeKr09a80PeRyBvrs
q99XpgFjD2G+bovpu1vaLzD6o/EdRPNoMZHHTyy/aCTUkTmcW6gCB9VdfKEx9O9kUlWhP/EXor55
WfEEf1kLE3InpKGxKQ1MtwOBybf+KEVTMGsyAXTnIqjBTMJkILHlt3ckaXEMW0ASnr0BxljpyDxn
rQCMSDNx+i3Fha9hYZLFCyQZlcD/o3Ugg78I7FalO4Z2VDTACtSFqe8ZVYSF3nqA8/JucPGl7c/x
4kiymzdDDLDyHm2uDuUroxaqoCuaD7LageSn4mvLL/1FXBIa2z9DuM842ypCxi922GgzdvrwjyMD
TWI0FeuUYAlr6AYqD6baanwO0EJYteiWlRNmUJ3ccgsIYBlx7/CR138O0fdpRHiD6SrC/F2PUvfb
7JIWLvgS8gxEddejUGJdEi607ZP+JVM9pK1kA8ZehyySSVY0FylWp6BS471hhI9gGFYwM6sQh0cQ
ZeT58L7ELUZnJNxYIO1fsJYTSeaY6ap9lBr0+7Gy0USwaO3hadjTHF1q3cHQbOrzd6BHPo0GSXnj
bEzd1L/5fEJRfyrdadJwh9uILNMAzZIbsT7AbOFEodO7GpBY24vzXe+CGb8p9M4J6qnQK/vNW1km
LhVItGDL8lqrtxaY+Ydez7zWbbcDeR3OrDVU2ypsvHSZMGMu+XdoTFd58WeT64705pi3EZ5EonHq
Y7+lecYcVC5zwe8htXG0rG0/aTgpB/jhHtU0Ah5MyGnICXsgSMUt54Pvx++PsTmqdhob+q2BD2Cd
xCwHGxqhWVW9oa+7v/kdBs2dmkVakHxZj/7qI4Ur5GGZ8JVy+6RDB5KjYn/wuLTllDGGM1+yNdh0
d6RLqkSylIjMoinuUOx8+tu/0ydI0rw+yH7PFSRqQDgDXsZkAD+/OT1Z37yFW4bsCVR0M0BQ0WQr
PXOxu9NyjBMbsSwKkeyCi9Dt9Qc4jAHBiXDzu79y4zaioL9egJVEpZmefkElovSNNFaLfrXqHu4b
mZeduf4EVumjsvRCDUUpRwNR4baBRcM+5ugPrYWcpiAQU9hqAQolNXGTdS9gJjY+8aBT/ezoXi0y
NDQO1ub21EsSmG7iw5TLwCW3tXX1OOXyBdo20Z0ZWxkSVcnj36jEmBWA4YlFN2PYlPhZcBwD1J7M
8IEtO/VvtPja6zhQ7n/CNunhayU8zSzyfvb1/T9ScNG3mE4FKkxZvWnWvacNaHjJ6j5kE9KYkhqX
oBm5QsXHMy7/J/8Ft98OSfMmj2eYWYcxI16yObLoMEx7UNzH2eItLpteLLrfEN9qXby6M7RQaSSp
NyOElwmqLCcC0reAsoaKecOSw7ibi7HMBUTmNUkNA1NPNGKCIAzEBao5QRBXgedpxL8nXWIiuLHP
BGIvLJcZ4c0Gg9/X+tv5BSZSDzBVWPjn1WdE96qlCxYwZQwgK2PZTfoI0ahmXvFc8eBMhU60qaii
2xTSw6AekWFNr9RQC5v+SknQCuMgc2BUI7opO8sYIrYFPxiPmd8y7IqmykHZ3X9gEKzjDE5QdBmM
aW8j3WOeU+8bY6DJO+RH3ZDWhr8S0Ga+4hlGEJZ9va89VaCJfbJfbaaQUbAa2S+QB69nMfQGlFmT
5UG97VL6vbOdTbIrI0BsxtPuHeQuMJOLJENrL6nmE7YYl10sScH3hPmJNoOIj0dR7g0+SZ/nf2Jg
4xja8Cv7OTT97vitQEuER1Ui6Zxg/892YSfebOH/VoTfuDTnP8pBTalGRWO3YyLbaNM6dlhRIiAh
qWHXQ+fGHEUBfWhXve+yolr9IXmnLMdFHxZO3T/XImkHBMOHL8o8JTPJ/mOF/aGBxINydYoVHlFt
o7dgBaWXsWwYaonzHU3cSzHe8grG7qzAFMQOVY39Qip4OjuMdoS+bsDdL9ZaYMMVcHCkHVv8CLNk
o8Oy1U5e92BvUSawDEt9dDMha4SO5GU/TeXGRXzVK9/jh9FIH1lKmDLieOFe/k9umBj5O9y1knnx
KN3U7OHrqKGCh5FRzeVjhpKoCHB8ZjLdjmPcT6WOyxVgMZGUkUd1lX6ghg7FrND6c0yN4dVCUGh4
PR8zna7h1xTC9Pnl2hwot0nU1+qqqHpBc/4biKilAcdwLvyqdraTEEMfCCVptt0MpemOOK1J3Ux+
f0AwqxLBYrghN+/nXAg4CLIsHWwPSFYOFXEUfVl7TBlx5wHOevX1eD8pzIX+pCO7ldKzjnWpJ8Ms
eb5KQ+RUWYwQuN8VQG+Mo7MK1R1Ypq4FNz3j2gdcAV2aNFWyGUxzAC24lbWOT6YdjlHpTVbWtyf5
sdtbVrhXtt45dKHBdwpdM+S+zn05uSlVLjDPDyD3XCNEd19JrMJjnSoMTfYK8H6xDMScV04FVsfT
sve780u9FIzGmTXNEKPaVjjjuE7cUIeQCni9GaAimXwekEA6zMWtV7ZdhwP+diE5K+IvjOsRKEH9
LZBsnc5ujIOLWyJnO2KcPnEUdwxtoDJDm+c6VveU2PevRx6LJfh5vJEYudnP6y6adYpRcIhpnHcq
hwyq4+NEY7aDMSUC/q/5yPfwPCPpoKhiLo7g1Z4UFFpuxeSbbqh4TmJY+ffR8twl/Z3bZq8QHJTa
yt44cRtSkfWos3mcOWIy/V15ypfcVUYhJG+q6fFK7RnKJ2tTj5MNrjykrUCI13bm8+yoDvuOZlAN
lRoPUrJe2qeNpnhthYwUzOnCwBsNayTn/aZM0vo+rTOGl/bqQNCIxows84AinOcAypptMMbw+zKM
BHkZLHkrpklcgkyFOhfTFdHZeEaAEmuo98YFMVyvUKUWk/Hb3/sVAGl3nKcl2nXqglyWdEFvd0SG
dH+58zhplWDKRzWimUHT7gKGuKM05Dngv7OeO0tOGwyTi30h1oiylHTXtmwNxxhvlval2YNFH43F
oxORYWXJd8UKB500Jr/mwzByCA56iwmRtEOPhm+2a+00Q5gKuKI00p1PzdYlrsY0xm671MpAI/oo
Yy3/Cdw/t+i15JeCG5FNU2sE6aAbTsH3wPYujCAxw8Yf0GHpX0zTdjdzPNLe8p15FEwEJJ+Gmyv7
KNVO0m2RUkhP5rU1SbhauVJeD/2Uva0wDrOWJcqHySuxZPDE1eMD8LchQR0M/P8I5ciy82mgcuJI
QN+yxGvw6S99YxEwJWpPsiFyKOMFiVwvlI0CzEnt7uGC70t6CP3Fu04VdT9GYfKQf9xFXj8lOyDb
IsWGMz6X8/lHzC5S565jaCyGR0zBUMoeRcVFrsmelRqzjoK/2MoZxiQcTkEU3NUX17JOhMUmR32V
4o8djHbUd8GBjx+KsfXP9sDIpNxQgRzc0VineTLUm0V6bEVStSB/VQ3f/1nxr/RuU8t1dYMvuRdD
GItROePRKeeVR6bgYq7myBAFYo3aPIVZYnM9+0vZ0yZiWpQHBNvXt+Zt3YW005cxwdzrk/0lNsoj
r8AKklp/BDcQbF/uFMNlkFDq5M9qI48sPkvXvlkwHVC3VfeC1Hndx3dOpOSR/3NTJujbXwio3GdE
4VPfu8HlVLk39BfPq/reNoUVpb6YPb9GI+J1NcjchVvKXJHdzGdxjVfa8t0//Ejofl8MdMS5MZ9k
3OyBGXjA90DOFcnUkuO36Y5bEUMaPJul3r6b0S4NNhHVpgJeJUfj1igKk3L+HPdzmx3TlStJVQi3
5HIVqbzz2magUz7Sy40JSqoZhiwWdadv9QcsFu2JwRp2habf3ZtOjX5vz664NvZAE336e/vJ198Y
N3AxzbPaK81N2wCs1y9+va47CGEiyWRYbRa4qkFeJRAkwapf47pS6oH0DjekHjrD3oTzKOBZZe9q
OUFhgT+uC2ZwUDdlTNFzlJKPoCim1cv4bAoJ0YcGr6GGrzDP/oRLH9kTgDAwn7gbPNHrlscQE2GU
Dw8WywIQ5CSDEVdQV8twS7OcUSs9YiFVKVpWgguy+fngXWfzc67MBC306PiM7WuObbDNWcYIAKq3
rndrSGF7Txk0StUOP0qKMOYLt+5gfT3inBYWMWrxDwyC99K5oG6h4prwxZVEyQ8WVPt/Ofl5W3XH
f98eOdN4JhCu8RIWnHMcvtKgMBnDSEv0gqTfjKH59lFQXYmnJp68XNw/rlV78G6r/eVuklUBbLtn
rej/vp8vfT46YdqKINyOI2ai7FH+KosDdo8RqEg7lqGU6PFOQbDcQtbB/XsgVharlv5RVoWEYcyc
1tey/80oB7obN0oQ8arNFryI9GhXqGJNkFiyV6AZoN6exkgeybQx+YUrC5aMTr6ynvpW6lbO42Hd
5cF79ldzUXvAmV2pYVS/IZ2V6w0Gi5Ld0uXliHJneWv8VOTNevfuT3KvcB4BpcYL7Lmf4qRanP3Y
ME4RRrwGUoAHuJPtWFWH8hoOXpsR62UBxqvroG21JjnnUnLfLVq0Tetv/5TOoUz1KfFmaJzEqBOz
IctzoWr+6Fw/eGTiqrrM8F9/D6ywHwCiiOCaw3Lm5gLM1xRHio1uEkW0X8xVhm8yESVQcuTYpETY
DLJECTTMIj2xMGnj6rv5FdgajHn0tt5gvQYAVwkfem9SeDBR8nIlBiMTixWoBJVSFtMr/6+Jv9ur
renf5ukib50qYvlMHCQyRTTPpF3dCEshmEq0/K26ZirV8NEz7sTXbg2bX4df7vC7ghBrh9MKxHxN
ku+ioFS++XUWGyqm+cAfxAWb6mZLi/emcDm/CHjwqQbsPUKnOwko27o2jlHEYNdQ8H3eQqtsudnh
tU6oX35F6AibySHAb1WmZRF4b+qQGgbbPHka1+ZKq3qPUmh5wVRCI14x53QejoQ2LxsekOvqf1Dd
kFYXcWLHPheRHFiY/Tos2S7JRUJv0L0Svgo4BIhtJ5iECA6MCoTdI8069WFc2LPmOZy5EHsZ4Z3y
5+ZvGpGwYbJ0aG3vceLx03sDak56x9KbkCthtHtzSsBDBDFcw/ug9fjdNo7o4rhWJwYnpKV2TIMG
+tJS1IC37ZkBH3rFum9Q44t9rInM4TabSB63JHcboX1RzDQP5vg+uZxvZZy80ipt8T3rKfMkiOJy
vl3p8Ks4spQXH4uLc8mhbc2aSLO85ioKjfuFnPnGHRhVKVL2jsr8K6z0r2lfI7OvP9wk/Bfols6W
Te6OPQ+TORKnrpBKLRjFZgs/JfZQ+EJaRoDKnMU3itfQtfCcpIh4YiWuh5E0t7Zmf6GFYy5lotSa
hUtdVGPZlJL1m4o6oeDBMfEFaH9P1CjtcOtk0A9tsCPe6r4V4S2WCvyXTIFtthR+f8CA+1hPbLMJ
KjH6/FFhs5Gy6StN1jawSpf7lXXSNL1qXKnMZMZb68NoSNidvbDltBSh4c4jT71qrzV1qG1cBN3g
ZKlfgqdWE5gMkHUkOXc93XPTIqmHu341xmtjvVv4EKwUaxBQZhE0Bn0naMMckp4d9jTeCCrBzYcA
MqyzHVJVilOhYfaWyQL+ojSFYOzUKJtogrn7lSifCdToPtl9ksH/NRnpn5WhpuMTJe68FKCIIGw9
WF2NyjWnryOuj9iL0nbIeq8eAiNY+ZYYDeXxHWLZaytPrKVINc9UkBFfC8TowwVkjgGPlx2dl5O8
GLCVoAAZx7R3HuOxCVuDm33w+KBcNY0e41VJKE9LXQcuINxPJtGABDEyfSHRW2vwcCL4vtq2KRXh
y9ikm04uJ5CP1jq7jF4qN/Oyf3JwEr2EsCN/tZP3kC8lpB5gKR6fzmyzAW04lfRoOQaz4F8I6dtT
oPS0Fa/26SsL4NZUsfSz1DXqhJ0KlJVQOb3JHHTTYlDDhMWoe5QePTfW5sAy7Bmof/gswb1BcsGd
4i5JdNLllK75iOAwr9BAsC6T387izUr73yrKAN7BRKyFgyGqYLH/uHM6LhtwMy/WTCFKG8YOg6RP
bFFgJko6ihZpS+fzFb0AFct7xQQvirrC5OL91VXLR9SuO3aMBrM4uxw+CLnp4qsz3UzkuJ5x/ASg
OxVRfH6yL8VvVCDftXsZ6MrkUV4Owowl3BGBA31ISpXQqYjbGxXW6MN+/gc+/UABfUQ9iSFG74bh
szQDFBq/K3Pfb/ufjBhmTPaLCju1PCYYZhRyhZjJXzfB950miOlvzxFKohVViWikS+rqPM2zQh0S
UvkdC6kpk7p61DsM6aUDDdxELSPAaf6dv1yT6nRXvmPHSqmOzUsPJsPG4R8cwHx3aO8Ofi/rr3oU
IU3nK1EymAzViBzwIeaoewB9/wh0DxUiFVOIWr6SiQ6w1AISqFemh0bpO6s7rl3cDNHrZrA2Q23z
7s5zQlhzPi9lsh4qsI6cR4G+iPLm8+WbEvwJmi0Ui3IxIL2qhlpUB/nSjXLCELjknI8isF5AgHrL
x9wq+xLkQXS9AzUr7+k3bbmJjtbiF/xeCX8JRq1CwybFmBgb6iz1/xSGF7enrr8a7dcbc4wuvfnX
0ZHYDj0JpMaRfol+IVzE9Nd5t5bFKTAc4u9HmOj09Tjjr1UQXaqChWiAXlICFCNEITJNcbs3SUat
hqd62E6lhtCv7l8SVz4uPRnJLTT/FECq/7qJBsg9KfOiv80Cpkjlk7ibd6s/HhlDN9XJxffEc2Vs
LVQS0YFJF5oazokHZUkMGnDfCT+DYKcyi20t2hnsVlCFbVbDHYFdWSLwxavRbpHi+SduUBTjpW/j
QjwR0lSRKbYevXSgez7ATyXc1OxBi0JmBLszN6o3mVPfeowLKtrUEaiy4+GvfA7nfryMArTwaYVC
pnxoDxa9eQfUa+n4NNCmRhYXsT1z3kK6n70kHWpimFq7HzphUuygqdBPD1ZUiuvoF3H6tj4kofO1
ZJG0HRMeMXe/xbNaWEcINv8TMMoAXAO9y8MXsbEr6910+KvCmi1MX58nZayjKtUUtSyauKaKPACP
cvvSC+4lXE2bApn4sRehQwiPJx9JtMjAPdoDx9YAL4zy06R/K0aicv42YttBg5HyEkbD8LSvzJsH
pxs1NqGANfdxBjRKuo8yPDoFIUyTtlPsRH+KALf0mJ2Fhv3fwkeZySffwNtwjHf1dFmAXdETDxgG
mFsVOMRInWHjX0Nnbm4WfKk/Ki/D1fXRmlclF7v68eAL5Wnj5nIFWA0R8DykRQT8mzU+l0b5oaes
P4DGfT22L8lmJXU9e0EfYCenSXTGL9RQN2Y3hMd4b8vRKNWWSUsC2za4128AuaFh+y/Tms0798/J
CGXgTFGnKzwkKatCHvl04v6JdPjHX4bNaBKqFUXzf6zEr+5mfHu8QnVJt4u7o1Urrvb/M4q8tNcu
gUH/XvRoPIqCwA0flveFvY6/zJYQPiEeatStxn1aDC0QD6OqZSB6siWywJqekvs9lOdeELJ6MV4T
IpmmpY+69Mnn9ChjIOiSHWl88oTKbwo/dkdBDJ4lQzIZhuKV0t1uowSXeQOU5lRppgW+3W2+ePxc
7EQazvVQTWQ7lVn/zTk4kGIul/tze9lPNsHpZhXySNNBmlS5OnqyxtCXjnzbc7zf2F80+ft2WBuu
ACJmt8K3rR3hwsxrxLMZYbR+bicENvAJVcMiPju0Lc6Gn/kxDY2NnVlkjqBgmsxw5uQizz+E9JR1
k8OtwAZ2kt1/p2e2gMEtqJhadOXImG779bXxutA3VSSOCFhrVUyXfJzoHclhTAIgJJ++7McO04cF
0v6iUSEtPxyz5hK+3OsB+lXwBlAsmle/UZk41NXYyeZNXZnEhCG1try4v9V6B/B3IRJ20sLNC9jh
Rr1dHPRlFGYSQhl63rEKyTCMF5G9ltqZ04JbYNEDW+fqEJuLKCwRAFh/JeIZ1kJAn/fGHPKOgA1A
+Zv0wxEW1ZggdlDpsLi0U6fHSyfof57gb2r+g4PM1ZcaHiKotitT3jmejobeMjV9rcHrO+aXVaoi
tna+RT1Dw30HqKxRlRJZcAagp75R1C6sD92KKTOKBHP0HyJ/7KpgCYuHgRDY5ypppxNTGaHe/AQO
27tVYVlTgGKP32pxQN0e2c4qkHbQKkibkfdJs2f+i1kR+ZjDgY5eSCtzeOx2MncdPk4GUTrs9BiH
IBm+yS398wnOIuNB5wuuOJN/8ulJ0P0AaHRZNx4SycXTgqu7eQq7IoZjP0irq88OiY9qdovaCaJD
rz3+MfUEx01HTjEcv5xBkM5pfEiG+E4wDydYvGhbbsUdRk0sloz64JxNu074xsHMxigJy+0/4tPG
2BbYlawBRWCATej9UKTiLhhIENwYP8WK+2hYMB/7KQ7YB6qklyMATTnqaCQyeJ4UyswwPWNME4hq
vS2k8CoM/fRbuggZlg5sMduji00EyOa5HVpHnzt0nQ3kg0QI5wcIZn+57vFmfIRfmq152dV/uizp
BJ5tFjQBEiYku/mfg/uVw1IE9w9/jA3XGel5/4C7HX/v/eSgzqXsCoXyWnTSsBaCBEBp0hBPbS5t
E+arjLtNmvu5JBsfy84ZntX8U0NyyKp+hpJRgpnwffYSPbk6IiOthc/q9kvNMXGZiXDBe/NwwYfK
vRuiQUgQPj9iNx8oxrSoltAy52DoyzEJz8t5DT8X+T2clz4+EaxV4tQCEHGvd+V6clJpwi6TdcbA
7wp1nKcMIaPsq1JzUP1FAfHL0Z+5/B1tvYKagsWFjIxn2OurNqbMzuY7yoNC0Izbsof8iU8E9et6
EG9WOtYAqICUWShXq9FOSNMUafsQC7fsGZIMq8/WU1vU9O5mRMgknXzn0h4ujdrbJZe7jd2/2DSQ
0UptfsnGUZmxR+LKyLB/NSGM1ZRHkXzZR4FNaTO/f3GyO7WxbOMUaKax0xgPfJMc0dTbq2/6gVXZ
GLhYhVsUoDkrelk7Sbl6MiuX/Qygv79yoPFOomQijlN+QfbdqqGxIOH56Zbq7vYLsctUgkldYAmh
ZG7gabxa/tW0uCoEVghDbFx3+2RJtyBEy33E0d6Wj3U+Edr5raR83KwfzV3ne9jE7JXca3auQxkr
3LdkWel+mrZ5LvLemWSF1qn2RNDEfUOuFIrYwhPipIAwEBUHR1Wywxfy2p7a0/oRIglfNHYrioCv
Efekzc4QAeMc3l9szVBO8AbzWi291UxWLEUHuldS5UW2hugeFcryYP7evaRMZMhMaIGJ9WtNykW8
DFrqBAxBO2V+4LHKW4qRnc/oykXgm5HY2aBUzTnOiFp3eqiDpTyqgoDypQYFiEdo+7xwD3DjfIth
EeTvAkicEhb1IdAtuLDayPbMj4W9NcUkO5GTJ65GZ/Gnwr7vzVSt+RyD14IgNMJhegNBouckDpOb
j2aKsr9aWN5dPd2B4oddWiPpT1yyubzFL5QULcNcVc64a/vrq1xC3Yp5q5/XzbZ/LLMy6O4oMZZ8
8F3LgRJ6mYxZoqoLcvezY9eR8yWZzcPTnAny8rPRtshQFYA6zEm6Rtx4ynCg9m0xqY1fSjVQjSr+
+lOU2/E7bDZMWpUDD/OU05Ukaim9iadao1555FK6Q5KRGaxN3mpRRbALFRYEYACjwZZwPLGP7uAY
jAZ4DfjXWWSXMrVWr0WX0kVs2i/4WBtnjNykc9/jSFmhPcjx3+lzZZCguRA+cYD1Qx7fpXpoqZyt
Z11z+m1KhRakcfk57qutN4ukhoSkzmyJA/Oq1dLkYhwfUwIneQsenBvwPmsrv/e3+41lG5jpoX8u
yyLrAorDd/O78O6DxMJKYwpNaAdTKfmOn2hMQmbVLd54mw2jN2B7IMghoYAfoXhQw1x1j/Xq1jP4
j5OAInV3l3wn2e4VkSlejNwsFh2UhzATxxPffy2HgXzYLkqnNejfzVRzZlBeqNeOULg/Rvn5AcBx
osDUGHqqOS/Ap5cezrMQlhVMx+UFQD4h34oq6K6Mi7EMuYK+JiBkM+AUM/PiV6RBjTJ98cOtR7av
MWFwQE5Sa07mc6Wpd3KDiWFqrKobOcjx/sx2KFLAKG8ktCTR6l+xQccsm/TcqUJZw7IgZTjKJSbU
rRGe0NK72MBUER9ZvMjltrj/dL/NeABa/6gsZGoj1viqZJmIym4zwTRiJT8O0LnpH84agAx/ky9K
gLFPjkinup7HhKCzMGAGxYA0elPDE3yH/yijFkfHztrM8lq0KshxGbj42dUd+hHajsd0iqv6SKZ2
s0Ez+d6FnPhpz59gyRso73PSk4i6Tbyu4LeR+pMGbp+y3L81HLw+IMVvSMFM76TWjm8hQuf9BE50
fMpv4AdvLZH7M5U3fmj555ZbzMcOH4BOiI+2uVYkKSh7l/RuVeK1hJIbHmRS+OoyB7l/UbWdc14L
z4GQ2FCOGfg5MVwABUmvFBQAYVHuEBWyiaQDp4z9PTkzRB/XuQ84dNSLjy6UtjnOAt9xtc5XTrgY
Y6bdlW6VkNxlQeKmLY8BXQweqVhJYzWtSijdH5swlO4Q8c2vz6zbQc15mqflwcoPt4TlmZvxBA+F
KIoaKk3zaEVMeqwfljxOMCfvrmjY0IrNx+yPUbrYGeEmK4qooHJRD3J4zHROPsvzpzVRlLo2m9As
/MR0Klezqz83Iu9w3HuYzghzCsuT0j4nbpJIy1ynTUPE2+3rey0XzR1AvX1Ra5qLB/xHZmMsvNbF
VlODEdJKidokdXezmYGnCodGrqGobio7p4x8/6qxesAxAWWyN0rV76PaCDtqcT73AFrRoHkM4S6c
BjtzeKKHCiBMqNZMplEMZo3898P8akMuUu+el640AwCqN9xzEZMQ5gJvyk27/aItabU+NMCBWpJU
euWW2kg+psybFJBnupBKNyo0wg6hrRUCWuZ3v0lK/Ec11bkBWLq8i2FPMLSOm9Nt8Q/QBjOoptmp
hw3bfIb5Qjs47s4cgPInqMKXWQSsY23+6O4D+ix6Bww/McDZS0hb6I4lNJUOR4a1puG2QR1uK7Bu
kzDeXyyj1XI/D9AZGPVSiA4fCFo7TkImTieh9j9iKGFNRmkccgxQ8SM7B2JqmUOcJmP4zvM4Sbbe
HsSzC2o3eNx8VaedYGbfB5XMp8BhsL/JKGmXnyj6WsTxn+4IWxFwBrB6AQxwolx4HjV/LO3GKvfX
ofsbxkYxZS3T8Sig0b2s6cRCHp1/XAhNptHCRfseIb6gdjomhCfZ85772EXxkwh01PCsg8AWJQZw
FvsgCRxWuI8K1oxSJDi9QRIOmmsnyN8l7+vtGUkOpQ3ZYVVWHSjE8THWAo59/8V4MRRqJvSBkuxG
I8R2K54pE4QHwN3vtiu5yO8zuX64bWiyjiZz+Zmn4F1zYkRk0L/vBjrBouHNlhjj/DN9faozefNo
Jz6XrXt/kULU26QXPQBV6mp8j98QSwzA+gKz1plvRMOeUZ8cVnNHmLUgn2A1RYgx3JuELFJDuBkQ
BwrDGad7MWzapuuKmUkjy3CmRbr+rhr6m/ntVOWa7mKH+L7jvORpaaotGQTTOV0HN54qeTi1K09n
pJqS20JMplPij2QIIPBhiAMC5UMjSuk339VEwhuY1Ft3QDo1Fwvd1F/FYRQi7bDHWSIMR95jXrnZ
wiyyi3R0n41f1MeFTc0pXILdPWiimRD/7lMCQA+Dk0LCcuEoKD0fuHMuO9vpKOiYJ+IDx/4bRvLE
HWQ4UDNa7KEiVWwxGG/uk4ohoEqIzTqPSVIZjRalSEoevoXE3Qdf2xXQDFrNPQuPn/Hg0itAciya
/Y0YFtccZ4g9nCG6GxRtiMBGCtyxxeL50rO0Qgm9FHA3VBYX/0PZqBLK4lnlBt3Zp3+47O9Vnwzw
aoSZOAVq/iLhPuuTdra/UYNXzuudKKT2DKEzjHDKUEA8srR6G4Z8P9ZWXaH/oA3a+jwjaXwv8Pe5
LuHo3eByGcxJLfYMyuB2Vu5i4LZs1JmtP+N5d5inKd6hs34PSvzS39wFvj6FM7SCKadorH1dTWZg
IlcYM+qMhcPxxUyVhHH3uzszFLhS5TBEMcF8DoNMJK1pYeuSUUFfuMFMOMLrRpUXJOmePH6AT99V
Uh4gfdznalMzylycpkVA9A6zLDJQ3a2RqeyZKRYMLTb29tto7mM3KRi10DbU2DbSs1Px8AZY5aQg
XDFs2Owt97UAq+OD0x96moiQNWXSBVhS0gIaVVWpLhtmVWV+mkJqK+JIlg2e/ueeqeauqZBOe5z5
U9/xhnwVAaAcQHUR94C3Gz1FxBTbE7Wbp5NnDyUhFDm4tOwCeXt5Eixp5tFqDTOa2oUWaOyF0KVd
eJj/8OaZHQYZr/KVr0ULKVDsp/IQen8ltg2xSt9EVqu9Iumj5D/Hmz9FBE4CEfT+XP7Y2ayqvYkG
mQq65h30rWqArMLoa9zd4DtCyZOcxN+2gIqDsh0MOZCs/VhNjF8fRzpLZ/CTQ+psKjZxVwNlD4rd
lR6XVVY6a2bnYuoY2I/0oPCeS81J50cS8CqRZDTyQNXwyCqSF9JYECeSH7HH/zABH4MNzbQjXLG8
4uuljd8I/puq1ijUgiRgiQtoF7r3Zepwoqka3jowop4EkeTO/wxdha7OtqI4tzG2/0byOMWv54/A
To08WrTekFwUFxwBtXPgT07uyvX/91wO6cDM98NL2o1dqGBG3c62havDPy1JL92wnJaMQC/ko6+Y
Hgo44NcpUJyRsZ4ttM99iIYshebGfL2Xt+qKVN4NKCu6EwpnRSb25ZBbB9KELikR/fv4qYt6ruag
7YzGppFvCzxSGip4SBYhS7KWz3F+yx5vhfDN0LIDoJLm+WGmEdcqxAIzVfEf4doHGF6nIbtC0LxT
Uaz+bU32xFcwkGCKYXSQl7mj94I/HkiYnVWB+TQEY7rMykQkRIguKiESI3NGB8yOCd4bfX206JGg
Z0zsM3AIJMw9lSgPHXcZ34twJAHlbOd8YoLsP5EOsoZ7NFa62mfaXx6qgeNsBdnWqAM9kW4SoX2K
l0z7RDXQQODbOwNJFAV4Z1cg7Wx09+hVfEMyK5gKESs1nazPix916AiJ+F1yNlblb3RX4+K5R+kl
znYFCTMn2RRBzGQMwjYLFwDVe4GLw0hvTF7tlP1LP7tbA64j31Uny8GTBTlQDik1rcxhzno0+Lji
tQhT8XWlJP5IfxDG/caiM+PUlvpY5dpuT+wmLOChkYOl2HvRRqGO0awMDyXEo/SLoie3mih3zIaF
aKVFyPkVijNCzGauHVhudvGlLuxYM0COr6Z3z1ei599DNJT3CzuQZE+rUUGTdvq4RAEPBZQJdgTG
pTkEKS+6i7vFx6A9RvyRhdSlC4AZxeODOZ3UviI2pg37CkHJe9zV0keZ0C0QCyh8APBgzFrGrtFw
t2wcWh/kmYkxGCqjGbcx/GqDxI8IdlBwJx5Bafav4RSttdk1dhMco2+CWt8JSaLMpLKamhanYeQt
9iUi4mUaTyzcEetdmLVizMY9ejmW37Fr6po0V3P1INJfmq8VoJTQa+C+emjbOD8+GPuK1ZA1M6a9
zSgalFvDPX/JWuifMNT16eH99gufO+yFVzZPn0TABpDIjr5oQ1hZMRZYPaD4eL2YbIUe8heCVkIo
dkJeCyW1e390ihf58TbwykBshs5vLhxoeuDF1KCHIcZnYQSH5SboQKmO6PkZTMUQC21A/JoZmbJQ
DGD4xDw5QNlZ4T8LP7EiUj0iKMPWTME56Nckc6kUXTQ8tNto3DmwPUoW6ZlgbsQpMOIBK451W+V2
vkaRKs/WSR610WPiVstLdjpxdL/ND87uClqi+roMb/iMaiTv6xY7JUNkILylxf+fquuCig6y/jWr
RKZ2yBzHhW0XhsZsaLmIiL1nx9+g2yROjYhFP439yXaxziuWZsfKg4L3ad6EzjAQixLRkSfuXx1H
a2NtfT5N/u+VYsAV1axyMsbug4bfxvolWILeZCTpTL0gZQI61PdJpYdhFWqlnXPZ8N8oG/Hvldd+
jC+GN+83plk1ZlsD7ITIj1y7dQSSCJ3MWbTfhGGdy4UmoC+mdRUHd9WRkXwyewO8YSzGDwiJHEuW
OzjTJp5yQv7+Lz85VkUflnNHmpHTNroRM0fsTQbFLwFzWFmLEzmLAZ6g3cu7gVmWZBMbPgl5qc3b
ObZFpGV6R2cV3RgFSfgw7OkUj98mkMS18fYK5+O7vmdR8g7FZtl5EkErN3iDVBdAJnA1LUsR2jlQ
0CyZ+rsm27x/fcDOXVBHO3mFknQc4skRsA6UqwtwZIKFMWJzkXbhpV1L3OnTKar2t4ZMeQHVA/pu
PHeHZeUFTjZ9Amm+axHrVnV3iV0wSXI8OIRI2ekSOHaIAZw97rEd0F+8aN4Xp+F9fDI6r5nVmM2c
uG0pi/rzZ/Q+3qSAVWPB3aZAbGZtQNLdBE/SH12EN+Xls9od6d0YwyH5YkQ7KyDqwHoi5Tuq6qon
O21mL0McyKcr7adMSbfGlRiAXFpsplaP9FXruym9ipiiv/Ug9kOJU6R7Aa65j1P/FlP3PvFQ38/M
8X6GQ27UcHGZWUG29tww9L8utDwfTuMOnhOfbU4/EQ+bXg0GPZ4wF+WAyKDivzV2B/PX7enWLZb4
ugMyFir7JcSlbNVHchjF7ysstI4UW9foZD7EiZhIHiYBZ3uN809zZhffwwn5cjnFPYE747IFzRDV
cUtCdWtpHkXpT3TVJzsuSXOQU0eGGiZLl85EaQARXrpvxFcMCrIGrJ/aTqccPfSrVUZT0rE6hzjM
H+TdHYC23VnfY3462YjAFlqa+txlctPS/KVqJ1d5TuRTolJkdbnYufp1ZF50D0tVY2z/YtZFZLgK
++FpEjuKdad1yGpkHUODmLDRy3ZroPAxvsN/AxrT28TNbtwijqAS1n2X1pHg93ThobEgrhDFBDgK
FhskWW/Q4M6LvNYrNQTR4+wFxdJLCvRRcXBLv0h8dNGoWmgYYY9KKaPY434f1wes0MqWQou8/1dB
fA84+dD0sRfC9NY1AR1r/beDrPg849n0Df2Ga/kbIhd6ODt6vcvhiEjMfJP4sgx4itXV092xhkXQ
2xarFc4+tKi1fRmbcuxXmgFJupIA/vYfBaN91ssT0QqYmLIsRGwy28wjcS9OlUFSMAkR5E6bPaHx
rsSm7wwLMjrmna4JeOgrI5FfwZgNk1R+uqRQcAPIus39G5+6kR6zViz+S/Olb0eJF1IAQhgKueWC
/0Xd1D5mUFssxdlBLeuJIUZ3aEfc4r/zP5jAZLdK1iPLDsJz44bx5alRA1PSnDkwIk13v3ev8zGH
d37wZShhZuMK3cGyDO2ZXGM60NdyyRF52P188TR/HkXjICLMWaAWqAiP+c1tO2mFIcVKAbZZLw/y
f3opwpG5aCH/DxLcg5ewf0wtEzgWqHDFVn65rG5iFwwweDJ/0YrCtBz3VKblilG6OkyDHGR5TzfJ
FIgYujPErf/s7MhkZ8ZpJvkbqxmp0oCKqo/yoTtha4r/MFlSVJl/j4u4Rg6NsXZDjK1xGyCydgwc
fLTip/Yh0LNqNzyzhLFUE4ArLLN+SXmnl+P2ojnv65xmWoBLAnWnWh7rjqlMaw4JQ/hnoX4b72Cq
HTJKFRFQs65ye8XBpm3t6f1nwet9XdIDWUgEsdN+PCOczDTpUzDjma93UNHV6izQUKgEvq8u1QvJ
oxa5k9CVYI0HBkGuz5+V+55pOKw9qRSwbVcHUTkl7XJ2DNiFRCZQezcFGkF6e+m4On6ZPyAgBP7s
B6mgg/zA2+o9ph+cgMPuRMcsOU77k1LrZSoKjxOv1fjazV3h+aClpmS+VE0Et0RO3eeZVfwvTGCy
nqF9D8v1lITuNcw8qkBgUNSVpltluSRk/U1ZqeNgwqvShhOOXGkGtLqM+TU4Tn2gHOP+NcBTf5Fq
jhMLSaMYn8uCKesNzqSJUYXR5i2LXVDnMKeasw2xXGehzHfgpxz7zSJUuIOxU3QlfL1+kGi6k1QU
wI+ZZKrzVudAmW3wwhBS7tksFtTtUZMrIuIa+Mx8Oz9wEXO8RoF+sGCVJMT9E44rTUihDvuiRHKG
kX0OQPhOpwPfEgjJ0Qrx4+Xu/uPu8ZzdZzUPb/5lNNLvYxFvErvs9O6A+C/5Wd2LVglW+eIApGoV
vUN3X7W1+3rqpFZEBzbKeB32TNfN45VE4j3HNGZEm5fFcfcpaNmKxqjyQ1cf7BcSkuKhoQxQWgLM
FDM9sZRrigom3GZXCiuUpv+dWnENFXH0l1vYH6Vv+K+nPcv2zyPu/ZFIJFIKB8HH4RiETOrnjWrY
kmtdS54UdGjGOsy40BgHyZn6onVhl5bu4wMH3VGw4CqZZOe5hD1ZwBzp6oLEwKB/nyn3jhIVcfij
LuwaLbkGJXS9DZjBK4Al2gbLKGBDkcnZ39JJImfTEUqonfXuAUbiV+vozLUI+KdgruHwo1a5L2/9
c1u6svB4qyKVOX3Fzg5S/lwOh9d8WjpPXd8R3iQIJegPjGf5c0bFS2byoR+9rbfvHTq14ciVoKVN
Zr+yvN+OyIrIynXAx0TsmxIiv8mZQpaZwB3RbUu3Emk3kLowaQ6F+FEY9akn0VRpbQbzPhTeGuyd
nBVRyan4QFzdwqmeaQMFSLIgwHYanLOn5QlIG6X4LCXnSSfp/uGWa6SAWQjnlZvSQBwFNnbJBw1L
cd8IUO+mON22BJu6aWNiCTRu5uX5QwLIQoYcjeUvuWHKmcGtMZmXdryZUKFw5A1f4KUX8Lxs7Yo0
/VS9nqslpZku6IfK+FKC0ix6ZztB16gQLOZQHF14vNKK6CuBGilWvPyiXNbzp5PgkP0ZTwPkTViH
cITk8k/Y2R+Vv3fNYT0JwAiy7/k5gzOfBzfMet6hTrEc/LgW13cOb5w9d9ZX+gH6Yp51GABotcA+
K4tjdBjYmtAMtu0bStux4M6XKalkBCUPa8Llt7M4ZZWs1zAw4A+mb1eMMoebYO6uIb/av7s4osZt
GLKcPMbxWHLodWucbsAVZ1fUDLZxbVr1kJyALvsuLm7vzMoHYBjTmPhdHMCoZYoGBquz/uG0+AUx
u8WMZQfmVPkOR/6Nq16vMUVmWMT5RgfQnHVs66ztnqFE3+K67hjJJZaqaqpdhuRStG65lbjw1rO0
ABHkMq0rhqm5O1jEmwOM9GbOr+XeBCYh7ynX+GERNAIRJ1PP1dycv8N0mDwVnYoqCxJgJcmT7uIT
1jCYmx+8nCU2Hzc3jhqWDMaxQ3sb5DMe2nMeo+jQY4uk48NMp/aUGeCQuaQbBvj28jyG7r060JWe
C4qBD11mN2MdoDzTG/k77yiVUGjsGfqFtgFDR8g+IOYVSJs9fJhLE9YlhyYCKs+2jymffAe1KNKg
a/sS2kHeEJHZOFqisXZlqOEZedP7mNGsAtwBK+ZS78EO8HjHEGl7ARB7JQ4TzE6kzh7V1glhxa+G
5+AK1TPrAn0XpxOdc5tgzrelL+gJJfmEMufKqu0cRR1aEOfzRC2ZzOmvddxHhmUy4G9iFbwy0rmL
3ViSt8Fr55g6y35M3D5hZjCIDG2gOlAl1/tWlbbktCA/0xXRiQRhyJToTa3V0C1WTwPspFJE8kyu
hVBlQMRtJp4Fx83O9GZLQC+AbHCXK5eo1t7Wv+PMx8MTVyFZMLA6gGXV2S4qBTe4cy+r08wrJpui
SrF6vxChQMr715CRXqrjwi+JOuqU09bEPDEIe5Z/zxSSPvUYQe1fUojqt1MUkvrkGF83dbrBGNrG
JsPbGbtaWx7LJngkMFxb7Lk8zBISeaT+SRGS7MIU2dMi9VoJfhNTaaqSZo2vSyAsnevadqffnd6G
TZlWZsL9u7XT4xNhbpNxTAWV7Nj/INt9c36YDJenfwuqhGCteWBZNVrAandb+Oq7OTWumKxtcil3
4fJHVBggAQVwJeXU9aDMjZXo2adA8Fs7XXCmKnd6Afiim+vb0KshdyB+sA6LfbjRqU5Z7k5sckhd
P6cu2KPnoLJUqBvGsw0vCHIdPpfm0EvPTmz3VPSFcuFmkf3EoDyfzQ4lllc9X6OenVayA3VW4D8g
mFuovx0QdLCGjELV4d9C40BAPqN/bBkdwEgqdTiq+FeEOd1A+sNxebXMkFvqBzvD6Hg/9qlvGpyF
ezOl9pKybjaUqF+qBlN46X+dhbufIRAYRPDsApX8Hy/UGBiM+tEKAY5KIB1zM6EkamNuqykjk0kc
W7uvrUI4p/B5cinpqfVgSpeuaJI4tCTN1ExntB7M7xWWRnYBqJrlHTN89tHbdGdJ866yMTgLS0Uj
QoZyevGswTFmDYMawJMyZcaCw+Yjp9+3V3o2PLit2JBxZXa+3nV1f0FNz7yyhrfVbDkAHtyAGI4G
E8xvxAhlTd8qmYzhj2VVZjOaLl5vIwGxDDte3ryBwUqc3Zb/EMeELyiMVcMc0Y8O4HDMAkIYe+GK
nNOBa+xD6rSrDCRjcq64mVE8lHJcvMngCRqOnnmnI9mGjAvPTLkXmindKqjy0O92X0CErK+xzFxG
VG85g/BxiFcfQ+Xuv3C2V3SRal9dQo+YpCLg9qp0a+VjJYynM4OWNr7i/v0CL5CGrRBCnbfXhX3e
gd28a8IXFYP1INhnVJX652UE8jNiePHGXTSeobPRUe5YEMrnrUPAbVZvSS3dHqI/CEDDUsBXWnBB
qnKkKfSDviYHeanz1W9PTADr0pJhTlP4KWK7xuXo3eyo2tIaYNb1Ras3xnuIjcsOLy/hqhwV7rMa
ZVkqb8nQNQ/dq9+0y7slMAfVjEUXYD47EbvP4tSXTKTB8fYIcaS8FZVRVvS7xEKG/Fd0NXj4bgHS
7W+08PuJo6e7qmnxaI4Cf6uyhQ+iPuZnywmvabJPRuD7E4QNLVBKbO1vxzznP2euWdqI3/FAef28
8T38XFnKNdDbs5BPU3KkLPk8mnu47gorV6SsYyQnCD8Cqgc0hAltdsRulN3AG2wCa8C4oPtDQPex
oSc0feJWsx9+Dlwkoj/KR3TzliMkRGG2Yf6x9ARKtSG9RGAJmpoEZu8t5DsOUAw5mSekpCWTS3qG
+hM4e7hoZQ16FJYgyjx8TUx3NDoh934jJxjmy0UTaCYGGSpXSZLPGo11UzjUN+hfIE1HjHvSH3x1
00j/ZdphTRcTYZHCMdg4LTpndfI2b4tvThT/XUPlALuAz8rBKpdw1nW1xUS8SClefGAdCul+TO7m
QTbS0nfQFgBxQR/mxPfjavbJH8yP3ZCbsPsJgw/Y0JGlqsA/QObS7rKEmPj4dLBmpI1P27mqKvLv
2BEOBZY+STQjxDlPvuFl70dv2SWR7xnCiUpvy6j5cbdn+GVfC5hR6kB97ikrdyrbfJY9H1Q5nODb
00+ZCwxVN/Hwim5qK1e5QWlw4qjmQFvpvEV+jwYMlG3lo5lyPRQzB5R7hqVoAg2eZYIVs7qJ6jv0
KqNczfhAzXcgm1KUB4AP+FMEBD0BjRKc0mc0P8j3gWKAWwfXShMm7IAdziKJ4mPWT1fIdz6fOPX0
CBv67pmdlfGzc/YUDtv+SEbebhUWmkZCXNXNT0/jN/4hbJzC++poyF2x9sXc4FAUVrz+A8sZwSNj
6uRKdxsrDrZiH+8IHdNsR5JqnAeqSRtriQnf4GDJ8TgmmvIlpiL+Ln/++bRKjFl8BVXSAgB2pFdv
F4rG4baS0gyrEw8ok9VJUzEE3uPU8JV7S491sAmPHqJE0GG4fkrVvqIOJ5iknBVZSKroQRqqSNBV
YTXAVsBPyIittN4xUbaZuqi5nPynzA+pdQjHqmsJjovz/GNR+K/Z5POs6LbpyeHugFWaGojOEN2E
d2V3newla5hprLFDmMatzfThuj7N29qdtnX0F1Kbmro/Chf1fdJGTkZWdBuZVUyhwecBU1N8IIRg
me6sP/P69qAh6hnQauaHWgYEsBiilNxjwz7VWZcK/FgDHcVQzqJkfvAycjKNlOhNrFKSiwqstbmi
KCdWtqW+mXbF+lLpXqQJlFXoJrkL7P0EY+4g381mJmiFQpE+3rs7k3fhXX3HKGzdl/gvjYua5X1u
BwEiDAXYsjDm8N1MwmpyahSGUqTyTL5Ya7pJyZPd8yZN/T0HSFhsZdWIKVI/Eh7CVSb5zlE/v07S
nZyX4arnek+NxPCVVBiaVibbZ63j5r1rdMjOFF2Wv1D/4wM0iKivmPmW1/Hx3M5rdQrdNQ9Ygkif
9K8ds85S6DbHFDKAtclCXqdPBbItELMdUuJueWSlLX77Y2QLlKM2DWviKOtTQtrXXFMuYTI/kPVI
3lSpoPVQc4quCGDz1vhoDgQBtqpsknaNPae9h8Ngj33k3PdwWWpoauQfCNOGZqRRaoqRkaKyA6u/
K7d/tGUuyRqzClHKQOXNYQVs1sEfOqjBWoDTfiWM9TrASPVj0sFi4v6q3sTLq01mMyTlLD+UU67G
+GHmnyOePy2K0ALonS4UVhMi+rg8osLJA9aizjYyuzacirIcyjl4nhG04DKRYvtH3+7xeI4ll7j5
sTvlwZbxZHkp95D9wwiBOu3vwYI1qlpm0M0g1AYJsFkq37PTjqPM8exC/iLdNKoHgmD5rTumu5t8
dFEYDDXulCzu4atMinWGe8F9vv1MwTNZ8EaZDvg7G7tPBT2klWTG/BjHk37Ib4GFzr+WjpOqV6TN
CH/IkG716hz4Q+71Ur4KgqDVzoh22U82mAHriZWwWX4udLRaj3yULQ+Pr6ohTdZs3C11vufPc+QG
7iFpSfvrCXIQO9yMDhQMf9q5PQvl4ABlAGvDsXeu5sBMwfNiaUiNi7QQNOHfXskbujx6PmR6BWTv
wFT9buOjAtrU2W15LCyy9SFvtKRJeZUhmGr4vabSD85hylnLRZCkiJafR16JsPIa2uznXMV7lbze
nhNgnW/Joa7etIETZdlaLfAHUzb/bjG0fD+EaW/eQSCeAin0pV4jC1aUyviE0+uO4BahP2PR+U38
S5F8YdtJ+wVXB22z2wMmWt4fMdW2YX3/q7GvmAkBCqhT2QoI9072RBBBPBqLJSbCMJvmw2s93UjL
NlP7Fh8Q8ZhO9HvG883lNHGnoIBkGUBEyc2+NM5PU0CLrFRU14MrbLQ1fgjYOTPG+Vey157SJPJH
wjnUKBKawlHtxjsHeukku58f0sa2u7nWd9Vs+tao2iOcouJwqQe5vHnqzV47EYIFNxYdHOuC14ao
N+Y0JOL8URMAz21QjUSdQ7dfL+KYBkp1p0ccstaSS/1uRnIYivsXDkTOwMjgSVZXgTuhdTzq63Zg
+Yl6wkmll4gu+YxQhZ5rUw0bDhhQwg3nRi7ZBfrmlvsKKwNbB89d8lT8DnFxiAtLeK5wAY4WpKjb
FlQST9YNig0lPIVWTyi8aIcA2tdxxvziZSas9A/Q3tuFyo35+5ATJc2q3RbdTtM96pWeXY4NBKQq
UIyel9e8oeZcLR1mwuoWDnRf+zH4ZBHyMi/1XaBQQ56me+6hnql45o2BBhKQWeW+9kpUlGWy8ieD
penB82KZXrqtu8hNS3OIbFqvjDMAfmHY6fX951hA7GnPl7NdNIJ35tiweHs3AcpzU0krZhs7ofS3
D5ZQjLF4d0pMeEj+wFZsnBE3V3EO3fRT+T20L8sSQDXeqJ53RYjXPs+ZqnYfjzcaZu/atky59wpa
dg9dZkbtmB5G1GiCmCjLL8aZaftRGpT4Xogy/1HTTsDmpKWdlB1BnA1ZGNxtrdhCKiU7MK+vj239
haSSFSklAtvINUzcZqBOB2DMe3wFycG/Sapt1xpiqTkUnUKz7QkdKht16vUQsaEdW6i54RMEoiIU
JKaQss4Z68AE2SRu3tWndq3WlcIjxdH/sQyrr8Big6zcGRTHeupZI11Od4woUM/7t4OKixxVv7O0
hY7ym5nb2qanz5LCEImq+VMUQj1PfkAhu6dIO3p3ip8ml3X7xijQqGwKSyfRepgEI2CpXA+/xtx9
apZRCyX0DhYVrzvL7KkE0MjsXfKbN/evPYFMuo5tq2dtR2EOxfUVeqeBF5oa+EKzNtMUpbWC4hgf
s6Hb4JRufLh7nL+WO+qX8yQPgDV+K9o8FXL2ZLhNm8gi9OjPyi+2K24yIA5dpOqevSiSHghGkLB3
DQPWsd8ANYU3PbXo/PZa1icUlBI2ZtXR+LiujlYAYOlvyNoeDcTSZSIBdzTEYM9kDpER/ZcCrLku
7rqmIJpFBtAqDoPjfvvGc2OUJjhA8Bhk7/KPGG1MCAZLBqY2PYPHVj32AQW4nMNJY9v9nqBCszJ8
C54H7DqAH24+0UBi1kcnoCMhWkz1jz4ge1PgkfS3Ww/L0cLaQRTgoG5Tj/ZdYc9+4j/nGEYBXORg
JrhrHzwbtFeXMcyfQuCfqrKWdvnLVZU+HLpCIeayxwupI0lSNGUzZfWFzk+Ok66w3Y52BRtExfr6
pzahuT/DaaVqmj9i+lJhfC0dhZyutLjtnThJ3Xaw8dEWLWzk/DFPv+vmEXOjN6gWtBE0SmhBzNB+
Q2Ged1Y7PoQSYcqJptwanDY+nNxVx5upb/HSsLEtmsniuTo0m5OtcUFsSUqzOUMKcUL8N1eLAr4j
/Bc/0hXa3ppGtZd+RCE2pixJzq3FRLRXzZfl2McZckh7MH1mbG1UE2jqMqfqW+VqOKmHHMD0iX4e
r/r+r/3mg0LHCSNeO0WF2jvwFCz3OT2UJ9RMy3gCiyAgUD9LrGrsrihEZkdG3BsY47plmMldWNZj
1eg0CuEdy1xxrLwHr+MtIP2mYlYB4sIXNVDsbUQJV05xF8+tsAx4BsPPdDPhpZ3A9Q/8tbDpCGaR
av2pvPWx0GDxk9VaQYYnWNS13osWO5XhBImPaD+Rq+GUvnQjk6iZQBMLEj5KzBCYewslW4iQ86vs
+fNnEzTMGTQSQt6nhzeQ4GKGXXnIrfKGXQlb/XWAOFB4oM2SvCxWIh69fTZo89/bO6Ky2wLtsayQ
m+0Rd7TWjnVHzSzbjG8X8qYmK+TjJAniZpaUG85No0rw4hjWpgPkNpk/r5n3l07o8JnoFnRIGRUw
BIGB+6k4rVxv5UQ8pZqfpGJSQKHow+WTBY4s/xq7V6t0vzmbERppX6YFtc/IkNcYOrm5PMM5gpLr
tM4D5rny8+7CKfFtYyImaWuYfa2L9F13s3nPZ/uIr3wpfxuONh/g6X6hjXMpE0sSWzLLasgv9Z4O
qlmG4TfmZLyJG8en2AJ68+C14F1EA0TshgHTOMdkmvOVSor5GaKgPWxT+AzYL8s6maupmp63E+eF
7zlI3eJwQoc1w47EOK4xkGHX83oVLw71TQGFY/ff8rElrKIpiz/3bmkZjN5HGbRG+jyl/TVx9wJq
1FW/SOk7xIQCAaLhCIDef9pnax9ZBQI975FCELHX5BAgC3cQiDUVHKwp3C4Vj1iXuVpCLLqaDikO
376gUlBTYgl0HrWj8OmRFQs4p2dXW8+QTpuHBvoas0Wr/Wo5GbV8su0Mma1m0sQnQW7/PL38pzY3
9OedM+n0woUb0QTTP9///Cv2FJPrpd3LUCc+0Vj8LbiJ0QoQaIkR+YIEapCtK8NHzXZ12qKxhy4P
8VxUPS8JEkHfI1LA8pO/eb2uZSrdxnndF6DJlVP1AFOZHYkNuQ/8zt7qtGrmfKC8lREhoyb77N2m
pqoZXgVYrLgSLwk8A92IMFFgx4J8evfq4xjd+GUh9XftGU0J0vBYavorjr9S9brlWsTunIxb0D5i
1gISDL1D8FQAlAY+GC7XVLycIFQzEAp69tsxFvhg0QBWWICGp6gG5Bc0KFN5Ja14qnl2XK0P9d1a
ZJoX1MfOtk8EZ+tasVTnccFiWwrAxOo/2BgxOxiSjQG2i9Z61pNyVeQxhCtHtwaXWfu6yfZI+pI3
1e++E0mq9xn6mi72hs47L1LOYD7QpqmHSTdp2hk+B2JV71i4GK0j53jyKh2GLRygRuoLXGHdMg1F
8uflXwfJdYNkS335sUXxeW+S26XUPiPX82gktTx51qK41KXDAHCiy9/e3GfcJibI8QMMjXUC0Llb
mwT1A7xTCHMgWCe5jzbauT1+8wQRFbgr6UHbD+hVrvNe2KmbFIQcOGg0YzEfGul7jsP8fRaQ79cC
cuM0ZxfkPxW7n+h7QailDoKUJGzIavoZZ+KpnH160UMBiaWbexvq7s5g1MZ/tw7jo6LLXBDvpcn4
+o35J20gna2ouQtt76NWCNKsZF8S/giVYOHjMP7FbFOw5FW3f82ZjPG4e6odrHab2hwbs5ERC0Dc
ycCzF41h3chV9R0NLx2rTKsF2rPROO1vxt2rqulHnWs+EH2xSGgx6ZR6CsdvRglKRnhtGiA11ocV
Yq0uH0ni8Xuk6C9MNUt+lC/WKubwplnhXVd0VkxG2RbjTDKQbMgl1ro7Qx6sQp3/NBxfMojT6pZC
9+3lnMDVJP5fNz3YVLhW0h/7W0y64mA9t3wjGlmZ+jpfE6G942FJVw7ui+0Bij2wAxnU2mCUlFGY
Io8YBTfyGHqpoC0slw+ZS+E0RrfTkACTs4WrSWjMJp1EEVAjpBbL/p/5+yKvc1zK8gLW9mIJN5wS
soJXpeGkR00gAmdnrf3a8fdoBotec2Id4f8EJoUeZ4OA/VADNBm6RNdHvJrshMlXDD8AfkRQgQZ5
AcBnbC0uYFOaoGMznaekqCfVqUupNA+DSG6PSwEt3t0CchFlZQ+Ek8HiSLhyl87Rg30ZIF8cb7n8
RuHL9xIe6JAJKM09XuhcYA6sh/jYnTf9csD8pUG/DFkTUGkVyHZoF4ptdZzAr+yBgUcT9v54/cC8
didl54xinG0uohoNP1mqJjozpD96L8jjF0jVk4AUsOTR1Y600wqldy9PdQoCzKDscLTxHIzWa6od
R6j9qRMhBo8riJ6xE3HjE2HFVHGLWWwMTpJxAPF/eOTQZf0k4JJk2l2cBWknwgHwGYmd4+T/XQTq
ehTfFKq4tIq/fplYFVSvRP/YQssq0mxqhbY8o/GtgGNPxP610B7E961ZGQzQ+4d0zzpHJ+t97IoM
8E/RtX2v1SRbZ2K0cCgOy62wiLeIXNf+d5lmoOX2OwSN0/8uocWl+bTsqmS3Q2xEzgscb04/nQPf
2xFPVuFQfBPkwfr8nTyZBNjzcYXZYeQ4TTwy/4ICZX5F8rgd/FX4OUGge6W43ESXQMg5mWCrTFBL
t3AYsDLthC+wUFmZxyrOXkNBX0z2NUVb5zSXTBcGak/PTM6LeAQlTp2qq5RpWKBIjsYOonD8IbdJ
h2z19mdGkPVtCzO9JC7dPf9mKUmX121KZ4tssUBTCkFRzMSJNO0o3C/5ukdvSHgWUa32gTbCnql7
TCyZCYfmu1NVYpQViCnSW8W+G2xl7Cdrq5EtXp5shidnhvgUVO1S30gQa5nt5VcTnunPd4JDNhk8
IriAIa3H8iB/ar8QWdLZtZocD710RQonrwb5C7e+hgEVfZDngwU8zp1vngXM64hAwDm2KbJ3kl4P
K17x68vzufF+5EpU4CsKZEvfqJV/jjC/JucO79oYeMoIRinWxfWXUTy+jorDcq+7S0SroEU+C5Zr
oe1COIH1BX/DwFKQ1EAcSToTT9YLBJVTu5WQGMQkUZESKBTv1WnJ3qVsuhnxN29yxgxhnuozsHAQ
NHkvB4koGMB+3DrPbp+wDELnUrq5bm7AFfZ12ez05Dr5Y7a0CiG1ueKy6TdlvCqEgZzppVImu81t
zjsOHsrxlt094yXM8phYsUAHtaq+26M+LuqFn2zGbH8COg6a+obIkeJAqk9hO9jB2ZAumX1nRSww
ia1Ut3wG1kxsPFITXmQYO4OlVwHmB9zIEEsKmoODvIF41BHIztQxRe8ErwZblMg1a6/94M1K0EdR
P7JwIr3FwVbbIn2w+uD0YKKTseJnefn+JwjqFJ9yEn+1d3IQsk+0dzC9P9XtSJrKekxUJrr+cz+W
U+UNY+Is8x4Ts1Ir24838Q033WKJZ8/gJh92FuY1hU3r6hF2udrUcvlxdT7ufhMgzW00iRxOs6tb
eqqU6SQn9+TVybo7oz6IKzIW36DXfTnRtlP6VS8Gn+vGoYFEb4Q1UCZ2tgxU0qFg/auF959sD0Ze
kGfM/eCZYIJYlnnZVdNaQwlO0Kb+PWM8Qr5aPRqAPJJtxlX+Ra72dkmqD/kVqMksm1q8SZABpSyl
qov48/nIZhW2VZBI72ISqPon6HjaAHQ2739JkGr/tq5c+nBQY6dA1GQe5eiGNfDVqV6Yn6Od605c
kwonQxlS5VvlkQ86+vx6zRhtZutuPP9WY3fpSpZ0jtYFubeEqBHfYX5mEelNOcy9YHD3k4N3spjb
9CldPglfohc6ZAfNqlxvTdmDu/kaC17rxAnJcPnIDE9SnKfck8XjRocW3aRGUf2tzdh8tqdiXv66
5Hyixi8s6VPbqclUt1Nd2xcOaqrdrmQ7iUKro6rvY66AEU9EYVcM23mCQ4Q7M4qn2D58GcTBEAaW
HkXHrih4DP9YUnA62V9mfyFwImGdaHBzSpv35m843700w1B2Biwl8azsL56wa/84W1Bhedx4MZTr
w1z/xR8jpGdKBEzggGeBhzihssETLPpAwbskg9Vw2VyykvX8fIjcHdEKg2jrs4YAmzKpTCauVdz/
XnHTHeF0Chojxym3o9XGcNvGATyHYQUpELdY/ImK3wbrqpv7Dasuwbb/aj2V1lh4RryuwNiWPrtc
iczuLs35ko/9IUZ+OiWp2DmPyiIjurNagRv6EaN9GWyTKHSBBkM9i1MPEuCBsJNFKqZAiqBh4Eic
iLDjz//0c9aaV8WqnZRFKBMhE4efB0bA8IPUrHHF2oHIdqx+sR2EIS4Y1XJsV9qCJcVc75cMsayQ
GrXWUeCozFGNShuYs2P8z0em1fhbi9KnTkSkeZUT/cPRvju8eGJk31m4s6ZJXJzAsjChvfAye+1a
Eta7h3KTMAT0veWMPeKPIQVLSqf4clcX/uzzOOaLjXScUiMHp27imtx82uDAjB+TihcRMwegHjyx
whbNUIy6GBkUE70xUhrCNCrZobNDzIj55j8N8w35AfbtQ3GtVrBlvff//KjVMZSMDGzU1l7f/GTN
/Qx8uH3KdP1vxduP+0DUGQmnnV9G4WXrzRutpaWY191SHkE72ARX4o6QC3c+JK4sk4ouj8M15A/v
kJzQWhIFUaCqD+OnOYdTBPrSejn+KAScJIyBaxkvp+vy9GPakqB5pkd3h+IOTL+2G5RmoSVC19/V
6M9uYKrlB3SUilzOTOSCp3DgtB3iYp8hhhd8vA4x1xhu2FZcnJFUYzOS6DkJR7ZptEyG5/3nhTXg
ugbWQR8iCc4JKsDTXWomZjIftimdePsztrDqi8Cb33KDJbMxarTZpAEobuMOjt8LQ+jxK8SNXDmq
PQbRCfbHZCvYaJAwJmfmj9rm3btbaoC91qc6zY9hkhsNw/wO5rL9ZksWnVbsYzsoQJmBndEUUZVA
+vCXFthYyXFyazbMN2oJk/RTCyO4DmSHBwHteSV9e9s045N9YdTRdz8c7wQMLyuBrYooHyOVTf6U
C7QsUqrrlNb8RAssJgA6gBkDc0Anvg6gC/PTWo+LBeqFNRr52oyGpdh/XvvtM93n+qUqdpF9nU7X
lqirky2UPE3cP/Y4vgAmupzFHLyxXqqLtJWvd3b6ZaYS0zz+6h8TeRzvofubvuiTRTSyorMffic2
Bby4vtR1X61yDWT0VC0ayt0oHgJb6oZTM6LooZPwDI1QjfjxS2MXafCGG10ynlhG3WREqWzSiVxH
suMsiNXamgRFWxHiD886dsFFkMhkzlh7xbix6zNrqGjByLDcuj9F3Y2Em3YsGhAXR+rC9rEXCIEU
RzCa56vKPMvTW91totjhhli4qojVRr7u/uVdRVeObLKHaM48J8r1tAaY4FWX16IeWcSMyl4NWqGB
XsHbkdOF1slppypglvpdqq4+EmV+pY15h1p44ZrvKnUH/ikrnVWVnDN6dEmvNtbhDfzvJMBczxXH
DYL2erJheAyJlMKYzGcrcXPOH4G7TxRIPiMUW8jjGG93YRUKKEOpkLABLBCwmbBuWlrRx2dcpjLU
r6ZFNI62b7/kjMFRk9QEn3dzWETqfNOnVuJexOWgdauaQDz8pF1BMVv5AqwKarnbXwyCJXUd3kPb
wJrPpsP2ZrFQ1HJAb4KzvXv+K7qgfptZiw4/5tx2Yq1lPYlRigrtLSNwwmmg/rIVjWNxZWbWU4C/
XUxfs0SDaKuCaREcPZo3s0xied5ZGl//wmO1bBX2RkKRy9TcsJChEkUOcRkC7uWnuKBxdqP3Ul8f
cOLSgxPW6qnBShw9Ft/irFzumIRwtQDcugLw7b8xXclLGLeRVYmoCGdc9EpbtNSAqdosLFXFOwW1
igRgajaKDQw/T+Ou0EbVEi8rxWW8D9k1JO9GVhIlY8QPsXtSTUPgLL9nxECcHWSGnRAUXVLCa5dy
rAX+myvh5CKT4Vc32wk1PX5WDu/Va99d2FzXpwCNaLKY53lPcrQy7RYUzG4ChWL2+Xn/v76weXC0
tbW2yJM76bgBHnIKHdVtfK8MK0JrRVCkaVJe09p8j5k3Q48Ph4awf98C5QajOFfCCY84K9SOvHml
O+pKUxN5XNwnJhjDM0pJCND3U/G4/YAOEzkZtzIF6oesDcMboCtr3h7DXVKs1wAUDs9DzxVhpEkV
oDzpu63I1QqfecRQBKofmg1JsYsomXZ0fu7n7unMpudrMth/SvfpUe+e6bO1OZorTtsEE0q2uCAu
fa5fQdbWEU3NRSxSPq1dCYskEe3u3ZRvWw4CVhu3NvAj19YWu6buPf+07C/eH523hm5vpm/L8PN5
K4BuywNsebDtzKd46vnwVezGlRslds0AvtsGYgjpEgeFLE/yOmPJTvLbjBMAarNVAM0lEosxqSMs
tarIV9HQEGGxVOGJGHTG0Vu/YE3my1t7TU+fG/NVJ5owDQnO84OcPXjgeu1Yly1iNSGZKMZSXXQS
keFvYdlXuFeeYkJ4bGVUauqmKmLMbwn0VyXLOHa1ZYJ4z423LHHkZd3tuyjBnuc4YzK1/GO1h7VK
ylf0N5+XY+y8nHosfZB/POACZ5uN8sR1ROA0E9877FjdcJLlIlneEfue6pWfmUfAlYQ8Ip4nybEC
gNO6jfACpiSBgBu2mmcoIf8Z5Ebq6k7tDjnQBmvVlTO3DRnp0lj6pPSNHuuE2sRgEZsLjDj/5P4S
RbSPy4IM/Nzbq6Bkxd6GWi5TlquqyG/HQGCUKWpzuc9VS1Oim0VU989L+wt7QbUV8xTAp1eF22UE
jSVqACBkliyzazPebkBi5B4JWIt+SR5IcHZchbqQHuclSwA53neZagiOkHFgbsx+2UEfa5B3jZgo
xtCKq6nDB5DT4X/d+NCHi2+WHjN99QbgRKFL3iPP1MR8qMlgAy1qEDTAc0qtTIQ14FES83GdlcTx
JNVBgjvc0hIYDaMTob09DbBUfCEqTBYes/shUlMxqffLdo6Ubp6FI0WbDYW/lABnoAqqJkEGuEy+
PHat+GwScI75pv+QV+MAQ9eVEJRP3NxGuYgZ58EjqAxF5TM7JvuatVt47INoE9IZpYDzfdC5x6mL
faF+T9juLKM8mcOvZ6OC0NYAl00IuErVSaKrb+WvF6Njs2Ilzk/AVo6SK4gIDY0n/odo8qErVn6m
g0Jk7mCyGh3Sjv0IspxGpvjgy2grdffZ3KC3Ten7ZY2SgYafsJlA8jaN6IblSfdLX7ZTkn0hKtcR
bop3nnB0HVcGI1/K/mO87VBa2Ei+GfK5xgaRZ3wJVClVi3bieCuR7grnPVluJwyZyKGHubpMkQ5a
gNEN82kWcZ2fGgiOdp1j/TTJwcaacZGVGMGO+MfG3YNgFoGYMcTvyZ5HNuF2KdwHGQ3oalEa9XVZ
SuCiRDa51H2xCdgorqGkyR5y3sPJOopwkelCbH34aSodNoQ7+kRmLJWCX0oYbulSZhJzspKVaQnn
gzCeOYo+xFOZ6Acw2KgojqbVlxuiEs+otpx9oNBurIXPRZxla5LCN79VCx1vrqNNGgAqPSBEX7gc
XDy+5fhzwzcDqpQ5dI3FjptSruiqXNLg1nJ5oCiBLpLaPiLghFklz9FRtBiNBdPozpX91D3TDthc
0jY6qZmdPlM9lNlg09Sdb5nZUaZkZapHoeLJafL/mBgIGWt0XPxxpFem6Nj5GP53uj9vHkQo7d4O
b5KXXbs6VNPkgr+qhjf2P3nvGi+hNfaTBGRwDdkTs1vLMvl4d0uXGqUv8S20wAU086YW/bWHbq67
veCKq7ASiZNwSfhGEjIRimNEpXS4P/8SOeOXltXJFiFgR5ZijjCaoxM98GjS7MvMRD46bYRqtuS4
X19G0EBQNfTPFu9O2UdNlGbQzO5Er4vZMjfpywTbvbsNUujaCtIqT3yvX7n4+4NiqlFBvnZXPNt5
DNpB5D5t2nW4KzE7gE4SXbBdFBF94tA+sAVYt658kGsHsFgfWsNUnZyLvdor4krBFgdnNxqAFf3H
fEckIuO0Oj0HaP4+vZTAyLOzguYOjAUCjHiU3L885axacDC6BaN5B+CQ9W8oUvmTb+fAy+SK94MZ
e0aqPBdhH9ezIdS4tZyq/C8uSrCneussQNVg+5NEKLEGXEafmQp6qE9wij8tf1RZuC8U5Ek3v6yS
+lSFGoofySl3dCpOfrYAg/SY3GA1lX9pBaMtE9S+1vSDTMYwDqYvXHiqMv9RwessIl7ExhY6P2RX
Cc8XnTz15LLTy0DlVQbAPMRCvhFgYzuSV/dw6vAxPZ+u26tnCQCTTa0t84hlcDyKCwarznpbXbgJ
7+Ltz6cDvyBc3I8g14ZhHZfc5KeuxsKC7QxNU109EPIa2vlxG1AQUU5xKfX6Vq85qXCP9B5tuYxX
IWD09J1bHeC3TOKKTPGf43zIIWkOyh/HdsaToJ644rGNjfoSxZdpsx40EGc6kcNd81X+AfbufuGG
zGWrPu1ltN5mKuvuHytxcGMcjkaC07RVuoxJMNUGFQ3ZTyg7wCE9yLklMEPvDEqLH/XcYyo1z/Ts
zVl3hx9R/mPB+QlsYG0jDCpyN4cpgpBUEXbXseuzMjJwrq9vJMNmPIDmIxbxHKlyGSg7KnmpUSEc
z1uGcxkZ2hA6x7LRTJELVLIJlEmY1K+k16NSZ0gg9huDB2FZWCC4jDappWiFf6LL7OCuQ9O2Fr0m
OY3eT346lSMoBlnNk2qMD/iiUzS65l2uZX8b5axyGO2WiW2g8J0NKZYnSWQBqQg5WCMhdtsbLKuD
JDrkejzZVJjFPSMalw+qjb/fh6kcMdRChAn1Vpk4ezXPbWLiKQ2bTibxYDNlvWD/Xp+OR4uQYi1A
tZzQXlpANKkdd2WGXpbFEJpd1wTarK+BeNAzerZvgAzni+skaDISkxZfe6ZmS4uwxFJB3nOdYx7g
Hw/tNdm7xDQHtmCQCkDdQA0w73KSgzEW1TtX6ifZEPaI2TUxzWjYXrtRmziN5X+7E8n9yVlOortV
GmbabvdcT0ZO1VE8vZrLFIlQ8x+OlfzioRYcRXySpUn1Ls9eHF8w7KFD83ILupjl2rVLuHvrsbVD
9R6qMFr76qvVBVpxeBT7ueZ9dfu8IhsoG0fSMZQgEtxn62fdEg5Gw0anVvSQ20JBpXpiPNIEPtrA
e4v8Ttc+f9m1AJkZ/166Gm7K6keUQxXoYc/tccsYIXMz2/Lu2WLev2ceDtYc9gBttOWNmdcg+/qh
D3XuKnUt/A/I9dEw472Uw7cD/PiaERxAM9eGf/gKEzX0cwWOOCFNayqf0Z5KwQPC4hBzM4Z0xCYp
pA1IowrAKEB/WQqdeBxnZXz3hiuGmBbwjeiAx2u/uot9pDZGhW4DfR1Bj4ZyMFQ3mRMysOmPPwN3
zLj9WFWqUNfbtCGiAyaI+ZuhpPFjo0JFlTuYZp6eLF6ElHV3hQgzb/MM6vKWOScoTStKAdOGWfIL
wWW7lPfr6LXTiy5WLQJ6TnziGRF4FEFOAXQeiOJeZadDauJS0VhhevlVCr8UJXN4jgVjbhgl+bT2
8IPX/v6MK+d8uKFJ9ML1YP6iHKxPK4pFnTeKbKHruwjFU/5cJ6f5vI0e0pj7e3WcKzYRDNIdd2+M
m+C+RxfgDxyAbJ2a0Le1KsRWxK5SAfOXGDz6E3r+jlXnGig0SOleNcLnywxwI+4r9Xhx5vZVpb/9
3mvyuovUXTDLTn5QYrtlfSTSWpycG/voUxRfT7HLzM2uS19KbJRGRyqcHCr53CwPBangkGHCnK7/
+5Fudi1toIZXS4PVQdSGvVzsOgce9imDRp5cfLOn5D7T5aXHXgQIDrS4zKrB09inKW+X5ZAKAB0G
DeoV3ioUjwpkoFyCyB20oQfFSSodRrBujfoS6nY54y/OeowHBEJSxNjE9Lp6EaTRXjMmGdbwnyD8
t7Zwz8vJGoPKsILnlNJgRpOh54kim7n7d+Atv5zqQDW0d5ndCksUA05s96dTGXx+hlZsqUxObL/D
ztQdnLnW8FJ78QBH+bI2nEw3S8xqrzf5uc2dBOjWS7OcHnuc5d0vT2s4ymscXtp+9n0GAROJN6w/
o6n0tNN6p15DGBXOf73Mzqs16dTfoutaP2GygXVAM4sakTWBovGuuJbJNQPdyJ+35pil27RyICCY
5hguASD7MIJGhrbK+FB7wLuQchuDwtmkuPZxHbU5k54MkfOmx3scx8L5Z2L1itvplCL4v/8hknc0
XknkFrtRzDFIrocLGQbyvaEIOaiY4K8Hn2GcTwrtFvAtHIPEiNea844IkCyZUZRJFEq2WwVkjWwJ
kVDLuXvkzf7uQnAFZxJpZ5Yc8P0XrUyptfZchxUd3LNEjeF7vK4iq3qcHWrFdhLjhF+2SZtujDVc
Z2TSVGydEJ/owCYSTup7qKyuqLB7OUdW1+Z5KsG9ooarM6X1swzJ9ez9fF/yzYjrN6Z6q8tJTMnN
RnU1C3WFzmz4H5RX7CdjlzIj4W3cfdo4VEFciEw3nE+KFOHCNZ2rmiud9posiq0a7LhdZoPCSw0Y
22oUQWbjksouQU9sZMySl/CsuIgP/SJMSkXZy8h+5FPeZF9OxvmWz3hPfkD/v6xX+/fozwQ2XFiD
vGrq0m0o/uYiEBtsbf9ZwHGRBv7pEr203L6VdKgMATAGa5Yv5BLYiy7TnYvRQqsBcnHmJlQulpyN
5InSSXMH69QgTVyRflOBAZXJmpHoAHZrZH1IAG465XjcpKutESrsAZeSN3LQOtbbu4P8cMkr03QC
Wxn2QqjJCoJbN9n0wqkhMsFiqEsQyR63cGH4u0dFq+q1nD4o6vzcNkh4Ee3VgJweXfIKG4hOW/LD
n3vh0RHqVZECSo5NuNPetT3iu9ZcfSZcw2RGk0mj3UZlBcEp8mZnrSAC8yps/C/M9Uozi+D7C0FC
UWe5LzX+Gkq3iogSynWMUkrgSPr4dJhWaH6Sal8r3Aig4jJp2pkytMjwKMDJIhYImBA12EL92nBM
cXjFgs08FUSv6f9AVRBwqQw/9ZjYS4Hs4ngL4JzmfIY4SeMp322IH7pAh9UIn+fZTdWTGSoGCCMJ
ROWCFIWZ9MLQ/31o4J75+HV0a2+m70YOmUUqb3dix1HxJ31CnTYiibxONcZeJPJFPlOnlYBBc1UM
QjqOs/aK9taWwTgbFk46k9K+fsaLBSeTmwb6lP38XqGCV5w0jXPjY0dKmYekIpSqLOZrbW3n0aB8
kE9jZGadO+/AIJGQk7Bz00Vjy/MubvXxju7P1szyuU+rEYCkghgknLOEN2ghc+nZ1suDrV38mlCL
y67w8d+xWOQt9Hh7bwHRXH7agrtuxlktLXPBH3D4XHbV3PpRV+8djlzOQR3oMHmQOJHGy+RoE6G2
fnFg4zXbbvQGACtAvpRHULFY4xhL6fpBU1NXEN8acHpduxhFUsi2p3nEIBWSbp89L7Wh1njVSfYX
eEA0zzayqhNxlvnjmFylqetJd8zsSM7kgbSn+heF22h7cNBHPo+OsLPVwNEPSdxcX5BZNWvpRTR3
5JrIf6aUDy1mtO7UZV24Bt7x3cA7FOszXyw/K8hOHpK9ux2z1sKd9o2n4ajTZqfII/P1Y1n3FmLP
vQcmSlag343zqKo+qfxvu4is3tcqtfxuHl2pqPpP4538kfwC4CvDSxllzxrn4aPMn9PLivV2J+1e
E1YVmL+wk4gO3F1BO+j3XtgmLBghoCyYQm29l5K+3DSHKBQJPszQOh5lnuL+SGYrIM1Nqt8t4OuU
uf2tbr27iiRDZ9AmSESuaBt5hg91kBo9sjD90jGR/9EAor7zH2HBHjFQtxvqg5LXn3MMeBR7wf4h
vI9XyzgU8on1FyQwrjYggKwCB1k+TWpTtzg/sYxWCFV7ffNAXZ13UlgkPVhXsS2r+C+U0mJj4fNN
0N9ACuDYmCwwd8SmFQJt6LfwUQ0aLLOOiVuKN/VIakoH8JJEFuHnDd3/l2JMm/S7EQmedAV0cPb0
+Wu2hNk+15XJxG0Svbo0KGl32fgWPVyjP+qlRdGitgyFITXd1Xl64UulyVWH87lzYZXTrZSC+sSN
X61t3+bW89EyDcK8bifzuqrX3nFxQUroE8678725yRguwm3vgRRzimwx6s6kOYqDqmMlMtwqCZqC
2upQbipDstlaWb8rGhUE4lkRaGZfBt+pCvZtuXfqiBTa3Q2VYGIyEiSSjNUWBzTeP8OwjJfXg3xs
WqLqS4mA3hzRZ7lncY1sJAcCa5bDL7a1uwl6+zQg7/LbPVb4XlAVPhD3qPns+UlGi/soMnER3MJ2
W8lSnmnavJ9yt3X4XYHuOhTHoYE+HFwGvyTpv3/eOg3oNO+pKPTTNkO8mqh1E62Q2q3umU39Y2Fq
UJF6/p8C/H3mUb5hTzrvVeO1OLl/AcmPFZ+GVzVvicisp0qf2IU+W4PkY0T9o9IiAL138GcYZK71
uS+97ysObJBCAXc9cGDGAWqt+OUnwe2Aff7kOLpt+JGKlYAxNY4kJXpLOAYUr39RKLb9HsiOqYu5
cOFM4g2IbukqcKHgiGOK7FAFhD9K6TJKjizvxqbMYq66SorSDK1gqyVQCv3cf40ul7cWUVo7jbTT
EDUViyOzVhQcALhr0nuxGhqO8qkQ8/1roD2MFkAKcrhN4IhgznsieUs4fORhP/pXBLt0T3cppefR
WBXOq83yDnv+gpCKFvmus59PdFwSrXjh1Z2NerjcTAa8ZiJAkx3JnnWvioJN595ATMfNZCHEePqA
8jXi85FHFrvE15s4tHHvw0aJUc1vycZRr9zU8t39uytUPjSznzni4NmSllnM1FkpiK/E51FyzTFj
I8mT+8JDDQikUY6QxDwg2hTW5PXXmyvyuHgX0AOyK02Q59qvLasAoMtJjVmrNFPFPKilXhLFGpxe
KUa+PEbcaqjrWke3zu5n/2aoJg8onBEpP+B/nnIG3juqwHWuhea3U6f1lCNhRY0MOMxbHBt3eCrW
UzBou10RgJOhpXml5C+pLNzge9cUfs887Eje/ZihhKSoDV8t9FVWK5gwxpIb+RouythW0hMjuL41
LLP+0DiRP55jouKfmZMTPbn6j6Yj9dpb8+Dsuyw/zyThU92b+251u7ptDueWxbHjTX1+fSpIPz+Y
bRTbGJBKfn0WH4yJ27OSxhSr9irMjXoeUmc0qon/dmXEYgX1OzIZtM8kyzHjl4A/SrsEXOcRdcpz
JuZfKkxwuUijyKQlbm/z+Yu9INpDC7Ho0ShbHwb1AVxFrzp/jb9b6FjWJu3Q+qxhmsv8InVP/Qtr
MIGlw1SzQ2TG3O75Q3RszJXCCbNOn6kvAFbGCwKP55ZBRQ4ZJWG3TkBBWUNx4J7Hkb7Iy3KoPZry
u5PgE0C++wftsBuWZcVcxUcCWuXHU1OJlNjAnBnLcYWfh4babDfdJkJ6iSYzjpMn11yCImY1A2S4
Oyf9/T2lIslVdLqkhaM0NXrUqXmrBOVdyTuUpDVk2I7CC3TXoKbP33Pi3R6MlV8zGimoPoMoSGxW
BXAQhqHfTAOYuSNMwbyD1i8yxkS78Lo2UXeQYS5xygWZo+lA4Gk9C87W1H9D4W2vaW90KJ4Y+/Bi
eJ/f09D3MJjuiiwn2hrG1ZLM6HGnhSps6Gfh0C0REIOBUNrqLU1g5S8YmPP9MQmYG7wkHq4P9ghu
VVio3G0PWTTzJYEtzrT5jNkUtKB4vDgnOiEcIXj5/CIWKE2JmKoJ0s/wQibPmI0iPsFTAyWjNFLv
JWh7GCq0MhbTtayqKpInQPDxob2IVON2zFP2hJTtCaGJdDKynm3x/izRljnT+fhJvpyDSguMTcXS
juLJkx0zNq9Jm6V88rIH2Q5gYz/AohGaAY1WiMY3slSN70/DQXVYt5pG/rMlcH52KWh+569C2vfu
i7qUd6mhwMbnU0al8sZq79HiBwDF453GSxLpt1/Mf4BFwJpOXBNS+3laNA/pMVRrWU2Lkg6UEuDj
gGm9t460MbTCkRoBzgHHIKta8Hp7lym0HxhoX1/gdGqH6/Z0Hlocnh/f/bhFPbepSPuEx53ODuwk
SC0v4QYJ/kNDYisfnX1dqOiUKgcBb9PcwHIy4C8gAa6bu/0vzLJWOvRpRuHhe1mEXZEmXy2SKZca
NKJ4VJ5x6o0jAAFZf1gnoHsTpuwM7LD5laZUEFHdh/dBqJLhTRuL6ENL3j85YM27l3YcbRIJbKWE
Tl3TMf6bRJ3AEPstX4RCNXlsiIlll/ehr/bpmrmGskxEjBb69+c0xArB3xgeCZYjMp+LQ2fX8Bs2
ejabMBwL4flSfBPEoVIL7IiEtXsXt2OASgggSTqtz2Q3cBLt7oMmXxGAMEDQ4XJ+SDOstR7UntZS
MrJ8Ei/BrkzWY+eQqRQG/eEtdiCdfzf9jjCg6M6JnvXD2M3vrKBBxJ7b94ckA1m0x1KRrQuyHhO0
K/ZRoKaFtXzg78bKxv0lhE2EfMYBIofE31VAwENVAdUAMv+lgiZP3QQXNuoWjQckBS8HYtYVRySt
SIlMn+oy3G/9dggdeWYvhbihtyljSzLNx7Vo9N62mL05fIqZge3eX7YKt7oqa7RZW1NaWT8OR4YF
RW8VXWkPNTA2buwhcHxCcHtaIL0RT/4qmJX35JkPvcs2XRYFxpQwQgrjhRNgLcvztdo/VDLXA7iu
iCA80P5nsNBKpamqgzcDtCusAAIdSlqTS2TQ68C5knX0t+Bn5APnpH0XCsMtHj1Q6kPz8hKRJsvm
krm/FbmBsJYP0p6f+uugYyjUOPIGm73/ZMGNGx1t7ej0Prc4cQWS/zAxu2vEutITUkFnCWzlYcAH
YVvEFWTpGKnchj2kSvzgZNlsV8AzobhyIC3ikmJJGLseoEuH1RyUVPC6cAd5Wr2xdttn9swvh6z9
y4SO5MMEB5c42fyCH9dxJTrXCaMJT04MtVXDUpmkifGXyAyITg7WOr/HrFrH3b51zy3EUGtKzRno
OFRWhqiB2nAeY/i4Hmp442UValyJUvCGzjsKZQYUrQczlSZ0AM0WGWSaqsABWnCcJ+ioGaK6a781
266VVQ6o1pnGGNw3uv4K2iBU8qK42ajhJPpiJCbCJT0LTvEzd5zL/vo8ytdjGzhJfKubdgNw6IbL
HvmacukncxOQ1HcvlsKUsuGKvszfv6U2CvpmZjEfk98ntLeckuqcgKC1lZNPbUEyitk0iBQ21jfC
LnMz7UHOo4Vrvvg43pTn34dhbAwyiRikFgKtVsjcgmaaebQ5xgPXb1iBgni0KE4cWZThuEGRHjr/
niCApX77lK4gfUivQvCOeqiq4zAcGDeImn+1SSkaJMK3c063Zbzp8yAkF9nsdyGmkTwO6CP+KLNv
pzrbF7RdGh5CI47Y98kpbV9kqzhSqtCSMp5ES2PWaVEjbJAEqZFioNYKrdpd0Khb0HTIgn4lAeVb
mtjGZ6VJj8xOk+ebRGXr9P263li+t3xUk0xclLYJ7MK9uU5x+NZCVqw6bMaooqOs943lvc37d9dZ
ZF5JFqE3qUVSQDIaAbMMJPbCUZy36YyA+jnXi/2GBdoeZKKju9ml/lcat+9RB0LSzuemcNu89XFf
Kkynh6MOmboYVSMVdkwS2h5I/fkUfdySvUlONc1dQQH526UzO/ChmwRhhJzkQW7b/swh4Lz+9wN+
k7FJmTa/GEhyjviPJwMH3S3JLEGjP8Bp/R6SjsqknvT7TMWFlbS0I+DKvEA0Jb/DRQp32DNF3VfX
xMh3m8UfUeuDbXkUxbff+2Si651Qs3kg3qE9H47O7A0OrHFaXGH5H7OsgtTsko43+C+zOSnTnBxj
KGqT5gUmKDjHHXNVafOi9/OjrfgKNPBAI7A1xz+zb3e1JwGP8d8WL7XYRUsOBupH4vJedmm84lMq
VLTBX5TxEABaAYenmSohuMXGKrpmHoqovQbEtQaH8BzoVaa4YHtxXZ5UoCOw/wdVF3EripDqRbww
I4KbQQD5WPBP+wk4cjj/J3+BDjTovyhLOUpE/mmJVmAh1off4kLQdwijdTeCit5PFktiPxiTtk/z
nEts1bXqIC5iLKuJhdUk/mFNgbpUUvPnTJtjNoxmFNFlH21Woa6XPU/Ch/fl/iY15PEq8MfZ2Opu
RZ0mh9AXcft/DNrY8skln+UWhge0bJASRQTgaaQK069OCZnscwDmA48T3zkKELKuQ6zYSDFLCS78
pb0SKrmJTgQvXrjBCMAf6/bKz1CaXjmAGV0m0i7NnS3dkNMg1N6n3AvQ32X3fS+GishgdqWie74z
fbYIswp3lZyN3gy+9UNLrVXi2aElqUY9yyXkdMfGIw8FzUuLXrbFbx7rG84ihJEdcVI3ZOwiUO9r
zfz7AhL5/jEX3BQUKpaOKIMoUnCJQI3rl64D/yKf/cGZuozBPLmrylaNTWY9WYsgB9DrBIzOsNqr
TExBGscWln13rqMhx2jIMsP4attL0CtDLcFxT2PF5Iq3c4yictlel4hNd46N7dQ6UWbHCUUrmMCi
2SKLMOfaVg+5hye0GLRNNmQXgHb6ruQLJYaUxA95+NjpaWtpII8RtDbJPjcLviKvbiMEhJV2XOAH
pg2kx3y/Kr3/1isoQ1S2fiZeLqGpf9XXYJ3Z70jRIBiuAd2K4PfjT9a/UZnDmJRqW0npGD0zUgOI
PmJBrUHe2cHIdK2sFVX1wF9AWtz2gF+7AADmvYmXJseYRJC11ixvjTnh2ds3X07kkF3oHDeM54TE
yBYEbTcuM8QWjbdPy5+zIUBXGZni7EO2xebsvHrVa9N/sY9iqi4+aYSoFw0xejzsjF9QOk1MKoB7
hdRH32nP36ClbY1ZXPoJrKJzNX977TW1e9oxdVputuq03gDqApGrKKA/5RRelKm7n+6+pDtOBwSF
0wi1b1NgjGej7WngrOfowuvR/NSXhKoTBjB2UKlhHqoOmJki7ojxtSun+T4HgNp7mY3RcFjcvMgf
epm0xvU0AE1arAfhG/C0/pUN7+b/CNug7aa7J2tMpXk0nsV+NG2QmPLgN9VO3sdftPRztE2wy69u
/tpiS+5dV15y4KRiurzLxjaCPCDuHq1WONbs0LbBugnlQZfMKOKdEeVdKWWaeOH1acQjzjr9PWvX
yqWyZ2zJgFrjKGBme8V9rBu/mcOZ6PNt13Kb6CDmu7oJfxo8tPBdTJPWJcWUDVlsDomCTQ6iqkgU
Am39hogX9knPIu0NXg3gP83xw1O58+rheQ7GzNfdkGQEoVU0dbFh949cEpyq2lqnTeDO9BpTsUo6
Ie6VNOeIOzXrTiVxIE4rjn5esF1CnN/I2nH00U6mt+XvxmrFci+vusQcVHapfz5baKn6zqEJ/9VS
flMR9v2FuGV5I2am6dpWyhkKzT/5adbDt3C702SZ7gVd4R8tQtT4fh/2IcNu3AKXNc44xmy8BukH
emlEq73SCk3LXrNfC698mYZ/y4U0MOsQPU7+VrK/jhji55cHxS8WoUOU6Cb2Nj6dw3sOGRSEJY3O
2fpHA9kgmEZGYZL5YyN2mEf85SFIxm97GikKNseBFPthPmK+Nqa+XpXI9P8eAu4lU+RXvuiily6E
EoekMbs2YSJjfL3viMloNGWEVfte+oRKhq8fR/bHv1oXP/4XRVuGFFXrSAqJg03hnMUK44dogMVm
lmePunXrSgEf7kOmUCWRJ0PapSjxhS0pAVYNy4fNM51OK1PML8b4Q78SspyKqW3BYmbqAW4/RCjL
RCLPxGsLSwbbTcXNn/Uyw5dKxsZE7pT0m2uMXoP55AKKv4j90Yxalu1Wm47JqYnFi2cxsBC559OV
FYXATn+0EuZ7foQnsz3v+Bu5yAQDEwIlAA/fKN2QN8ladHwmBi1X0HcX8Cj+rmffq721dDa68sGA
qlLFxw9SDHYkkTLdfV/Lg09Rf8HdjT7B8wBQ1/pTWoqzTsEKX4fA+Ds66eDTqnkbe2L97Qljwd0r
UWLBKNKXCgz93MuUTTc3Q8pcfTkIPP0tBfvPHMB4/dueH6Q4Rf4aS3x1L3I/9iItNv9W15vrOqqT
+KAOt+OhQ0Pz1mvtHIgmip+ctOtk1fYyqpbUrVV4nS8RalQ7Tipqbl2HoZszTDvvrz2HMbf2x8QQ
tQFw0YBRx+kvDVOO7ZoDLNgkxCi3k70+Ji5IQF785CKf2Fo93h97G4yuH6YcXC5Amn1gmR+qDmdV
3B19eVR/7dStPQFe+x5TAX+5K1eGfuj2uO/oqqBAqdY7nmAo57Nex8YPkkEPhiRf8yTa+SlMx7SP
UfImzKhIVONznEF6xNBlBpNZI5usLyL0ZOv+oTvzZKFRV0JS1n4h1+5nSCmQ9zcu9XNtUhCf0P7j
d4QDIZAYutQJIpwCLBftmJdRJ4r5BABNoxWe2ohJy67h3ljKQlknrF8uF832D7X+m8QjVJIHmlTc
rOCnHuGSVEh324o99ryClVpr8rGNdvObfTjov9BhFGF2lnP9JgigjvvJhXhkJ5yJ3+aop2bVe9A5
IbVJr3SVyptjBeZqOu62b92//kGwoRGRlIc8ToimbPuBQ2EEW2QYY5t9NyZ6IVjfft3A6+7OR1WZ
5R3LpFfp8qeInZrh0HC/4/1WufIWNH7CZFaD6TQyOpwznuluaz+cIqZhDxaTwzCBTQeo15KuiAet
GZZSJfGQ+iYFZLOpCYiP/JRZHDedNSL3BROUAbnDD1uiBbZDfR1vcmosZAfisJ49SafLYYRl6oJD
IgC60r8Dw5YWRhbw2T+W0HwQzVrBCbU2PKq4vMz2NAHSxbyLe0pFIwdJuq4hwvZTb3CF+FNAMBLD
xDIELOJCGKh1g9nWkKjgAg53drgbcpdemkFG5QTNFSUltOr/cIFZSIBcL5vcTmByflVAmXzOL8Bf
GcS1BhvJG3chSGz6PpPIO+lR4+FOtMBhhIhG3TvR+mnb8ctbET4/gt4pqke/8krjvbc48xNSIei+
5nhicS7j7hD6N3jzByr/G2t6r12twSWZJPmGLJgfvyXFv1Zu9cSqzf3zaHWWHjyHYLwrwwuDb1TI
LXomth34GGwTJl+8AyZv5f73P+OmbAZXGbHD0mEkIMmLwGzi+0xMZ+FB9vzjtvesUh0fCqvWYzxV
hLwsMxEfd2wGhTYVxKlBXEvUlgOUrwQhW7A0g0U+cWW4+UsQL1xrbddCEygFnm3uAkPu7MHSqsgD
HUZdfjl9un0jhziIub18CCmLDEbVSyPYPK3cXDHadVkir9ja17biFv5uEJzHuuefz+Ots6GLpEM/
6/zQqCyszaWewp98aBOITHPKnmob1KskOG7sKiqelz1QqUQqkO5eTACT4n8Jh6ZkqUDTvdhA2oaG
JDVnTad0ZOSQk2Y+k72O+5tEZfXfQ9g77LA9DsxZnb1nx/nHzjsi8tHLre6ZP/ckDU4tsfZ+h/TC
ggOsP4RZUOdShJ55z3TD+O39cHbXZX4tmWfJS2QRdI7uKz8M4jqBIlsViLRihDVF2bo0auihGN7J
UrceoDlqnaT9ARu7kv6z5ILEZn+YXovwCq2VuV+2lfl50jouxYlUYSlRStBqEMmkz/7QYIKuwC+W
OdwHGyUMmNczRKC9iUxCC5lqeHpX0Y7QczwW68vBZPr3PVdYhDL24RXG8yJnjE4N0lUJL6jKdCj9
F1G0/Etc38fK8U/Jo/tezwUUg4nBViz16yq0VFfYcyabq9+kfG6xnm0jHpj9yHLZnczAiqG/a8B9
M/Z9pslJbMqvMngkTdk7So6/bqBzEC3fyW0vCVFWJLDdN8ED7kMBY9A9g7ashz0V2rEID+aHLmzQ
xIK+0Xz7KojbbXyZ6iCfJRhj+8r5CvmDDXQprVQiQC5JckBaexWQAKaNPvXg0SrZ9RXUh8Y5sbIm
ceghhNgdEnt+RQo2PcIlI0+ROcjgeNn/OV5QEpWrt5lgDxFJz1MzP3dpLJ9o5TB+eafH0796BwqN
ongq79Ut/Fej9sZ1ITFbmCwMP0kkPuFIgZnXmp/4LKCt5bP4fVXwBTf2n8m9OpoKXTInBQjkuDNR
WGLUnf9s0WYBvvd8dK+U/QlYND8k1vN4C4MdGcGAoviMlpHwcSuyid+Id9aKPpc9DGHE53sBKN/t
Uor3fo6kSY9xTBrYrswntllb5zyiqBlxv83O3mvM6gsZ84sazFIDEXsz5E6VnAoCo8yKFnCqnF1l
1K7xqxSDw8MvAYGncrr6kmnY/j8f2Hb+qWM/iA8s1L3wS7wXw7lHjwtIWSWH4Zo2sNWEBx0l47tO
EJ+RsiXMHlBFPC6v6lEERWwxrfEmrWjFUjLXt7pCBJjODBe4rlGgJgmHBnDHT78avmA3jaLxii17
hilnf4ciYlS5ZUTDXIO2g34iGMOiFvEGx+xGtp9hvkkT3RKiaz3e7slkoq58VEGVNgCAlQGr8UPu
jg2XIZBVlgaAcTzuC9TXvtrQv3GppPWTxbOljABVeidSOaj+RTjOULV4MamqS1PBW5beTuSllEwv
8DAwntQXGW7PnJbwtPWlAbX7ldPKB0GKcd47GYbZli8J7O3aF6IHH578DRpbcsgpczP/f6gT7cN7
30y7YHA3uWVWGMeaV4nhwY218xrQqrGWFVL9bzEYMOAG0BL6LljROwTNoe8G2oe6Gjco2R/6WWQ5
tBB2miGHLw3GFO/JUBgZTJzgkMa9EEIHUz4PDxb/uUy3/yrJM78yHQi6GcQ3HDZKLVHT1J+0ZJlA
pg2dVz2nyfUY4KnqjP2w0Y2nwKWOM6aWo5xkvgsWyed93ta8rfMnSk2Oo0TzetFzUmUjgB6uRXae
W7KLj4OEIsVJfcGehYidrGhb4mqmGKLiVSUSc1thw2S6vOg6daKB+n+cgKUkbf7kHhM/qUlr/NFU
ZsB4k/yTjNy/PPrjfAjF2RN5VI8R4JUbAfEnI810+AAVOYn4BoBK8LV3ZYjjFhqN+zexMJcuVS4b
jHhU1QVSLGJodfshG77ep7ENvC1PGjdPh/pMXf9elQg6UTx0DIpfjvepwdTNiLGgL3XPcvzRJWA0
+/vH4w8x9E4c+HqvatRUPnGiZn/3zhmC6gRugZ+/byZP49HwFr1ozo1kMA170Vb0fx8I5i0vCm1I
YNgo6HCCarECPlvA/3rccYPGr9nnfofEhbSX/NvK7mIMsWONziXr3kfTVvoHAxSejttfVGSWPD2J
Uy/bOz5BVbRyI3gqpXScROtkF/YtNorHCdzn+RnBXZT8YuvAP67iMIV5ZfWDPsiDAtrCjxxHswu2
4W/euK+X4H5E2f5f/U8U6C3EmTSSaqPaj/RNRr5D5zuNA+apkFUVKa0xHGpFeh1eTtM2mW5JaK05
SRdbs2uIDZzUvnx+cRC/bdvpizpy+S5Es7UwppqPMk4flUyJosVolOXljEKLYqkLzqHuAoFAGSi4
rWDgndiVVkyxw8NmvugSwxcSZwZVIFrBpVFeEKM2GGiJb1faZwne+OIA1jWncdHDa9cH73BAi2xi
3p1Wpg1aKfoCJO8OfGzwmVlWhHTW8MQBLSu8hZuFTvXrOnSG6CXOmJHPrMwg5uD9n6s9yUbfA0iU
R6wJEIPbG/DK34psm/FgwPYcnuw9GOdnxxEG7RnljX6TlKOrQD4enRM7dmhVFsnBguwXwG3U0Jgy
ZvqrwitcYqa1p5Hf0T/83UhBpaSZm8WsGT4g81cg/NVhUg/4FHfwIpItxLkNOYdWMfR6tcLd1kFm
zhMZp8qr/zqu8igtvzbfT/nxPtjZbzWYL3PmIj5uDbCBIeGqtYJK/iEdKVHxGQfdtgThMJwrTlaI
r1D9Tfx5BOuGDbRQzV9b8/UDkx8azoxyfsrGuUQJ4eFe1M03dB5YO8sTCQkL07ImNXRnxmwMKMT7
27RfEDet7q6lLGo8aNRDgg1oZ51U9lIkO9O9pxeJTYa9WW61IQdrh0//SetSmm2nVa853r0bLnHG
NN/LNqVZbmhL7HTLP1xRNxOCY/6tl20/ADMtWBs+oHzGMq79GuT6Teo1eWz7gndiB+84RC1OIS58
AU4rEYjHVXsKYfTnpCfyjFVoFTnuTYz9BJOeT096CTRtUyS8Yf54SobOfcDRNRzKryKRvAzPKrx5
FSkR/wG/9co4C2VR2khIo3X5GbMQqb4FsE4xe2bifY5FkAGyhYhLd22dCS/2jGKjPErBQLCOebH9
JvWd2LuKNooAnGA/M/68zYVjVtSMLvEbZj/qTNGLMgprgJu15NciSrtv4OfOKi0EAxfjAihW0Gvd
RG04Z3NLh2Fl6DCOxtwQVJcU7oIAnyzIZIpyKXKF53FGDFVrxlm1yJX2H5mUBeBNdZUcIZDsDC2i
N4VX+acktC9qMSnNtuoEpCI0GP05X7BG2zNxS1XT0CbfYER3kr/A9ftpCiE6B+1Vqx6LnpFPudPI
mqwabIvkPw9Gd90RJLPlYqzVQw8F/Ypfb07la6Q+lL3XHjJWuRBrz0ovdyCO8Q5f9naNJeRBobEk
Te3mHuWknMLn3LzHZpVz/jGqy7Xv+wHwBdZXi72uymSF61eotLcSX3vNeiGocWY9IWt87Xu8jc7B
ksQC5sVAAfFjeqWxQGG5+3td9bcx+qLRb0c3ymaUngi9+Vrwb1UZJzKaSEFuZX53EkdrnbbxXfF1
jBzKvrU/xuP17Yvv0Tlayku/OYVc1zlw033uF9//IAkmhkjhw0/10vE31NEGqPmSAiosdUEt7C7E
+XEm9U3/T/qEV514N19ERLBYe2FbJSHqk1a1/JxqOHrc7tvNkZ+pSwHS06neaJqjoJW7L1Ox6PXm
1lMSyhhIAFCptcRDJYsm6esqeG1yYBuArDj6JSvM2EksG73+z9t+n+vrvbpFtLqXCEY8wqzfou/A
llC76/7yxpcZ7VVzhsQ0GvBBSPPHo6HsMbhgU7ArrdX6K0KOix8V6ZOCsXVsaWwhfhijvCgxT+0y
qMS0iDcZHGkvG4ydb5sDVt1Q4GscdgzPWkivBoLXHjj0E1L1Nk0XdGR2oUGBLeYGiXvltO5Q+2u1
8EdqU70F6nGcWNeLeifGmAaQB3GHEy/C2q3UdrM/6BVCm/AFW2CP5Lc+GFIN2by42eticMLDE/+7
Stevz6c2KHAuWoISaW1N85WqZcA34bdqBBY7pPoIOL40SzQUcTNIHs1qz0Ba+jhs2e+GhLnFT0pQ
+uzoMZt7IOeTtGhmklm0w1epWq8vxdlk4d0hT2+1d8d71PHGaTigLjfHsh99or06KmjC8OaoEaal
8p/t7mSysaltemI4VCWy6uRT0VvdOHQF62GUNLahQkRUR+ig2o/QopiiYONMrNK7do//gWC0DfTS
8RY2mAay85JVtwX+RM3nNk5OKpIrTm+07SVY1fIoNBr7pqhtEkXv7SlCYpn0R/xKUnidOghxlOP5
hsXpZS/hoa4yjkCojV8ww4TSRWnJQnx5A4WQukLc1CHxO4x4RBipXg4xS2zu9C+YDA0RcbzFJSYM
9o//Ct8mXEG348mlk/7nHdIDmfIEL/rEDvxHuhanwswgYeEqinFZQWdQ9S8eSPPTvu8DKG1IXEKw
mt9pPUy80ra5sxJHkBxRZ5EbKpeivzoWTzMNPtZZ26516CFrBwRwYKXdMhCH5BTQAL2ucXSDjB6b
rUv+kODnnoHVNGFsimse/IlpWeoqh6OqmZj1xPJ3M9cnQ6hbWC1N0sMy0Zw4nEm1AzZoXIWVtTNZ
B4cAY+gDiziOTlddezq+e/yKScin93NbI5PPjTgrjNrXvW3H4kdABgldSb7pBq1+Y8TxmrwPsNMz
1w8+I72weLkSc1hCdA6zsWHLvEylMti6e+DsCYqXGyYkILCod6rs4XoKdEcLZsfNXZLEacDlAxvL
zmE6tIWutxVf5VVtcB0D/11wKIOIZ95/Mxyf+6659jaCO/kIfyCwtpqtJpOULOhOVtPXF7h1FftO
vzEgpM/i/TrFk983409d0UHtcxnzZRGqnyhwHKSfvEbAWyd7n6h4cTBwK6VTyx3VfNS8c6u5mtwj
Bd1clyrM4TO70e5BrVmlK37gZeURgIwqm2we4b3JYywGy7pi44nt0LyJZlBWBv1Xy2eteDYR3ESx
CR78LbGHEuOfVdwaTKOObKd+Kdv3Q5jV86LgOYYm3fsJr6sb/H8yH7TDih35fw0wCkkvjSXqWbz4
pNcfvWzpt177t9NkVh0Gpmu/VS2yDyVYVETUJzCPhpL0DVxFdel1qRhVH425oflbs2rYqzZQzyj+
Jb9sfRK3HTshnFE3D0SnYWFvkuQmhbUnMJG1OMx2T3QH4I6UZ/lw2f+K/I8ab4NUhrDx4VzBVFAu
Wvl/HPGuhxeu+vBl6p7r1enNiHhaRumgPOySJfHoMfeRnVzYCEMJbjMzJaOlrebmtXLJPEFDgU/E
PsEVxff3DdAHGLNpYeko3iqWXqwiwb1vWaBnfZIOqmgeZoYZj8sZd9NDYN4kjwf8b2MHXOj3eCUL
n/hnWfpMk6YDB2CUnKDWjWgV8tiBhRCs1ynewQvcCxeGmwHtvdeYTXL6C8DIOqZO/JoB28sXC4Rs
1pZ76JXpc8KfBHL7rBdysKgo6BEp2gpvEQeXektnMLg462hDji7HaNUJrw6qgcPQJWQxKcg503d+
l5zAdJpySbnYrA6vPqTZaTnmdKuYqa1/SEw7ssZMlCoiD9TsoCGorZz8P7ea3yKqFlVUaWrhho84
Gpsz0I2zEcJVqXgllU2x+ns8tGxdCh6TPTHY+HnY0nvzZt1zuJM7Tvi7EwCLv3xYWFF3iNJ7iu+t
Bl8/jRgR4CMTJGWgRMMzp5hQYd82gTJAfDdAOgt1z2HSMBwqzqIMi4l1VCpNeGMLtwlr45CksWeD
7MyAQJIGI7zY7LHZtWfrQgXWEnQLYzimd0kd3AX18iigyDjH8/homL1to4IWxQnxL1hbpqMixG45
6qrPxd1czXNx5B7JUitTMaFEAm/8jHLkOe018bwD1Vjke/7fSRXXhyzLf2r19FuM47txG0j3CMUt
bhFbImb6Lz89lnqTPQnOaXdeqxPaJYZgChCeDngDyu6EmLJWDPMhO+3HSeLKbX3pUzOnY7T+RkPT
IBJlFyusba5buDIi4xUMuT4CnpYR+J87nHNGNLFt4vr6I27mVnhnoJ1q+K2EJnnLt/WqgU9x912T
V0LGjhf3MEFSEbXC48I+4Whoe9wq56iYlth9+xdefz1QqcG6j1OE2R9he/5QkMRhCsB3x8PKVE4R
XBJ3ujue9u71KpU93A+AnSeOqdRxx5ls9ev+hs/Wx2g3RVq0cSb9CuIEqkDLN2eZJpSzuW5Frocs
ZYr4AfvkY7vUCls4ftEzY1YpcHrmWGTWT8iI6JHPnCHmfDpyPLcfb37S41BjOqy2rx2zrI4pKoCU
VbSxL4ru9uBYyKvo7GCTcHxErlswhrUIeiPzDl/SkS3UBnimDOk4yd7ciNSFPuV0bQGX1sd8c8wj
olOxK5KnUovuFvODrWP4qdL8nAjfvpxs3plvJWg9cb3S8wG8JQMImP3Dlt2UmNaoshkS64E+/4N8
zimBJ15nkdP1sGd18vjCdXVbKqhWmuW/FvRyHB7liiSmEp6/u7rC96vxK/tSzgbjMLlJYK1UcjdF
kTXouo1tOAteOXNesM2UmeGT7m8oiOoZa2M7gdnLmFQXdt4c1cmS5GtyAGs+pKve58em7hTY4+Fz
tP8vOaTXbvkC+l3/Ep0ahe1HozRHDrCxfvUuVioKoAJoK8XrxVOk+lvL0A7zaa6cycZ+UZDYuwaE
tvma5ArGEt4hXbX10alIBySauS6ozCY+CJBLTSiOezGDCmGnz+0TpM0xnePmyl+YWDCO6sZvkfAP
23HaLlvzktEFu5IWijI253EE/bRoRZtHnXmHRaGZa4YOjHU+vLHKkMP8jHv7DUVuv/mXGrbiQS2m
X2PO/o/sTvPMe56DKjoWZsOh1UQJXT6eDZtT1Nxtu1+uIx4+Pc+F9st2WyxajLGelFtGshfNV/0H
TckBRXdPXH8Sc7hUzyM28uJW1ZmmTSFUvqxi2xk0iPvUF9oM/ZxCcIcchKclxbdJtHuvRqibpf6d
uU3iU/E+5bQmEi2oZSENJKDvziG4bfTXtthBSWgbF7e3TNvHO1kvVAG1ZkwMbwx0cAUXzfxJmBDT
rue1BIMC+Iq18KV/tt3rNnFruVqL5ZYh9Qx+vnVppf2y1HNewHnEYIYRDS38to40EpUlTqjsaKXa
KKH9xd58qiksw1O+o4KR7pBgDI0bfG1+4VqzrjbQdUbh/9EocpTXguBHwQi8vu/eh6+nmj/ix8ET
T1UGt8xwkmuSroilo1HUIKOGsYHU6wc+PlwFRN00SJLeHJ8cJhtGIm+Ta6tfX2LZEZixADXhO4Tl
8xdYPQkaOzspBf4tqSApiLgf53DogeV21WuEPat/YjJ6aW8MW/BFTt6EpcmRsZoUEEzFRsMFpaMK
Gb+AkqD41OuqsRPleYFIeeDmoNYMMwaiqv+MhX96bQCS+l85BIaw/97zrWfHbRP4QMIXjlTfJbbq
G3diJQRl43d+g4XVejNLuq/UynCLHYDtpm9/ugeC9wP56lVWO++0b8JioHw91KR+pRotDXfHBy0i
IFHvQ/ZKmuKba5COX67r7y/qz1Dp4TDAwtK4QzWJZ8pELvKfn5VFTz0fHCWnzOuGaEBZZZxC1+5b
pIdW7xCS2JEDNNoVoM2RtcJrhRzxMkLpBWyK+kqbe37Ku734Ic9pPf7u5keddGIzyqLDEHL+csD6
U6rduJ9qG4R87CvIc5df62HBg/4LIK4dB9w9zbVXqDmKtrl9WxIc80bGPzA1QnFl/dQ13HbITq+/
CAZG2FQInwyzHRABXbN2F6ZMQUmeG6UGf71VMglCZ6SHa4OvGpFaFnAEKa0oIs1sAzj4BkvFbRFE
DVqYz1g4f3dMXMtacjQ1YB8/VEeafk9QnadMp1sAZcHd84cENUV79elTHXkKApdtP3lpoO0uFOBK
aYL1VlUM/vel4Lq1cwJqOIpW2OJ/P0Z/B2j5sHXGva48MGpaEz3010HVPTkA9yAwo/AEE7itIwyT
rTplkvhDnEf4Gnh8F/L0Dua3cNgPulojEuYKQNxvuv0PDMyx6Pf1H58pAtFFEmu87684I0S1QJXh
vq/WCgIJlxTy7t+3Ogvl/SlKBfLHL/BUijHXMmzNJp1zoos+7XbmN4w4YbgVr21rrks3WPwHytOb
5BSJRmAR38PXGIRl3OviEJqghyoQmC7ik+BaNgCWUIuaw0SKO5kUxghzsVNqoCwVaL9s6Ex5RlPb
rifyEuq3QNnEX0+GGQ4v5qYq8IiEjNBC/mDTbDgY8NXariWasfo8WAfqMFFnp2CtkdJvfkrxlEE2
ROQYEJb2JkTjlYJ/XlJJjjt3cJKXhxHVjkMnBCseURm6GmUgnNXWpP+BwIc10SofIsRcou2lThn4
T1HEznZNv5NnCPJqqnCSBPkUPPC2FHyoAv/+SJjdj/0RnVcPR+0mc7OlE3ydONVmjqBod4UTVD8Z
YVfYf9oKm7a4lMYkgDyuhSSGEIwvxcCXB47PYBU4Pq7BVUpvM83gwvDnkv+KOK4ImbhubEpm0dnk
Re2uh1tBD0W8jYIgAm7Qn8n3ssyYf8FVLIOJ9psnLw4UxIiIzb4wW0/XZKPq4grUfgfBlDr30BAe
djMSHeC6o/vjA8/ZOcy7/qVilRiD2FfVP+zO4Tu4GapiHahsVc12DzVLZ7aIzSQ2uioHOTND/9ln
tHpWZqetryVwqWNkSLfKcB1ixm5CB4jhRvQCycQCiCdgoTL0d4qWKBlWYHzDjxC+8x1o98KOiI3F
IluU3XVxW1FM7EDT4jSh0/ZJM2aq16QjlLCFlpsKPWFI10OxkEM/32QI6QaeFNXgq0pWDiZoPKe3
LJrKUZZzabRpvAxXToItfQqI+5Pbs9dy504vMGZShY+5OOqhnPGxrWzPBpoo0fxeWNv6JxCj21Dz
Clq6mEWGKxMzDPLmuxeQcWvlPJeILuJMpI+kfwRYeGpGNm3X+KG9CAJJsmdwiRIUZoZ9Qq1kUPOz
PoAlMbbiVmpArwRKWRkcfVj+7P0NGiFePfyvnRXCNdKFwOohVHAATO6BDNZV3Vrtjym5vXZ59AOG
3Kint6Yufh5/bPx29TZeeoDZdQTHnGZrggqmBhs9gxiQjm3yJKE0Ueyp9luhCXzlmbO93ez733cL
VobkwnnWQ+Gk/BwBxP24e7/NkiCloVPrOWuhN6dCYmdH9kpr2ftk6ODqkQmYgW8qBj22LPRlthX9
GpA9Su31PV1brGzhuuBHWdMJ7oRD2HaPtZrVdm0eup1nSkkJ5PMMNuA+xIG6C7sXbaQ4JqQjkWFx
evXOWSFOqYK3yU91cYWAzyQro69ObRTRt0n8W3Flx3iDYCL7oLTcF2MBT8cZiOH55EvgXwtsDHQn
letn6/3b5rDhW94IcAMLFgohXpHqTfs0WSVxRxDYfd3l1VhdOD5T7bQELT209JnQvRuB3P/8zdxt
cYlPpKq/kYi1YaB/cuTSip5HDC/U73110EsngcmO4lQopmrTglnd7s1dpLKTg+z9vyc5+J+HlLgG
FI7x522oe2pR4WoC07o2Pcbqh8dUDLBrKo5KQRdWXjpOk9w+G+7Segt0v5LnakCQkLNHPx6dlhsb
XMWPccXuTM99Q3ptwNaT5/e8QbKh0/TW00QSKy7IapvvScKBvxoaQbSU5DdfFShfT1k+LFUR/WjK
D7yuWgz1mC8N40AaKxUV6yVHfKhsLGYJcJLEf3cEPaybQfw0RgBpcc6qbdoyZs4UZQPKso0MUXqY
b/FCk6jSFR1UywlAYWV+zMrg2tzu1b6PUIZpRu2zl5nqXt8jLt1iiTiFKBAcpPVVZG79L5K0jNQK
Pbp2NhEpjce2URMcr/G3JNQ//+AQEn59aGtwFNaHqoGBx7vytjl8L5mXGJ1sRNps0F7Hwr3lBcP+
fQhdc488U1MpEY24U/zWmaQUSo4/octi2FKgwDqp+3XpppCod4KFzckTpV5ZfnyMliqzyPQUQF1D
qwHrGk1ja/GpuKDhrsXqmNviT/aHiNZ33yp1EbhFQbd8p8ICeqk6vut9PuBvEU1piH/oKgQTGeuO
K6ybwycdvyDgFJhTmeivUsvwc3HkADmzlH6bJNdjuACsgFojnQQp+XrquxpRnhRckIeTT8+n+kn8
OQwc9JTx4Dlpiu28rCYkiKITOUTGKsVEBYlBXTk7f6hbq9QY+H31P8gaNknjMMFoNHSFO2SkQB5r
zZqbul7HpZCxLf9QjDehEfh7dPbutc8HELupPuVEBhAn7oKSnz/S3JuqDFbx0UvgLgBJ24qdKBIV
Rhi5X94Brcc8K3Mrao0bLXO640ryXmuJxYoQ0THcopMtpVzzMuly9fK0KH8W/9yrPAmUyYBdfMVp
OzN4lzVPbOvBgxcENDwcvJYaoQiQgB8huJZm15KwUuN5JRa0YohcjYFOufwdEpyXjf1qa16whg8a
HjFKy2DCWcuLPbHJ4qn78hudjZhYM2bCovqWv5kL0lWmwbA+ucyAHL86IkpF5/te5clmDeoO2JGC
Bz2YjH00dOnf1WJV67gtQXoewVqhPP0RelS4H9Pa5SpOf8CjH1FzEoIIM9YBc4bi9de/HdCHnFDm
oF+t1paTVB+CRBlnH+nB22YmFqrCr6q0eM/kvrbJHwHWkFyDmKIV3CdhMuZlyFDT1Da7sSj7qwqp
+BY93zi6SSykWML2gGKWleXu1C3cpI+TdUh4JDtWCUAZ60oWNzlwMrULyJvrIqV81xLdme72bjqn
fon/fdSRAhxnRM4OO1YVITzKvWgCvykPn6tiDMMG7qVc+hjpATPfeoSqBms4/BWLRW/dO58Cijx9
n/NPD5QTgeyshnKh0cNhC2nkACLD0Ga/7aLMmk8ZkA1Q9ij9niG0ewQXf/HVlPTSyt5Q7Ji8yd8A
aaC/LsucIxo4wdyA8g84dhe5FMCjbfVIrd0OvuXEmgo848s5ZAKVhYd4kQmBHS8lIngyYB7Nr/PN
W8rr4FaEaIhyiRLGzqdG9hsEeF5wdHVbqXg3QjGBgAmREPEy/5/kKxCFI1PDPD8Bt0qrZDrM3Qf8
S0z5wh35DEsNqXOOstxKny1ccNOztLISjBghxxpTTB3+0qIsi33suDGnzJ7MBxeGfXkQwxizk5V7
ZVWQyandZizevgvaNNIQ7tfXQk1O+Z79x/ruk6BT/WKib7TLv4Xe+6Lo6tmT4b3BkS7SXR3TkKyR
n3Ew/068K+Cj3c96cW47xbWbb3doyD2BZq5gKcJY5zxHB45X4dtWjgH6KKdFsPzZSMQFEZoFzAhW
iN8IpWXIxG2awcwYgiyLbXdLI5Z8wwNJv2NeIemBReWqxUMTRqjWrKfQWGo5EmxcFcVYd7AydXx0
j8Hsklwj7cNEKjbrfRmTGPo5oTAeXK/69UI6cSE+0V2VWB2+x8sqsVpguNL0+X+7ppjqlrlpxLfv
VZEI/HF0zP37oCbpMnjuRPuvjuzwW8aAcqvacqNQIMhPlpCxFfz9MpeMR0geXx5pWD9gfCLnsUg9
w5KjHa+VMZ2eIcH++BECrHmTJqw0yc0HShL/7RChvsw6ezKAnkVzOAHryb2KWysWHRtVo85oSUPe
wre5bCe/8PgSdWNf2cZ70Z3t7/Sg4ScXD6uro4XobGVPZ7ZIrkNOJlmuwssFsKZmD9yJMiy3UdMv
qg2pVCl81+rzFR8qCXn4u6D4/I3gIEYqVD9SYIOQ/V4kcNaCI6TUUfGpP7w51EHYojS8jCJP07jV
ScVcNyfFLyKYysnVHKzZJVdYR3KLQuC+HInU0D5iLH8iRvRx74wtGIAZFZ0PJXWTy/LMmvJp+f56
nEV2fJ9ZWkpuorXTQUxPKYppznmV4DuWbMsKzfXdRqLMz9GQuXpVvZSFg+bojvCe61m6uxPk2dx/
8iur6NfTm0zf8FntwYFRPxaL8dBA9+ePxBE/QeQTEU9rFIwkc5T/ctk6xiJv+DwuE38aaaIweaOF
zi5S2p9lW9oIQlxsYHMeAysvyh9SqoQQ0a/KSVHZgS6JY7tgJaUyyhdc7t0xzqzJrZs6hEX2jrKe
jhZcY4H/ko2yP2jlyrGeqANTfHfk3zYGpZXWYyV7Aq8A46OJKHqWX9ROyy+bC+6U0UJbB+v9tpqK
LOHzevml8V8PHtbr4fppUryEbpBvD1XUkwLn29zrGL/mwO2HHRIpltq5K0+Sald4NA/60yuIf1T3
PWxT6VtS+nClObQnYe7UvHqpAnv+LZpfqsjSi3mU5GB+jmm91OXxUTM5xARe1gOW8xg6P5J5mt9j
lCZcSmNnUn3O5yemlXsp9VMnoKdMHqQc7sxX+izQR7qaV8txZ8GdOGDu3aMtxbuiGo0lneAcSpfX
vG/FDe6IsFe2qJ/b/3zWjleKINC+umrXpT1YTMF9WLiimOYjIe0oUmiHBHDHeS5JzRY0Hdytctd1
9UhbXjBha9Fs5bgZ+tP6hNixPI+73kT22W/YqLSHB9f36d9TCq1hW6v3EUbOwj0ogxoSQRVoU5EM
iH/vWOUCEtP+swHbAAnej6WPH6luDwewzRQM8kmalSoaG5pPXgTCVvydkBkINe3PuO6ccoTHg8wA
cE11iI2vzXYubZqcmZ9HHgTZkRpE1HpCXRpJLOG+lSxtldv1MFk2Lv4M/CvWVkLnWutfE5guT9mT
EjLiCRJRz4oLfvWj9kvyXl2TsxvroNiREOC7NNH+z3ouy1ngXvZ1+YVitm6ig8Lp6mcZWSYWQkK5
7GFnD+wd+rOwg6JMT7No4pHitabaBcR56dQ5OsqKTd894JacxyRIsuJf6LSKpSd11/Ejfcf2oheN
d37nA7iYO0oC9I8YDTjrtxaY4BsfmRJUnX6OnsfjNRHEMrmlV7fodwEEfYLHvRxgvFSQtETRR2dz
npSncNU0Q0rlhrvLNzpMqawf4Hp19vmx4qxerRrckffddiUU2L3B58XB2pXNTEhaOjz7LXfFtOoY
71xr/uNVZcH4cZWxAmUD6aXCOQjKhKIsFBan81WKUoGmB/58Akh9IzhXEeMVYdUxFraTT1P8shBQ
I0Qh5XfNIcl7wKYkO8O4Kc7J0HyWvQgkCEYbM2n1FNW+Obmjdl9uClblkYQhxZHXaLljVU1PByFy
C+2Nvk2qeOenR6ClBbGEp7OgEDMRhyuouo5XKAbfptoygRwzvECQvEzq7hLxtpQ5GfFS+oQtsZmD
oUsaNAevMlEgGd7tYfLUkPIgS0sGXmrUiiw6x/Y8+JgaZ7o5o7OAOEarcb6S3oXJSTiH/ZRkbpAD
hf3zvcrWzE8W3XHK6QgBQ0cN19EdzQLNA0SkeXVaTkHGqiZz1q3mIq2lNJuZLK3FK6j7RMmWcbCf
T40ttfY58wS38zLmm7hqONcw3WAgG9Cqc4A68mlCEBab0JOm7v/+CMw3ZS1gF/crSJzDWIBMgfeM
t5r8qfiomYSkbQrngoLilzaXDpjOFvXQYIzKofa6mDUZj87XjnEpyPwk/uGFgjG/+23ZxLJa8H5A
SbDwcvidyyUVN/vM7JLrJWQ70xv0lsiv/W+1bi+8zaD04gtM8lLwzGwTRQ34DXh868mMEY3K2dZY
ySpjxsjKtNhb7kEMfl1bK+GTxptFoY0M21NLhFk5N9gWejWSk8Pl8QEcoGWj266XxqBh/NwqtkF0
L0PDZmJMXo6VrvTz7s5QaSjWxhyGbUvb4gq6qaNlaaWwdaci7TXvHeAVYgi0HEk77XCjoWWupol/
Uk2NBC/Y2pAxMbHWKuYJ6CpoyzTkIo8+EmDemwn0++hYm/REHlFZS9snVJTqqDR5PTOAKcsgORfm
QTYOgTGEZUoVgSRl5dS+u176H3dN/lRKpzpForyEv2XOoFS7bEcImwdMOmvcvZQ3yoHCa5iWlaCw
g6ghv8533tehqBZKBsImKp8pNKdrKpAfzXRaTRgua+YiBBN5MLmkXmMvzpchCVV6c8wRzDqC5aKH
4qMGG/1iGWcfaZHEkJNdEjGkClyHYjvUEoV8iN1DqxSdXfwe9BpAGHAKbK4LpMpmTlXzBKYO1obs
RuVeriUgAkq4KkZMOcyHzifPupQCl2xEoHONGIJOc9QRqg6vhexNScgN+Qqp/nB4eto6tgkG1fbf
pIlGn4N7gMAdPBTkjXOqTMMs5yNUz2ogfDohTKFwP+wQ6EJjXYcZSJJV+Da0XcOercai1nH8uppC
kqXeJCXJzdNEnuh7tMMD6ya7IZq/0YeFjBEGC7eVjpJeS2LHGJwoNg2qI1UkrvpkVqEW9PQWhs3x
x9TMQfAgKhct6ylMErzV9CKePWFz+WCj/7NsGVqYPxfInmLSRnMeXpTB8JB7FbB3LkOKINdinuVa
zlabIj5nrjg8Js16cXElwyOQqc4T5mUnM1TkiqQiedYPSYNZtUE18CeOSz1oQiS5z1WW8V66mOog
FamvkQy81XC0o2Brhk272k+JCau13NyZQMhBmqeDA4eRpfe5Tq8kOII/HdlckALCp2ysV2idtSix
KISHNXXtmFUMrksnAa9ym2u0LeZ7LK0Oh02BfiGFuK3u6N+1l3ClV883ryCgJqnR2X/YGIWc0efj
3Fd97aue8fwBaRlRErNc7u3ZUdQl57MMXgKOrmJX35nlDO1WSZw5U+LNzQ2Gzuu27jzDkfMJbS9+
d5HXkxPV+OCQGXnDSZbEWFKgfMOfUogpPAFiVCiLYdVlKls2grCV8x8JxES3UO+Ux4/nVdUi7hbO
X4A+Hpkn3qOBWF9lNrAMGdkczzpKdDV9Avm2+Iw4nvErJeq+YoCBkHOEjx3SGA7OmtO8ORWQfi5q
3LPExD3sLsXITHAHsisVJXLF8EeUKh9sTvL1aaw9zG0QVGyH5HY9hu++tQCCVQ7yTNgjhYkITrEe
JhFVpECwtLuF4udA7WwjhPw0LW9/0gAWr8tPaL0Hi1CrSLqOsM2NXTEal+OFoXD4sfkOVZ8iQTuU
jSQkfg+ysKghOUjXJtCyXMzy22M92bHwwWyW1P6nP4Sq+aRxoiLJsKpZtFxr1obBVTOzbAkma8Te
kz37F32hf7qDY1BtLc3PgKRNAPHK9CWM3YqoGcCPdTaOs5gP4dMcW0LSTMyhVNMVl11FCjxOkDVF
qSFfSqzcTqUNaO4qncrxmPSQDA0iZ5ST7/0mehit4lsg/sA5SiJpHHved55Ti5CWcRrW65kFMbqM
9jDCbj1L3TiHInJBnXNsZvgqEUZgw/9ZMJMmp+apfOZXtNNl9TRNeBlUW/h4YjkxWOw8EXBFQrHj
R6LBUQLw2CFQiRqxP86InXWzGSx2CWeapVrKWWvgyl+zf9z274TG5bjW7b0d8KCsaKtHMXPacCgc
h8a54aU/9zVNjBM82znx/Nxr7mT3dzLIL226Vtir+7rIC8iYBTi2izrmFy2EHX6XJjmBl5lJA8S2
Q0JZkE2Vi1mDsvk2Yl4VExUxmKSsP8raopBUgzdU+wM1wtc5k+1ExgWPfghMxzO/gwD6PgAil/4e
r4nrUvt9HiaEhT+oyoPHLiIbkkfYxwX9vg+OawKZju0LeJ6ovGE7NBLO1/w1MfAsmtMJ+2kYkpEo
u8dPqeQu3mdDGhtJSWiGc+erpKvbOrXAXZ5P8SSTu0GxR9wclrJ1XN7YTrRiE+8T3On7mo4jf7hL
62NfhVFAGDJIumKoBM0U+6pp9SjAd9PcgDosyARcs91Kmcuqn19NfD+94GQdDyRsj+LrpJEIe8xd
NgPzDFQ1tMNK5ovK3zqZ2Ik9XgX+ejolivc4OfSbH5t7Acj+eisHqjL5FBhWGqiCe7GlkA7EzUYM
LIvgsVgO0C9gx6ED+nyxK/NXFyZVO+hyRsXX7hzApwitT1irjxKbMarjhglVuX3TqQjALa63vEwG
rVo8cWSHXPEQAdvcuDI/aXYSkNXWrdDHr0NQyoelW49xyrvVgUUAsfUtR4yuJnb1J3RPQTg443Y9
WCK2QLx8Q4sSBtmh5pkRItfSEoznTjhPRJ3krUM/CT6OsYPAzvltEzEEODv6wM2W9pJg+IKCUitJ
JjqjH68NOwVM9L/iAjgwS7sFILl0GYC5BTImZAC11c9jZknzZT1iLcmZgiaHzNIQKrtkqJK8nT63
fxby7XEVqsxFDOG9V1f2tJWgb9R7u4BQryzV8xOprUU9gXgANKpQCrtg6B7l1qfKW3zWWUxF1e45
pabo6Ho5MPsm1iwzupP3NNHD0+hqfGX5VU/Rl2NnGMdgWpJ6ORApvdwakLE7k7urlVLV4fRrdGuK
kCbMfFtH/MkpSCvOo/Ugfi1ZZrVR9pENI1WS4qk4LQ/0VfcrDTzCOB2M/nncHK8eb1RF/Z/s2gCr
v5l0whS7OzBVcjkaIS6+Of4bglSRnEk+sqyML8oQTjlysxt7FxuGvRj8PyAeKof7MCWdlK/j/H8A
BFKnnPrAp1TpjgrtAxrJwKIGbO4ZSybFUoP2RWZUv52ZMwzxziWaEzXOVBfmRy3aNRYzSFksUcTF
WVa1W+u4bHQAMU6/nNB+vjRpJjEpdil2GKFQdOK0A6Md9dhF56y4c5w7YKhLdU7oVNYRAX/2XD6u
0FMR1XuucqaOPkdUeh7pkHXKp2L+LBxeUpXpWRCNtvvP8zpa+KJBM3Y1re1U2bf+wo5Njp3RlLbQ
jffXyKqzq8Fz6dSlaroceeAMRlguqYKpFO/F077VD1VGETzXOPQ3sqtuG5f5zKeSIuXEsBg611M0
bDBrBdqAUEoe/jNUnVKDnXSeRSeRKK3czdhFQ36LefM3bO93joXFs+R7qinojnKB/O4LkNfnytQ+
CLQ9btcFTXJSauAEDwUKHMQvi5PBfPFn8av8QBxMsxV0zqh278M8IRKtaRXORFlwiWQXXr/W1kh0
VCj/JxS2ux4cp9fejccwYceKOfwPQpVwi5Av19LH1wu/jrr7GkhNfFY7Bm4Qzm6+kMq5a4CAd8mb
pj2VAcBdbPITctl8vdvzdK9YIiurYb7elu9iL1C0tyyZKYqEi4Noz0hOTXWkNRnEoWAKrtODoa+i
7lB1ntigOSuU4apFoLkuCkH4yE2ItZiv3FDqCBpbswdj11BvMoGZGao3DhdclE3jhWmS9xKCHj1t
S8XHeO0zvsN85AYQ7hJMoxmwbTSndxenCFXXnjR7ItDUOjxAlCJXY6brelLK/ySPrmISEB5yEt+c
z+FS/NtEjoIUL9tDiuAH80BgxXkvNQToCgaavl7/6xIKNZAeJ9t5omqW5V58WpLZJ56MHdF5fOKU
HZDL0KIYjaHH3OC2+G1iyFIPSXhAXh46C5L/QDtzGNiInjZVCg51JGPdhmMKLqEmnXKFEIm5ZPxG
qRYhfMgW2EEXp/0arFqAUeEY1GUebhdNGVmq0qBVBjlnleC+GJuWXnHUaUxwl97h0PMLZ/BYJQ7U
8/SJxVGO7ZFzZK+89U/avCWBdGSDs2vX89RnTz2wjbkvUdtKCBKT7ltuL80QSLofFRsclGT0Or1o
5B3EPyCOmNcfjuDcoydZYbUCoGXFqB+WCgV9Mbg1u3taf8mCwtT6Wz73bRqy1pDU1QWptAMnryZH
5brv+1FBRb0UULbRsvW912o377erov5qJEZc5IQQw9Wvn3DCCOr98tF7uwcGL9xn0xewr4XfOizz
7yNNpIr7nLybYCxkonSs1uqJ7HMCD0eooF+5AvWj4yLC1QYRtDu1z9luiRRcz9yv0jDTgXWMSW7y
p2gqDHWKKellHeMpwoQbyh7yTLXBsy3GssG6yvXsmtqyH9qSDpdusQUc7JbWEHLAJhdw8N57QW1R
kUY8YvEFtuUJ4EmXdcVwribya9aEPdKCZrFPiEJoOmx27CKqnLlwY727xN9taw5AX6+r/TRyYZ4y
7OosBVA2tdPnLrPHlLvS6wbZkgdDHper1U0QS89SI+z3wlulGgmS+wG0C0U+Ly7+VpIx5zVPubc0
C0wBFHj2wU/cLI+8jAEaF/pkK15LfpOxPRXsJnDuycEy7d/bTdb6Q99PDA6SRVUPit2j3LMkHsfp
crgyzqPd8R3E8cAg6SqiqemB7zZr4Yz3zpmNceXkpW31WNfillGHvnVM7BMXIjO1WCPAwEi+fMwF
VnrgqdIEbsad9k7WBuPFLp8LWxYXIKzd+wNg4su0SX9IbHMg/uWY64NoSwLfMlh3NL+2ewVvy6Qa
4RPuyOVXUfPOhD67DQb2+FAURDxuKc6mFCB4nIgvoFG31z2DBnCk2qDn/QNqijwh7XfUcaiiHTSd
yj0XiBnwerSsgW2pms5EyO+M0FwN4lrtmrU/PAbrOpuTCqPJSO0AjoRaRgBY4BcZGYsd5gZgfkFC
XTnwPzp9QIZuRLcXIuV4gEHeZ9oLD1eIHGExRL9pc5wMXEsIYzO07PeZUnjskZ20QG7mjJc65Ac0
TUltC9U4wwNVzm++QbCUfiw8npQfk2had938tPtTglv05SDKOKodIySX2+5wTQGRZjOQX7rPILPv
+mYgEOLBGqqVgzeMPe68VNrbdhAEOXBY9Hu71/CxoJrXnAcqyyfcARI7iXpC6Sa+kEtIj+ZYhEjn
cWglZFIR7hDgFttRFZJPciKKdn4/bILvYV4az4JiSIXIWgkD+ErAOd2UM+CVlatpc9nh3sOcSlyH
JI2aTL2Mc/a8BhLGKxnKV8J6jfP5RmlnSTlBNXbb/MfiboYerrRt9L190h5yaxVZWh1Z3RCo3+r2
POzbVJJ66IiptQjWtj64hTslaiKLGCYmSwJKG+0ewzf78eSk5Q/IMLjbAr9HlkAQuE1r5WYDpCHV
O/jcfKRv0APHsKY3r5wIV92tXe8ePhVNVBVgQ/owgtwjA5hM/PgiuAQzrBEynu1+MNM4VK6lOALb
kvdywOkXimDG0ZTS/4QYzuIEYC5x7jsLilpNdLoKK4prgaJ9K51wnClUhVjt7PBu0Du4w6hQoSRb
SItEgV7avMHa3FRq6snIT0Vam9/q4TlNSLVrCfdVfSR40xQ1KP7Sxx2f6ThjYwre8OGxPH0bKSSK
ejGPfdZDV1f9C8W9TyZdCBgRuSprJKwfYAm5HIcB4Pb6u8TSyS8ogzobZnp1PtCJb+YxA6Oni1Ai
hqrk4jEaWQ/k3CvDd6W1Hr/f/f1W5+PqM95k2OmN/kqQ0u7iYGPV8iRJGBdhb+Cs10LMPGC1fGWt
lTZjuJqOH0reY1/meDjOCX1H0Pf5+uixj7hmd1KJWEJmHhq9GQDKNxf62myKXarZeQdtPR7naFlm
9xFi8k2NId3gEQAUcudcrI7MXG2av2a2dl09zp+TaIkpQx3oQi7/WyWxNY2qRBWi0lkfUDQ+r6cr
hnwqbW+2KqzPkCIfND4x2uqGxn5SEF87rqNk5t74Kp4rEuNw5RRGjMfDGZKrdzeQaqTeqE17O5Y+
H/KLYVuO2L9S+VM9JKFrw/42F+bGXNij/KkSsAlcgqVxjfLGh+xW2CDOOpUliOOKUgx3eUiYz7qM
Wkj067GUVNMjuAkKY07Mv9FUCuy5wpCiz4FrS3P/XfwAu/dDtQ4PH7ZdLv0ENujmbeCfQX6W8MMJ
OczLBkzWhU7yEBJKCkjYOLoboduLB+0B8CS1PvYZ9yPncIBEmh/0fW7k9SXPb5rv789l0Ffl1CMb
uig11Ju4ygdj94SpJAOAyJAEs1L5YU3rrLviVAr4vX9L6LuofmWcpiKys3cA0mFkW2RZL+3dDNkz
K59I04h8QxTBOPZc6nMxFoU84PXDnG8tOHOT6zjN+2/x8Biv+RPmIAG2XphV91xKR1s0KZJeN9FP
nbIoQnqI2yHSO0hJi/gQVDTjBmXPPw2cG1XFqGcSYdhy4OkK6FJ9wCC3LsboYwocD1XNZfmXIpQS
Nru0ijRDyrPf1dtP3wDffIsqv81xk7+U/sYbRT/VdKLfi9fsGx9QPHTR+wkbz4norTyDC1/Xwgqe
Hq6HUM02E6EooRBN/5EwoCYlx3AdL0rhRJVYNmdFPrjnTDiR69QbwCADnZA7ySlLIhfpQuO3J6Q8
ZIiIUi4KDZ8tzQFZLj2wfkYZxttQrOObGqDKzuQ+xLtG4chwmMA7zBezojlMHwgz0Gn1boAEfxbD
CR0g1so8t3ENvi6c0XzXZRtpk4F6M8wzX9bFYxSACWQiKKTAOexa5JD1JstoijXZ3LRYqVpT8xXT
Up85IY8QaA0gy6QsQRcEZzmHDwZg08/mFLh0sW3U48YTaIowXAwOvBNBedJ3qVZn1kYAQt2WhLIK
taL7onRTTvoomQm7KrsrfSAERKSaXBFVDYuxD/sQmJ05kIMHUtlM1T8j6T0MuoNrWWWQYmLKzMfz
7cJGZBxFajNEfbfHgNTYdrPxGgVGFB4D88Yh0m4usMnBhe95YP7Jpq4iyXirw/xXsBYNns4JEB/0
qWKvRp2QVZ3zdJI1RBAj7zrGuplD373OY/MxW6G7qTXBrvmE9cev2HGd7mnLwcKmT/Q9pE7vJo8P
pJhuHNK0bMJ2F76J0dgiBVlN45qkdiwlHciFJAad9imlSo8NlFsekloLJLomSV+Hzj7aetLP45kW
d2xpQikmXLZtbLTCWDzTtEWen1DPSer7YMiMSla/SXYjubn1FcwFJ1m1BWHq+ApWWiuYssHvabFa
0dYJetdXq4GEQIZ705bo7OZro7iknthRfxhLML640NqNW1n4i6pM6ZV4fGEXJapNLFWY3OA6iKse
MvQ5c4O4mOY5Et+FIv7XyH0vDeyFbd5K1iVBgCIQEom8KyhEJKdDEcNEIIwDAOvi/yeI88rL4RiQ
vDxxdL8DSeoEUtTfK2Vg9oVq9YKnjHEu+5SDzVbYoDFwrRbGR1GgVaTAvBgWRip+uODsJ8Pb2FYJ
w+spRb9fg7p64ud9tqVv/i0ZfkUDVfms4EiVYyQFOlCeWZVRh0o1zxXbt7oQvOTGtK+Zi0n0j1mC
eHqFM+HJv++ShmbaGISjO0B3TgfqhlY2hILR2b2wYs0+QBdOOoQ8NKxn02646ODR/DWgu8vGc25S
GiI6Oi95X6VG8X01d37DMjj6nrWzOTxhjft6j79lvh8KtHyyhEh/DHnSihHPAMkHJ4dm77VmaJ4x
bQ3W0EN/OxA+lRZuvfdqFwfql+UsIZ4wYPYTWqmzPq3GQGkK0hxgyTGBh0lNVix3EPGNHi17diMf
A8s16WPwn61VbDVLftULOqes5mqoy/PKKrquFahds+Ruy7wHLEt8tKVwEbRZ4Wma/ORLBZ8zvXfn
o7tfk7rUN+k5+/4RRcMqjf5CNzgw++AYT9HtKfaziOFcKK8REcSO347viB09KmXUCx16/da32NwH
bJ16BMBTHdnxiR9eh68mgdzt2zRkvxRpY5+tb1GMffc6FXaUkyu5uJDk7aSwa0V9FLWY/mCjieWY
7loaw4F3U58S+d/YZTVrUMaG8ttE/I5R0inAtzWL4nbe651nJW/PdFUZw0Z+66u6lfM3jVB6HkYR
TEIEj6HD920BmuXOUtxONAsVhMjcriYkzlarlYeCKIyQHdJwV+BAqzO7DhiuJIAzsrYc6Ue/Swo6
Ye330fbtMhUSVEDnn/cyhthwELWi0jd+zzu4u51D8YtB35kaQAa7rvp84yK1TTc5eqz21RmfGHe7
L+N78+C9LCQjAcWFmd46RdL0LY8RAwcvWPs5VTiYj8gfKIr/EQe2PUx7OeClxe6uWh9uDgZwJz9g
kmULFyCa8i7zwjVJ+N3CbNTSbJEea7ooMHFtMEhoJ24GSdNePbbCJruscSft2ZM1n/6iuj6kHtQe
AGYXQC8fqx7nwXVdPkDZQqKjwOxyWvVSPqoJ79zmBnS+024e6e00lM4PLIsiCoFqdyJgs+BH7KVT
1w/eFgb/jOQhq8dKpjvVwrQBLzVt7Uz2UNw9aUfLZASY6z31sHh4yB/pe6jp1O+cB1157UFrxKn0
yFJH5zogM+nrp+JhCQGzurrK1DYsAofF62rsfgtt5/3elyEGPy969gy+k+PZPX8ktddtIhZjS3Oy
zNHh5NUHqQ/xg9W+PjRK8d1nGQPqwukWoDEm3/ryQ0JmQ94o8tzVVi5qchXKO4cDWtA75DxCn4co
aNUK5ll9+9oAriW+tYJosB9wsVvQ58+HE5s5cGbkU+3aWQ1ZFiy0j62NxunDa1FkXHWJ0HzQwcey
DfGnjVeeN26DMIUyYTw3PcpfJQzwA+dd0ympwmCcpktJbmTwwO+xowa1q4wlU5eyj2vQco/Kh2e9
zYRBz1kqiHN9/IFp5DbJ3RGdyH3w5R50x8u88QIpaPYpG1PLJ5DeetwPRtxJVkEnAUETFx3kAfwm
G+TcrqSbM6UBpHYuOOnmj5nODa8xVOAMARaAfa3GU6+Uy/l4DhcjLxlQSVdZmZaOj4XC5wmtLvWS
gfaIOxNXz8oB4lMxNOXKNd+yEqc8TOLU5w3+Mpk47Rtj/DcLf57yolLEA6m/u4WNVNJnqGvLiGBO
L+vwfx9U32DKTghcsLPyqa6n5s5SGEF876529+phLHGox4Y19Qi0AAHA2asuAMvDAm4ZqKBdEA4j
rhPZ+vYi8UZqZ58Xqo0qyMOuZV/b9j8KlH+nnrNSUL4mzW+yzULL3fzPQg/32dmefIcYaHkM5B9u
RhGZOzh4yZRU6kHlv327GPFqP7eLWvH5mq/DZBFLdZCcH30wA9sCnW0Ag0uHK4smj9UKoHkBNU3L
TkisrLCihLFjWZPdYVl7w2loQt63egb3gMpBu2AsH8n7yxFtHdilPF8CuUUgJPIcdGm0r5XLfGV6
SmUTzrCIbBV8v5oN6N1OqDOlgd2JGhPbjYKxI+qBwwV8G/UHuFA7AC1KGG6kEmYKhVEUEBehEBN2
5Ux+vifsVaoB6EloSsyfivXHgikY6NnVMiidh9ym4x5n+ZJ3ZAKQ+j4tlGCS43Hv3SF8c/o2UyGN
iwbpVOf9jTuNMgDKPeRWTrDvwIYy0lA+/F2J87XUful6///oXZ1VcJSoj4y9ARcVbOT/lw3jvYyP
yT2juH1CDXaPSUVWasrtrl8YRzHiqdw/qy147GnmLwDwugWu8dSrmwgHSQ4hi2TLw73VmqWslTOs
nRBpxPeRc6G+YQmMsznq+5m/EoFbQgciZwDz31jV1JlpjbXR/EJHi8DLE/rh8rPsn+L/iIzvBVo5
3GaGiD2BU5Mo9ZAmOwaLSjug1HsCX/Q6Mx8FwXAdCBrsm7eFLNVPbVTPSxK3Z+g25Eig3WAO2IUf
yIwh7LYJDj5PLBnKvPFiYMWKPMswea3EsiPPNfic6gpAtSEngxLyeyAoZTDvTMQkT+nItTtWXEJC
5CkF5Q6UCFdwsUiDUvvP/UyGJuiZrBFBcetDqcFuYsLWcJU2nuNdLDGyGJpvFSJfXHoBPbGFEEAN
MwA3mAebrkMlvO8fFPY+oZ7id+m2T/cXx/+723qn5KD6WHIZLRoLGEZfQvMlqeXha2mK7bNFrpKV
uI5tvsKEE+i1tSj3a/O2+2NvPZ+bnzIv8XUGDFoiJDbSqU48Vynm/wruupNKd026lgoBeCdzCX3K
gVSt2swT5W0QF92HA4R9uym6bc4kQjzjWfupyqE/C9cFdzKLwveLg0Wz4yqjYVtYJSfpDnVXkpkF
ZpvRnNXY1zY6g+hQ2vGjascsa6+srEOyHQYaC26N3xekrT0lN5HrWmw4TzPa681aS9ISrvx41BY8
GIAVLiRYirOn2BulIj7SehOZBGnJIsP79kYYMbnV5lYYYJYnbeICZpWkliqorT//ainWBK3xe6zS
mBo+7jXGIERes9OOLk7/+2JitbgizqbfAi18UmRUfckGSmcEc4A5BVgn89xnTKaiUjd9Hz3XU42E
zl4tjAK0W+tZogvhtnktP8Pw5CccwTT4NVcj046Mby6zjwaj/4OC/bGGaHtX34d+VPu/9BCLH2B/
SprGDPnTA3Hk3ihQuPD8ctvy1f8YKRWGgChqalXagl+03u5gyWZ3oEPAu5KGQmBPPFC7BB/rU03z
IKSlexw/GKpNi+ulAOjuI+96qFdjJKf0RzoqKScviSvY3fHf3JoH+1CGX5LO1FtkL9Lr0m0EuQqf
IyuM6K1cmAc2ZKwwRsWFFfPsNJA8KMIvL9CO3aN7uplYEMPdRiVQ3xbLWftxudML3nqV3bK5OVLK
QaxpZJYyrcC+W1U6s3RRRwKxKCnd2uhSc0Y+uAZo4cuCygDZ64OaADIyaFyM8jQ/OUmWIG+8Ji04
GrVx822XkLUTrSOrbb4ifEfr2GzJxTZkxPMd314MFcLf1bk1BbqlhxVOohWckqaSkkQsViJ+maTb
zD3lPE3YttGiRa85EhSPB5BuRa6cjxkIan/lkIiATSwcc6+oHI2EoxCs5AnMwHstivek9Pr8dCgk
aCqKwsGxCwPm8FtTBXhgWZfUdGe1kS+nv06yZlHjtwWdWqmsx7ZZeP3Qi4+TLYLKNEn+AAn16mBX
akSNkHHU60sy6HfbRmvwmuvHm/527NsDWuhVDO9iwioOmNSlh+/AltYagup2zsPD5oZVlfONKovx
oEvzl5F6fkbpB9ECSSCh237PJ4ODG+hj5O1R5rmiGERczR0XT3Qu84hI7ql37YTntpbt6c/MtF/2
2mTPcZd2bXjqTLkEMUAZWW87W2QJ4iKAro59NcRctFGS8pCfESsAyS8EyrkAcKKN3Yrnp8HF+QCO
YrQCAMnplQdt2esVlNBBwBB0vxBEU7T+i2wkzVzwvs+zW/gh73+m6VYLh0TU4egdKmTeB0u6x9Kf
KtX8HXPBqcqYT5t5bUyCsalR6kFxH3VvL1h2KJ6EpfaA+TJfSDRaOVnN2uUYP/acSCPHFKMyppjm
/eeaHhuZkrIvN8/f4fj5e8Z9TjoSyT8hDO3WaLmg6UfOLKYLOb1XdG/iZ7rnQ0dyXB0S8q4i2td8
KlW+5BeJNgIRMw08f1Mn2dfb74WY4Z1LDWEIHaGIdL3kQHeqOzo7v/2zr7/qFyHG5nzxE2rg1xB3
TC2ul3bVPoJ2/JRnac6eZR+ovquwEWCcvha2EApAHRmQ9MfK5yeWzRSTyEYVKkHZ59YddpImxigc
Q+291thZZ9lJRv/KI4cawVP924Y0tNeYcDd1ydtFsNTAzN4TL5zFMfWFwQZn6T+/WVuUOTeWQkoe
hhijI8qzBGdOR/6J8WGoudT9UXC689tQG6a2wi7Qr/QYa4/eS9uG/9lrvkSNuJhylMKITQsu3Vvy
kviQt0YOroEpE7fA3gw1TMU24NxBFQW5naaAZH9vKx0sFqFkl20g9W990BxHM4gnCRazxwciMG2L
A10j1adfnjEJ1eC+/0fMi2nUzj169JwQAM0xVGWCwSGwAigprfFpX8iHioxKvmymwr0TkPT2CNjk
ekWToQdxHzJGYddglhXp0sMjMDy3UYhAJIXJMj5IdagWUrea9GKbXxwk1blgKdjTdTPJbgVC1ouB
mzHqrqbbIslwPYGkR7LWeckQ1rXcriJ2JY0jMSAT2QPestLSLD6K73dMFOnv5qMOfWx1lz+GYFte
Y/5HvetRvJdVmLmFLV7dm8l7yUDDmlybZEWqE+RNyXc94W0IoqtZGsvsTVBsgQixaIfb4ucfGfGy
MFIsK5DZRprqfzHXCFNH5o/Ff789AIwD1VqGiXYWjHUdvBl2pbE7FVFEZOUuXEUguyHdBkM0oI4v
SxGJaeQyoT7+rZ155imqNjkEmbFKKBV9Chm1dbSqA/TQ28tTmDOAjASd9CuInQsciktNat0UpVmq
TRu48joPlM6IiejF124eS15MDgQlw8JPxkA2m4xzdk22yX1YAcB1K7CgyRxqjF8KNEErxEe3TJAX
T/4+fF6e8I2YzFzjSfyafAXj3CfDeVs69QSOPuCo9CYz+kazOE88zpwueWwspczI5ZZ27+6jwDAu
6vbZ+dDKY6omsu0gmYSt2Pqjf2HRtLGh+Nc2ns5apSsaO/eeCmTGKmb/LFHoEXaQVZ+TMBGCYoqQ
MsXzkw0GHVZWct+OcyRTKqI62RKSDQK8OLPxi6lLKNTj/BXwchmG3VcHTrc+CB64fkW4tyzzQjIP
AeoMwFjvdF0uobH4/D0M+96OC3k8+86R3UJitoJh/NBI7sAm5iTIy/wUHYp3uvrs59ENbqzfpp6b
/tF/KLEnHvG4IPDXN6uzbVh2T+lMLcqi7xVDY/OspwkLFpm095DElZhhQ4fePzAu2Oza1kJ1aS7I
ZPjoXxRWaOBC8tpvR4DKSESsTfC7lEAu/1BzFXy6NZlurzh0+RgtPAcCY1Muk9HKX8AhYyQIn5F4
VuwUXQ+bZLDuYDZI+JeC0J7yblKTPwbCCqDTK9VrOjomCT6yj8SsfXFZFCGu0vjFsFw07qBvCulf
tzn29Zb9EojF7oKxlltQRY92sofvsnEIKVLekGJ/unI2cVr6+9pY6OYYPgxASWmB3ygjDANAjTBn
kcmI6dQpciboUuA9WWI0wH31AbdK6xql6eqM/NvzkEi4ymL/WDTTHRujZbOpbbs29c7SL88FUKZB
hAWGOQG6arOsajcX1l/AdxfaboJnNIQXLT8gxJIePxmaDVljwqX39efoiU2O3JCFobwWyyXthjuc
BGYfovX0CuZwAT9u+d9P3iquBlippSNHUi5b9WfX9Qrdwe0G5+kEunEK5m3sa3lWnhNrTs4hNjra
oetSuebK0azo82PvOA6PbknoVUnB4oLHeAMH1GyFo4a7HCPMQX9mmx1kF3HtlK8ZD3OvRXXAD7WY
PPbvoXO0fZlOJhfFp9Oz9L6yD2MRSyQoYckEsL+FZJeJdFcDBLJ/uVPeN/8TVIaRQH8NzGCVBOD3
cWgyWcFP6nHElrWnTLOIg/cSKseA71WynRaUHM+qTzMplk3xg237+G7w35dHvq18/1b0gUAXOnFm
ttih54nnap49o172l43uo/PKAasWepJ4zH0fuSZcCKwQYqQFT5UofNmWgGSbkrvDW5uBwP1R9Q+c
mrUjKqw5gmEt3xVPcFcWyzXOP74+a5X5NjgkekGF9lZHcKn3Vt8CqUVJx8gVOpiAAADg+IlvrdY/
Qljl9sEmmHAoLtgVDI2loEevV4+P82o09vkOhIMQJi/F7ZgrCsw3uVZbOIub98KMNoIPRsmHU6n/
KkAq1FAxtuY4TIk6204tHvyzp86rMo1naYDaynaQpQS34c8eyayewgKaNxDFNHftqAELePJHbIHV
KamY0zYYWvjARO0YvLwViYo0hGCe12IToiYSxCWM3NukhB1EurAmUl/rq0QUSBC2vxiYCiDgLOBF
eYJecEId/LQH//J+Eahdi9HPh+iokH3BVplL+/MfC4YpfrAKCGUdF4ZT2RAQlaodVieydReiIkYy
i/GuySaJQyj6BogfF1feinteLqTwKBSDtaWGQv0ax6dkK7jVI7GVxHXS1sHFsCN6JhePEaAmLodV
1M8YNsJrKDYBZj0c78oAtrAnfZSBdCmzxYhw2Bje21wdjN5aJQBlqphQdYjbvR1Okw5KM8sCZZ7F
jVBFGCDZyU+VGdqka4dj0/e0LGowVmKL/gMWHux3rGNU6BuwBrA3x9cG6hnieaQZpYMEqMuSk0PW
pqKXU2UryaQluTQP9szW9tEzYCTdcYY5TyzmhIyIHqaYzKikqJFQPKoYDcuha4B9t3BjyW4GS873
aPaUp/CofOdCLLwj9egYVO9ecYOGowcYw7J4THHfiJrReJTNtMMvTqlAu/El3f3aTdNKz9kEd682
JAWhprpNjC+O3OPD4T4ZBRwPDEecwDxkVW5e2JxK8uVjazg50fQE9M3xmIiPkOeUoNR9nFYK34g6
WcN5YH9/q0qcBp8yo0ixN98xytP4YLwOgqy+v4h98GYooMM6A9JGMy1DBxdq4/9iLHQyJSc9M36k
aiKmilbkZeArMBrKGy+7pLeVcKaiPv9mlWpJV3TI/mzZwqDCmz/rUZjY9Im7u3poyNrfz1jkzHsd
gLLVBZ7lD8zvU2/Ku0pfBZ2Iy6u6o371dHnGsQEMA9A0Ccn60+o0iuyK/9lOoZq6ZwVXrGhkgtbs
lKGz/N6ZLk2HXk9loQU8vvwRfqmXKcpwlq9hwkup71xoyPb/6c/zzpdrwkHuoLTnhRAJ2Izrkcek
UFbUnrz3XFworoYWQ1TXyGuukEl6B45W9tOd1SCkz27Nj1J6yIzSURn/1g7mN64a1OWMEWaYfA/T
Rp5hj1mcQ+w8/FFwzVk/gWO6K9c8zZ28JdwtC85d32hHitFWGbBQ6c3764DZiuiW2F4oVGld6Zdb
bnGl+LVH6jHz5/0M1zhVzlHSRaDd9SIM3Z0ywcUwwnbzH8o5Pmned3o5ztQauQaCwCkfy8mqxrfG
kypQgkHk+We4PNJOb9kVRr7H+6gcj0UhPj3pTPVw0dS5T7jli0QR1B6WpSdo5faJ7f5uB64+boLX
BQAqFkLcxL3hgPFpMTkfIQfMfUYQEQptryM3rYKizcUOZcoVRxhx+ESxvqr9HUFf/j21G3ljfovU
1F1s4e70X9UpfJkJM6Xxj+y0GfXyNZ9snEdVbNc/pbvjTq1OJZ9jWpfoFXfeRVznROeYCJUic7rH
ONtB5Kg+NXCodgQs4dlLlhXN0aLiNGxhoeuWvBr6lmT1k+yVB8vKHkRfYDsp3hUMvVlxrCZY4e5b
Iemya7mGVUCr0bkkrD3SDZL2dv+fOlG/gmyIZ0cLjL5d9yvFJTcRa5fE7wJQCJN8i2IoCpijEBk2
nkDA8j6ZpN2geQ/19deQoObTiIZGzsboRA0pTsF4xcqVM55nZOEA6WjolPfuNtnIrW0e62IMSp0R
MduE0WqCTlnZsQkn9mBSFIPyUCbI9MUI3ccIac3VySTtxKjNUQuaj46BzgssLuJc8yfASVd1vtnP
1n8dB+2Y18cz/Udgql/o/MrdIh3eCFj7poM7qksPXCMx199bvFAggayYkvQ54wLGtMkZuz2MMwtk
CasL/KbGJTgqjl/WKziqNXV9a9dOQsnwPzf2l9OFjuLKrLVxmSNcE+4+cLEBiAv7oF7aq8ly1Ry6
PKckr9i/iqToYz4GTPmwV3lOgeJRB08yU0xdaVJRHuZZeGbqL/tOWsabDKw0Waui82LtHN2FCFFN
0zsCEdCsUnHjXIsvwnmjw1dOMTNVSZ0cQSaLkNR14UutlxAs6ikRrAMws8H4eYIUVUQPO0gCYwbs
0dZKds3xzAmht12h6WZfZ2+JK5CYbcPdean0eehZhIEB188sCW9WmzCPkygz2R+2Bw7haFHJl21K
CNMZxGurJ5uccgBAFcVX/s0hbfMN3Ohy1cbsD8cUh9DTmNl+7ut5H/bQJnfRCpNfNgedQSi6ATZS
FMg0y3UNYZr6UsD1zU3cLLbS1scolVW9SIdaKI4sejuD+C17kyB3cIgV/netlqttU6syeeAzwMR3
AMx/YlHyE1oqdCRC9jYPmLjC4s2or+Q/juMYwhCFngaF/QbA+NpGfzYLwuu8J3+xsxJY8VHiq72M
W6IWDt4W2QrIadNYSY59+0LdXq5JFY/iNFTOtmbsOzbVHXNTVC2kx5q/FbGMZSlFWX0Bs0mX9fyg
rVhzD7xylWrl424wXquhuvQY1muBkcwS3vCLJri9HlDXX2k9dn0ERiW82cB19QJJH2eRrWJEHa+8
76Vs4lvefLGYnu6XiFAFLetjobIJgogllfBekCmR4rrnEx+Mq84NPylD/DZOZF5V1oFFJrWMRr2w
KKOCDjLIIcNZTIIH9MK5iI6t4SFqc6fQTDFQijb2Pu+rmHNsmAoeRtCt2DPTiyTpiNqN77vAU3LW
bruWJOjpPSRmAxUTk1sRSf4oSbc6E2AF0J4iglPDudkKEW5j1JOqu7yfKpTPTyV1TrSaqspqBn1Z
hHlEZW8KZanExp4747sELU7k0QlxshLHGmiI1BSeorRks/KGmayf8jCLifmM8EGSWpnUSCBkkLZy
TS6KJLoPFnKeaPxBJ8ZvReUAu77HgWNK+9Pdk0XgjF+6xJW0nBXrPojnYvR0N4Q0vuuHA9boPPDK
JPzHOUBreszxE7wQ2qniPfPbs+Wks0fJcuuivk/3j3jAmBvz8XRn7JkSkXGhhERYgKKdhZtRPYd0
tC/W0AOz5ijaZ77Usp9avk5igalaRPBRR82Fydq+bLg2puwD7+0S3jsmh/gN3OzhCrVZUvXrma8R
hvDngf3LJy/RkJCkVWoNn3V7vujuWQAHJzKcQPwrqEKkjJXu5g59gGUYAjsT+y5AJsz/CrDq8lK+
3FnfXxE1bUkfADmF93jbS4IV1X2bqyJqRnDz5VvpZgNoYmtoLMF2K0eVakvpXTe5Z82gpAXn9fgG
4ZZfG3uQJVNM0HaqRT+gqkbalwFjbak1obQrBgy+PBMxRuTaCGGhs1POVx36iEbzUTU2CNDNMeHz
2fqhXrDpsdNZSd1D5RJ9FcqEj/WJR7XK2wS5gSmsXUeKvNhbI5kQg7b/odpkaqVtkmkkTbLeOiQK
Xn2hlzY/yrWJK3/3PHdqByCRbxriP7mUQNMC3NuqYFV2DXc/pAqCn17fMamSkzVA+kyfKu0ZwEQn
UV5lf0xCy5dgy3NxYvuKTXFTuvL8eAPnszRNl3PnmJPVgPb25MQoQR+/jlP/mIiU7ji5mOufJNZ2
TzZNgeb6wtqRyivDDhJ1V8NJ9XrzBfR2zxWNMCJnB+Ph7Fv+8rCXfYVx7JXvnxds8Kevb0P7rFrj
HTcz5rWrmP3lv8EKwpILUsN8K83RsnzL1OVf0tudd0VUAt+9tPPaOKr2+OUZA93rYS2XP+wS0Fxs
gpE+QwV6jmL7wTrooProfCtPW04GAsdWYhSfTWuy2BqDW7dTXam9MgXw3DoQSWZIFHKtpZSXTWvc
KoOi9sb9FaYQVohPDVsXN0eEEZ2EN72xFCq1vy9PqHm7RurmQc2WoQgHhgZ0lzr2ADou+CNbtNyh
3YsMxrdDlUt0mPdAH18efikO0FdRaEb767s8K/RCL1Y4Rb9+BV+gUnrui7m1L2OAz8ZOMJbufLZb
z49RRrG14iy/y0tnCiYIjk+gUo1QmWBjl9K19gRCAWnTTAfKDhBcLCFfTTvypPZpUQsIfRpjaMe+
GFzc4zF3+wBDjce/1st02Hfqg4JS0wU6CUh9aitOzFeE4zMuz+jLXsHU5xpEWFCdhmN9OhW3S2oz
xzGewIdBVM1hSLSXV4gYXXS9roTr+xbqLA2Q72Y17IoB4aaanb3gFfm50Uw44Pn7A0PCErtTfH+5
Flq3oUQ4aQ6K73aA3fUakRL2fxjXlhxaJXWabbVnJyDM52XEY/VlpNOIDrcyRRp7HLRzU3khG5bB
GRiKNQKUYXfW1riNqAi2xrfQ8wg4kTsqtzTmgNyxerprC7G8C6jpq9CEQRD5YaXNzXtRJvdYDHcx
CpH6bTD3UJi/cx8dUNp+GoyfUbHDC5ZKrTF57/XcucR2qCA5+JK2TTE6fv+yCxEA1LQrBoI+MfAF
EAzTP3+6O2Ln3rfPeyUYIB2nr1m/LQyimDcyewi0+iHZxYpAW3LhHqSNBJPr3BnZ7ww1pGbXL5wp
/UrkfbI4fAEjiCS9OgOFRkbC7gf0+r+L9xh5/mL3YpK1xVE3tUoW896duV0ugVJbmrlQ1Z4fOmbG
+7L+RsQsFhJRs1EoFG/ziQvCrbbxhsy6Gy9fENo59dUkJltCKJH7fp9pU4aHNEzR8JB7yfoOp7wD
aX+BTNKMn74t2uDdCKgevBljQul5TYYr9QM/utPO6ENIP8WEyJLsxIdfR1gv4PvGwekghVw+J0Tm
oDdeh4LhsP4z14S5fW/ny9QSMRMhVh9Esswt/kSEqzs37WssM4FObunUnTH2V+1hxm+Rpf2RXfxL
jGCIGe1WZ42/ZugBlLxNp1jr/L5tl6sLxWZfBTbwFNzXSBgFwl9ohbMYFRpFcK8v09HN5NuByuvA
VeBv/jCx5fP9gHFwyNmRbrsWGAwP81QBfNACeLEbsJGxsnXYXhcAzAfB8ysij+o9MpB0cORNdBOQ
ydUBMZtQqusl4S5a3XiupFcNdg8/Ymnqlo5Loq6SgZCug3gOvJ3NkbgrHix7SWuAFHSSa6YkaNKy
qdLt1dfet7irpyYM8Mz3J9SleMNW05PeKjy7XKec73QiJWkUrVi++sTZty4feIeM4NCEakNADjTk
ThwJFXUZ8Vnk4nqOVkCFVqEGS0X7HZ8eCxuxJOxsdAE4fGury/ebqvJBqPDcA0lLi3pimw8Og9aS
prjMFJ3CRae9P/0Qc+ikeShTP3CFqr3gSgHVFkIYKHq8RHhNzZihzHamhbrzSp5xoMVYANWsny99
Picp4mJwjjr/0YO4EtesQ0NgBmFw1nlc25zcEeEMMed7sWA129eV7MfkZm+xEo1Q1MnoP2kwkqVC
OnGfbGKV49CFMF8JYN09eVtwL4dsHBCZr40Rn45bC76fMzeI101RctuvFeDnm/kClQ/Zqku8O2iL
8eR9cSdTOtxF7IJUpNflm7ejiXQ781zqmBGjDGEPwvQzy3bE8E51Lrb3Tx3RpMV8loxx3rlUd+zB
Tjg9uPmMfpXQcE6xF11qGtAD6J5XWIXVj9Kz0+AR59fUyoh2BeJkNqsTRGZwVswdq9/pKoylmXRj
6nUYyRtiVXAYN4nYVxFh9rbTjbSoTxHuAYW1A9XeHXoMdqoNOwC1AKy+rwvMgX1tmJhHwiIk8TJU
kh3vXr9zmw+qCioz6yJPdjofGfyRjz0Ok6xFmDWi0V2ikvrvUPW+ugwx5rm9zFCOsJDxByk0zom/
xwNH6kr3Pij6DsRUf6C7yaOA/X3efCMqYu1//80ygWvk+WnFGXmZb3jeGZx3dBJ1SXfFT3t9txh2
tzJJqrdMTGUO4gnSnd5Uu7uBpp6Xrxzo3DOmtr1IA5dTPFpXQbFPtRVjySEz0cei9QrkLf1dewaL
+5VXDIE91cmoCAv+q+rkOuXn/2Kv+LNteNqbyZdEvUt+3oj6WPZ+veo+COKyQwc382sAB2+If2xj
j4L0FChVCbvgMQoVjRQEMvFD5wjdMcdVCNV6TUvneanbESvadV4WqWkGGyB357I5aVy1dM3nq+S/
l9AqpA/mUTCCM37wSf6MLfg46kO80rqotFANMU4GF0P6JpN7a2YK9XlLH2+yndX+9ErqfsoSYScX
3O07gpODlihGksBJ2NVNvbNH5rOYLyh3LRf4PKdjbMFSbWmTuLnJrsEqoHmz3V14MCLE2/tsDJXc
EHsLTtnwLLMUEaEwpYcqoX8hoDplfTCUieVHaWlwUZc2itQ/z8WKSdWPU1FzuVkKGTu0FCLY53bY
yBWjho9+pdkP0+6zaR/eLCV1ig7WUnj4dhNGNspS9IIJBtjCbYErCgsbSdTqiawNt4k66AkY1cl6
SF0zQOfwBY6K+oVHRrgij/QOZlQW+B/c6VfgHOdQSwhgNBoUxqKvgMm7IJPu/A+sJlHQSXulsRL0
lUoFSPQ7BFYNerCFd8vZTKZv+R+e1rcnJfyRoSu0OmSCqFS3X5YMSxo0HBPVmzuIVLAgizTij073
gGqrIdUyULAAA54LpigehtzzvcKTtVrDqGuJ32Ap0TG/KA4WuoMeQvFyAWuYR3sSi4NDiTucwgsR
EfJt5gc+lqCBEpytuxQ5qo12lH7lzgDV1QhigVVxdboHPkUtA3WXYvtxYpHzhjz+pY6AQTsVTSoV
oXS5FUuK4iXc00PfUL0SGLFD2diqcTk56LJfWBec5gdsER3Zdjwa4P+STnekRe7lIs251uPsA/Mt
NeViwiHdNPkR9yKpoFThClHQles6t8WiSCSV8PVuajlwohG2tlzKvhC7mmvSf6rBQ7h8a+Y3XJdF
s9oGJnfK2z5KuGj301MjaGdaH6nbNBnmvZU76baA3bUoV5i5KzkpFdu/JpJ97mLwVBtw2GIyFsCc
+w4CrOMu4p+WmDrXtJ9QzMhtBfd2MtPOWO9/dTXq0U8ak9s5cVksQiJMDu5A4wpPgKA2ModhegJ4
eN981PIYDoaXGbiKQIpSNlx3xG/DC1h3yAAOcHeS61GGH2TLUZiZqis9Hdhk5heTrgUodNuVPD/e
F8raPDBzF0QhxAVlqTBHpq/by6ut47o7m7mQDj05LOhinWwkD8WrcSoQ1iHYZU/Rv+FcfpeGyU34
4uoa1Auayq3IGSBq133qa9tQpTTQq0K1QY76NkQ10st3I8vFeo/mbo0R7rKk8NXtIYYiXCuywWVN
f7ClfBOyJd8kEnuLSab4JFFIlCLEcCVT9tEcNFSHm4lV7EiQ7bmBE9Kvz58tr68I+9jkVgIWA2Ra
26Pvegx45ep/Q7A48T0irY15Rn8NP4eUFur8CM9p/NzLs8RRu9WJXFi4i3yJKisgulzED7XgbR2c
oLmvLOJ63C8dvAuFA+4IO3rqgzvuNwx7YJkTt1z30Eja1xY5E+u4/ttMshsBwoK4St2Uihz6DeyB
qPn5e+HkpKBAfsHr4eaFkY7ilXoyxmj+yzW7bDA7lQanUgVgUl3vONzvWPY/GwD+o9dVdcjlEBKn
OE4ep77kjK8hiUE23vXj80Uuuz9Ll8qwQPp0Z5yG2H8fSHoAl0m4mU7LQ5q2IDLiRG8g2Kw4Yqi5
Qxbob+fx9WgPt14EoG6dSjDqN3HbJfRQIRXibMUDejU83eyamXQ5/WsLS9f1bQAPhD0kHxGNNQ8B
G3iWr+NCRmiD0SLcgmqc0++z9Vd4I9vnzQrRSgDvv8eNo5tWMZwf0nmbes84SbxpK8enuGfotmXR
2zh9vSKH39JilTexMbNWQ0mQkXB4rIllD2Xtp8D04UgVgXERabrAbYWgv/d+n0ncIVxkm69eHcgR
gy2iM7mhkIZ+HXEIoKJNbJ6/WdXx+E7hUQMzxBNwq5qCNa5sVe5/YHHFkqXw6bvyDK7Mv6ATpSdq
fOTmCup87J4swaokwjgWpk2Fg95tA9jQMHBfFoEFlWtk+TRU/bljmlzO+G97Ott/aHRzZ8OXgF45
qmAw5pKxG6DO8jxmHCAYQwjKzfT4jznPyaauuPa7I3tBQB3d0TNKIBO2fAOPCICYThVrOGHLsVpY
fYo1i/+WmhsS94Z472KIN6N7/RytUeRNS6bj24FOrFugHAmVFFqzLTW7EVamqy317o8Pxre0ITE6
PJtePB1GVs/OVAQeu04LtGyIFoDRaJcSqNs0CTSGq3KpPU3WTT6t6f/MtzQhxdO9ZhIhPCDmmNh7
fIiR072vn1x8l0wiphU8znk4wdMRk1Glu/3mu5F53RKV5U0jbiL6DO1SSRbw76k6HbboM0nLWLZg
XrbhWVrsnACvGeniEgWXyFQX2Se7ffhZZ6qTMOHTf5Z0pyfKtydAwsVZe8EmU4vEYbJ8+ovqoK/i
5/2Dd4lBKFakHTQjjo/cXK0LiLntsYJ0VtCi/FtxeL9U9R+zQ4495QeEM7UajNGzUxbF+xGmG1xg
mWMRXlmNAsrFJJ/TK6iktYHcvdhKpgVUMV3GXVF3KJ11xtUWCHHY4T/bcEEZt6UUBP5tXs0pM9MX
YkexzdP7+cGyfrSIV9VRLwlYe40WCySqKbilPaNX+tSihl+X8WohTzR5Iqw2F7pOUGhWS6PZWN0t
vxojJlVJqclbgi7nV0pmqzEBbk0WCG/Y4jbqyutiuc+eIbGle/WMLCbHsa5et6EHrwkf1/HdbLpp
zq3GaKwXPDybFqcviIygtW5p7dQVZ8+VDeK+dsM2fl8XzzM+KJq3dqPnKKnGqgqgP3uPOYQeNpwA
Qvi+MZZdDvcJamV9RXplWoIzXp+lrREo8Zf/i4VlBihPL5/YysfMJ7S4UBnBn98B2hULkZyWVCPo
4ovUs8N+b12EzZizDa0zIZhfZV/duU4Re5B60RyB79gpBlnAeaFE7RCovb0AFbxJWZO/3x1qm+7h
W1NucYACP+J+YGaMoxDQsgEn0WQz1R1Vjwgjd1lC4BNr8QQdN4uX8t2bDh71/5iJ5MusISu9lwz5
j3ojSSz2nUGk9zVPRLitFFR8HPcCNiJLe8mNuA/n9Mh8Z9jUxFseVeEv5QSOWRB0aj0DZ6/9wkU8
fZfU50EDBFihdjp7nplSn9PaBt3FnwRBDpuHNOEExrWcJuQFghrHCQeHJNTorD0Z0yN1SSAvl0yA
ll8Tb0Km2543YzWgUb7HaIaj7GIfRh/7UBXqGGs1yWJqBk/v8Rx3vWURgHD/nExzpJdsQXDVflWv
Wr7ATYwK3kuRKZ7AETSWJPtau0dkcOOI0ymmAZPlFFo7p0+2QWh73tUDasn0mR0nLfw3Y1GSYYgE
b10fTAIgLcmW00htHculuWlI/rL1AL4pM2Nd2UQlmBYYje+rhaowk+RoRbRP/XjPmva3tjcXtll9
nQPTxfDGxD3KtmbLPq+pzin0se0nlaUx+3CX8U1S9ylFQrK628Ep7MZbXNMlpLQdYbCFiogxpafC
b7mJFhzgvp7uuTv0JGenumodWU70jMmzCvtplCAOZXF0g/ribf2NRcM2q3YN4Jm3DgUZZxAF9hUA
vJu9RfYq8PkPlthzKuHunLM7aAwHK76r79vmquIyjAo/RmFNUdpsf+a/Q3EN71YjwyUJ5sXE7WDe
KK3vV5EfYUoDHKrUUnvDWTY8wH5CAGqQZUIn8h8pTmQk570ejiEP6ZqHWYf28vefUlW3qMvwtqXu
WsnQm4aum72+4vAB95ewJ+444OAzBE1HwhslmfUWr3DjjAIw+X3h8zdJq7lWmFRPFuh0wY+pSgiu
7s0le5SNWxO4i/rtHCk8w58rCxKbV1qAHJbPCgJ2QMz51RRX9T8Mqdo4lyp8YYdqmnd+b+MhC5lo
Fx3bW2xkssZmPCd1C1dBXTLZZlOgSKZEiSDxIjXfOy590xS0NE0s8ttILiiFlauN7aMETjeYIa2i
JsHvMVMZnn1JMn785Yyr/BKCEG3s6DwhlrwDPXuIr0vx1rK+YxSmGnKSj7iFTDK2YtLdyyAVpC0u
cCjrvHd262WxjeixdycwxwuNkYZQPxdEq/AbMchN50oBMP6VpR9V1f1gyegFJV226svXEaZ2bpVZ
8713qFvzp5C0hh8Wq6bVSg9nYfLSJ39T357ZEZYAE4fsR8znXcAyz7ahXjxUlBA8rN/xMDe4y05m
/ihcH0520tw1cxf00dOfx5cAG3eOs8ZWoyerJryzweN2EC+9tdd/ThNKyy/iq8RLf/Z+Li5StpPW
VBRcRRbMGOorVIBWXKtOtjrKxRcfaAa2wfIR4QraSni++K6XyElCsztKvOeWuz7CqeHVf0vD5Tau
l5cs83HSPMVwYDiSupR4HPFw1EkU6wzPIDZB4iXkOl5rXfubwKk2ukUDKhXwcDv9Om8byCNCCg2T
eF3FDZf1yRmzqjdMF2mh/ZP2StIgun7uzZC9RbMxjZQ10HXwsxyyk7vglq8LxNw9nzvKqc0DWtQt
bV37uShlHLimI5EF7v0cusrmNXpMBDK4oVQ9Nz1jcTcq1Ju7C8eLBht0tizgngMDBxG4VG8xFENR
8kqmqzRRSux4SnG1mnEWTz0qA4kN6UTnBAtAAqh3VyQIUn8ejOQ4yWyeseUB+jpLtOFN0tchtsH+
jaIsseQl31SzV7Vefn6ZJsUsvajlBn5tFykS9uouLME/Pd4djl38dCrAGSu0YZ/N2o8RHdVwr0Mn
JEOqwZc9M+bN5vcB7j5FoaZUiUOhbW+FVxrWGqxNOnZmT4LE+tofjcWRHwU04g6bY1O7bGCfKd1i
bfNsDz+j529iMsU9KG3i3XdK6QX29rfA5jcCP60UQIOdgXl3CHs1EHV5VTkE43yvp3pC/jYQrG8i
SY9aLTzqHU7G42RySAwJrAIPpkkqRL0Ld8FIJHQu+9Es228y3XLpHrsUfGDhQzW8+NZmK0gybakj
Hhu/zftfCPvbhUN8cxAU6AXp8u8oeEZ9dd8n/RIdieDmwGsM6+xKSgthlYcZTKb62sl+boLuYMxp
YgANkEJJwiTxsLeQmwK6Qrg2CfiBII4iaM1darKwH3ShxYKwqPUDumq0ZNAsXkICcL5UrvWtqniJ
i1FyQCYxuGm8AKLSayD0rm+1Pv3EzRfe7AuuADnjhYH0oTcTbWs0v2d39fabeOO6mHCyiuUKKQjJ
kXuzMAtK+LQ9x8eZMkHT3/jbJqVLB31CpqrTmHN6QNP98rK+66IlzQgpYeM+zZbQDlhDkgiKGBZp
lfee7TLiIitWa7AO8csxXLDl5yYjWz9v2ZG1P5yzP0BRJbHVZxWQ3Y1Bb/NvXBoJCkZPHmjtYpGg
pxRkoIVT3hxu/MarEjZhVNxrvRMn7/FBPN9MDewGbV0JoH5P0GoCEc8T3ec7JsbntyYNoHbcysSF
3OSbgEJmGfPdTyBbdAWjUEDDmjkyjLijcXsi3lNTR2fXrhUhoLk+8paBogcdzmwO6rog5edbOoch
z9yGV2XyzxGsyPLgeFgpSxVp9FfQmDuYzsskLrVRQGVzs4bkYX4LNWiGF6FTf6saNdKLjwGUWaie
eesL+mzzsFhymX7O6J32iYmKsUoPC+sxapO0e59ApkrCFklyeCs1crBA6pC4YXyfG9ERmJwHyaNt
VEGFl5Bumj8Cabu+5zjGezttHXFz8JrbjQTxRvFt7xPvo7W+vFXG3MJXvaCLey29iV0LQyXgA2P7
vQt3il49O5khgexRKDw1NQNWV5mpzV8nBmzsJ+QKnwmwnLDmuVtepfWIgCDzQnTJTlIW8uAYf3Ib
MPiAWmzzeZkZhF3Qg2W+kyPkQ+DIxgW9kixtuDAygcObdlop3imnXNcefODBHAZ/kAgli0hwL7Xr
++WZRmKmMSd/PCU4AKQtYYs31g4c0r4+5FIe20zN4FLK7V54+VK9rjadMNSUdfxk2IyqCaL147li
n866FY22BTprEobsRUB1kTD62LJUeKgjl3KkB91dG/JnvMA+MCssnqFZct7YKeu39AZ8LReS6y5q
TAuIgBWX1Nsb/Nv9n3jj8IVez9GpcqAqZE3mf5vvxVQVZ1qn+pQ46U6ylcsr028CHSfPOIMYrKV7
s7wgxbx8hpzi1ZFU79g5xiN1SW4euduXxQYhdhLIrNJSWP2yjYd6BPCS1FWOovn4/B0TdrKMNNRa
78YoYeuW93xj4cQ0HiQarSpwzcvXkKInxP0+l/PjPwgIBrSS+yZau1rEXxKIKyYPyNN06ctUN9gJ
e5BCSGrvZUM9IDUkyditYYYm7dOTNpkZnb7lt9urbaYUX9icvO7ez4YcsiQd1TUujgF7dyKoHorX
78VJJL6Rrph1oyy6+np3MPHMOroGvyorcbzzQMOtm4InaEkVw4jjqlY2hgxcVp+bEAUAT9X6246j
v4fGA6SdoCHjl7BUDssMbcD+255uUqXDhBkdqbyyGWokiHP3UOb6blueueUP7B1QkDId+bHC7w3e
V0/7D8SVnb8UeAnsezyPrLqHsASv5oaf5brkcfcCE1y9tq0+lbjL9IIL+Lr+iG+oXOY1VpSsTV4I
0l8hOP0Imp2n5CzEC6MYC35qgPVM1Zjby10xv6fxBGsiOZV3Sc7nuv2Y/ropaJjp7ZSFJOrnUkPa
bLVHLlX2uR9zf3bABQGbYW3nhRCQkX2eBuz9QdrMdmLEn5K07KreWRytIW8oTXVgOOSGbP4SIUlL
9UoXVgYHsqNv9Wd7Rj6xRpokJsvOUvK85ctA6GTwmB3SbX7Yq1Shw7/eLKlluaYrWenI4WqopZdf
4qH+N8yAoxg4TsoQvIsSaZTayg0kPy42Tqr5Yy+4J8dj5FkBdiTlzHNwkevzYskiGTbxsHhgWtxF
c3sB0hMr1eilWfxXIiYw5qiFmT+1RJzmEuSxqIngVQoBaaAOgPbuYWSW2XLKHoKmyLSXfVA9H+T6
wqNiXaSejhSLSk78kqobGMt5Ez7yrSs5PxNpTREJUKBLmaEEiUa3EbYPHU3igPmCCkexH/AzHjHi
PboXcu6NTN992m4cHxJRqEYrRMrtauIjlfXLs7+D3xqiVGiKe/Ud/geJOQ2WUEO7NjKHcJbbFyn7
4OpGFaHzTuLJqiXmGkUHOhPDXNWUjJI0vBz6MRiHmGVzzwLlrGg+ONCUX0ZdrBnjawdE6Lz/zBPv
sLGHcqYAiNMF91d1gxzZfrHyyGzARhbvIRZI8V0g8dke4+P7yv06FYFgEpCcZuJUAjCXC9nS6c+o
r8erGepmPlxseY00Z+dq0XS8XF1tJeP5xYuyeYtbgOGz39maVJhdfMGm6ylVul0deWw7frKKULI4
FrsCXnAJKgch6tGtASh7HGjqa1T1dmpM0mkefC5Phv2ReCqejwXiWIr3Su4krL2BwHX5u2Mu+bGE
TTpuuLkBuWNv/Gs8NrmEN/YXjTSk1PctUoOCmLqhH82BwIaZSdRyVHtSirjIM3HjPJ+xrdKWc1qm
u0WQnDV2X8gcDjTWJImE3TmGEfVuZzJDUc8iKhpatIyVkKfCVzM5mw0gA6WpK4/bgNWY3VL2TffH
xVYiOiqSfqhQ02s3MJPYNViknBVMth3VtBSa1t7XG8+34eSsbGwtuZmEmjJk2GObMYjSEjwSyh0b
9814QDRFvFQ8jSDjhpj+hVK3BVDXa57KBFlQYVXOg+iAgkLE2bGcpumnCQ1IUQzxcgRrDJCDEE4R
BBIsDP0Ymr7ZySceZDHsJ89fPcrpAEcXKpORjD6GhHsji2dag2wdOXrtl6rvTeUQoEeTx8gn0OxO
AvgXYG+FrMdi01r81SiT0pcwxIlMjDjHMV5zb4OkYzRMQFmiR+vkr6xNBebpRk02BHTsMw8PqgRF
p1yAKBIp6dakdSFARKAwYWk0Ux8qL0IRvTSDbDGNTKBI4rktsOlT1rgj7FdQKny/xng3szWVDIEe
/XcES4pDAjzN1k8BY8Ruk+YIRVYupvCnfLvmtVt2nTgdEwZAaYGTYy7FYFb5Dsc1Mfr153kEsonX
ASh4hEOrcxqMICuvaWdpBw7TmTpe+5LoAHOlhnyf4Y39rbbYJIhTZMUzIr52YFh1az/ZpntGHX83
BnJtQjkYTnWkxWCHWrFny6p8lObRB+HWVpODIK8Y6lQMX13Tc2z5r9JF1XDqjbbnsTUXGmdZgfUG
YagHx9dxsiQ3mafd7MbT2+DrNKYRDz7DSdMKl9KljcOSE3ws8N0sNKFS4URx1jAn1gqBloyzVY+b
EpGp/5wGN/GJ2qGsYpft0JY6lShDdXu9E7lge5Fx+YltlaaXXtcy0kBFEntzhuKbUazVv2iRKUCg
E6DHHUdsMnR0AVS3EnaVcyN711s3YrwrKUw63BPn1ZpEW4796Wy9JcAilBX/pHqCTTi9aGb0/NUf
cXwgyyhsS3HhnUadS+v07t+bSmF+IO2aCxOK+S01U49/ec5BTrN2H5whxshWuTgnwEfSlPTtNokG
taEZmb3s3kZAS3S7CZv65sGW/z/lsbNglXXILuNHDd7ok/9MVkFtZu8Dw861SRAzZ6mkraaDwSyM
0bsLVmOTjnfvYySJJP7X/NkEz3a1eX6iihAHlvmPF/jkRPTbL+DZb6Xp1mNjsaIyKtyX1GOGNG1u
YtN+zhbepMOTi+Z1qCR4Kt3c/fvaPbBmrRf8CmA2w1tfOvC/wA4c44pMTBQRmAzOW20NnAInWSa2
kBb3JZkzDoeUIPHPBAbFSjOcru+IHz/LmfXB21s0jEhNcqbcI1yMIO8cnAij3pZR1zO6U2onev3Q
oGrwa6flCUM+jQbKh7OVjb8Ovf/sligXD4PR/1dsOeT5K5jCqoxEdIcy9xEa2L8n8Ev97nqAEFFG
mE1kT/u7sgQGzJMvhkRtN3xE+V+LJWVJZq8lJr8sapc3cSIvhcb8EXL4lIbgDZbZORpa/LcAQF4u
1LGcRURFe8I6Sxl3RSNOfK5lC7mkctRZ+FOOErNho3T5enOrObjYDVjO1HGJJ7BVCybnWbMC1QEE
K6j6YTkyni5VlVcPRC7rtxcOU/8/SqAm7ybllO00r7qo7oOJ1C1PiKmPDvsRMwpL+D2x+DqkRY+x
B5s5SASh3YaQI6dvp66E4ACItMch31Ba1am0gf8IAkOZYdjVpCeK9xruRHBCjuEeIE2X201uziwz
UuweI40CDea/vUIiKlBIofVWsjBj4NgWL1wolbNu+oAhOOLjFpeBqHYGcTVayZ7HVBHSHDVTMTQc
au4HkW3AKgOSD4rlaRBh9XSU41jcE6BrqrwTIg9x/b/BLQLAOZhud25nncuoF/yj9RIpcpPgIuKR
Hr90sUcYwsHxJUe1P+pMV7kWf7YuPmlzCKzqqyzXVEaHf3l7hDr6HEAhfHGNHXnb6LVbxdsJLcPW
vBfWHaV/3NxVMV9VGzBzMg+w5x68IqpZSO+vo6RF7x2VX8Aj4Cxnk83zsCWjv44VqDNrds5HdaJy
sYoVATEcvUuemDPZyuhL1o1tOBqw6OEuo6NHiHti5KOUILtriw82qfGOgOcpRz8J6iDY2aXrDU9c
Sxz0ubUosbCtY6Rre/uUbFZdz4zeYoR1V0xR7teTpeKdrX3Rh60c5gxEw8oSy69Eb4pVS9Wk3hMe
vMtAtBG8wkHJ6YFq31sZQaxwGC8NGO4RRZ8fnd5K+LjDKHTU+ZEeKp/zosUdh2Tr+FZ8KRWIVtMB
2NYZEPGSnu2/KKW1Qa4tAqDsVEVMI6x8JnmxLLQ3jaZWjpoWc8xdDSGsiOge4NO5Fp+bsLX7BOZH
NT+PTyJnuyJIN6jfYJMfOOOPKxOtN8RouUyfaoX7xfxiGv+8bco26S+D+IL0bXwmbHJouzli0SHL
pPXo5re1I2hHIOyqL9m2NWN4dqYjAW6OxRon94M/3zRUoTR6eSGKus0ndbqcEXC5Q318K/agibho
AszdShGcsfMYooQA5AgnuEh04qj4RCw8/93dUpeXcGNp3Kiys/8ckvEexvqW+UXJ+BqAPJ9QIEYN
TUOICRIBQfGHZQ9Pn8W2q0Mijwyz/CMsbtbur4weHIVjtvDl9WRPKxfG1DNydH7lasRFcP73RI6g
SMz2ZREceeGfF8qbkdcYH3DHpmSllgEHNcMpvBMVt8Wj2f9DMS86uEKdqWCbGOLZ0QvtKxPJ3awV
9g9P8rEnBPGA6Qdmd7RkgcE3kNwJbX0XHouvUN/ofgYorOsgLbhik0LELODv0bBF/jh9H3dSy0Uh
u3ygxGi/VBJmwgS8VQHEvJy/AlOEHCjsK6nvPZmsz9sQ0md5xohhlBKmJM2J2WsFIE28xkmMrI48
F3HwTsW+WN140a5vvkgngxcURJ3/RoRtxGdzmVDdT+XH0RcYydCvA/vdxKJc7P+PiUojC7ABXk73
UoFAWJ2vVRNBGvfhg4okuiD3G3FTwvYg8MzXOJJBYM4fAfXZk22q2AIUuJPv0AWSOjOsxXnpfF3i
U/OsQNrNRQusZ6HUefOl3bZyykRPVcw0Ho2S/U0FqnsKBcgk+wPMUXUPD+k6QOHedi7sovAgHGLd
CsqDa3HSjiA2S79aNBm9Bm++Lwqb8ycn2fwlZKDoX5TMWK2CZEEk2B35hc7AVSENvClnYQvfd+h7
huIvZxNtry/T9u/SFPu9xtHlEAplbePcDALEmQtD7xQp6c+RgCVS1T5VyFCZdN0ZyY/CpjugHmu7
F+gHoP8vZzHWRT/hp8gd5L97fC9Chsf23PtRAgnEjeDMupV30ER8oWF3gEjUiJoMtePTn0Z6YJam
QnGiVpD0UOCdCri3OYjY9vf/l1t8AoXY7dc3sWgv2XtgqALBQBS5huQ36z8gS5j7Elt7D9Hr1kBw
eVO+WNQdaNFG2kYQ+VIfxwVtsCVJZdoM7oC2545dV4YOMvc8pC3sJU9OU/EcOE3YHCQGAhVgTq1a
8l8rW55kcK3n66zh7eXUG53K8uh6EiMnCruKbYqt1LXjiRJrzItCARDU0TpUdvcyIFWZCPTOb7Wc
nGCuNqLvXCLiAd7xrMOuLIbfZbun91vZ7xMy+tv6NRkfGJN5iYg1cnB+iK5aoB5onLhmsZP+k/gt
vCqSnnOreEsoS9PbfhqKyQ/ZCxAWRGDiYPxxvRk3XsQupN5JGNteJfWMQWXXgniIUwiKyrqQuPad
ZGLVSbWPI8H5cjiHhNPiiE+n8dBpaY6ygE/hBbL4rB8lA7OXW1Lniwp5C9WQ1tLIwUSK97k4mQ3E
tYrB+hIFPVKKlJo3JE7aUpxHttYmrchh+wj+f+zpY8Sp1bVjO1DRkOjb3BidX9HNAoAtL4qil35v
IpxzUGuyubiJR43Cy4ViFjBwRESfBfeOvbM/yiyp5EpzU79Sr3A+AdZZsAmc/aREyZlP40gdpqZx
7bHYCEQV4Fv6KL7iWjjuhDE1N0DMxqZGCBS+AxWOr4K9gDvnghDLlLm50zaZ9bTjgRjCaxtMccqm
26bE3nJDYN6NsK4qI9oq9X41hE53112yNKUcI/rs+ziApTPyUbToi5D9TH3agcRU/p55yLzs6XFS
MCFraqCx/jbp30IGtV1G6vlDlRtCOPljmwX2jl870MvSF/Vo20fBMrRi6jX5dqU0lUOf0slPTn4D
u9GfyY0/20qMWeusVvcSJ7Xh19e5DlFONVVWV3nAJX2jyv2AKeN+qVTBWBHSFmKtTO33dqhOcisq
LiAngqQy4xTnz5UhDKgo2mWqyHuopB3xQcw2y/f8cUldXJSo4X1Y+7940gCcBRbR2szWMcAYWHfO
Izv6Cbh9f3FAtW3C+d8auoqwVVm9GCuopKkWkTRaovL+eiPhijReOlDclUDKxnI3eA1d+tB2EUkQ
jMRvShS48HHRKFIBJdDV8NzqfrVHTi1jFWzv1l9HKsHiUSGXRQGm3XPnJ0qGqlEiVLv+Bq5Ffiig
osgUPCKoVYNipNWLSJFogknrP65KGEy0Enz2RmAMgBqVLA/SjVXu0NhNC1yOjJCDFTUAkrTrm+7n
ThRPTQTbrPFEqnlIPFPRWMqKrnjwwHKEYP9suaWQMRHBnL2rKAJm6OCFNgYSNSdhhA0GhxjP9Xwy
a1LcE6wPAdMT5sar+EaRZ6J2Wlbl4Gk0XoES4t0oaP5197FWf0lyE4gIRhE+e3E6JtgWJZ1w4Neb
3Ra+2Z7UZxpL1uBP2gLnNw7FsEvsxsH4zThB2JlHKXNethQ9Q4Uy2nrzkmtgmNWj3Jfb8IfKdcPE
9MqF95ZqB9p/Blm7RnaWmCQ9DZTdwW2puy/tzejVukPaUf6MPCzqlB3sAGqRV6YSZVzyyLnYfojq
6pXoSrgu2xx4tkSlzKlYRyRinYq5ulvkDS0SmN96zE1aOEprkck5kLWqpMOAQewyFAkzgdIy9puH
/IaSJhSafS6h5+0BbQZX3LSy6LmLfSjCMEX15HzipPW14UwJEoG4iiz4zH05631APtsYxQSLAmJI
mRnNz0iVWlPKJvlKppemEu2jS96EuAqfpQfp58oOIIcRF3Pfi1VrN2gsrXAa4179teyu1yj8Xfza
+RQJZ+LYbA7wV3Dn7cQuyls94VIY56lyJneCYCSXk5zVIQnY4j3xchRrJd5wyuZVY1ildBjHKbki
qxjEeErA3wcqcWv9VfeC0+WYW3Xe05Xepb+U0XW591B6k18WG5yHynlhfFXxc8oitpe/A9ycJ9gq
DUuIaSJyugdM9Rpz7e0oLPwYaNTVgiV/jqDUelBHWaJ+/TOMNHZrN6lY6P3ylMCaezwXW8Xg8JCf
YMLzwrmrxvtPrkrafQL9WpJDtmlVIakQSzpspVMEMicFulHqySlyvPRrYfEXvvPxBa2g5ldfJSI4
uTd3SOc3E5pwTmEDGLIxc/or0vwvmNJVPc8OcKvOiFr8D+WPWLQAbSt28x+AefwGb0q5pl+Ha1B/
igS5kEICQOZhez/iJM/Gb+4T19cvtaro+l9wL4BkiLOIFvGdKOTlZe/Hk+O9vAuUlI97ZWIhmWRH
5Z2D7JfNP+jYp/oNjTywHXGik3kII+s4HneMCF3NO9jQyebyONQnr8Pki6aI0zlSu4sCpOXVeqnj
6QdO6cPOOgbHPdC3q2zp30VxcycDdc737X5+RXu9occb/7GKf1g9PaQKEpEC6h2ZaWvZ3KUfvXF5
GMmla9SelQJK8jJB1AnklG1ouOqLDqbCM5D3qQtw4Vn30UII/C/1h4eGwrR68hmNj1ivZNC+M4pm
+CmOTZNXSSqZVN3xaSUyHG1jh/iLOZE1I+BqDMeeTe2cgIXKZ7PhwZt+I6KpSjtzZNvT7jsFYsVZ
YqMjI8BdxItlB9MA6bX+r2AyFY7pJ/mM35MqGeoKLyUPZonMD92CciJnjkSIQAkevnDGe5DfVotC
NY0RUpto/76g+KePR9yLhnXlEHIwSfirFfroNhH9jpcJTgOMuZ37y2aQf7w87Ah3rMidoNyYmQPD
1ubGpSSzpBmx4gLmK6XNXyK3BkXDh5NmqurdR7IcsPQJ9g6FltapPcnNoeDxxB8u3Dlj9vMEIuE1
xlw7XrgZlQunpiWyITW7353IRShccfvO4S+3Ar4tYBMtkXxZNXxBZhWvH4qCdV3ATiNhJKVPq14G
nCc/Sy7G8PTzXayxA6XbPkL8WmmfbiA8X/7sL9zynSIZcoyuGAOvuTOhoc69mw0h3At1eTE6CDHA
qGk+c+0B1R9g0CJ0b9BGH6oHbx0IWxlk1zqqEjUJ8PzHW70uT/xPSh1EEtwIMZCJuCMwylVq2DVD
rHEkKfcqS1eKu7Iy5zKCbvnP6n4BrudS4jaSLxwhcxxgdhUpADxfhuWGGP5Oq2JO9OY7vmvDke3Y
GEfVSyh2vy8NzRA2l8AdQxl0ekpjGN0Yp8AIH3sAerb9POZOhlmHaP7nwXg5Id3odn0aW9e+x2bW
PUk9M/kAgS+hCj5pv4N+4B7bOhTaRDoodzPJqUknyPEE+qtmnq8dpKTMUwrcaIB2KsWSyEksxlgy
yYrrczQy1vThxKeqqzBryak8wQeZ5w9PdaFGDfT8sHoXMoP3LrjDdsssSv95MwuIdd1PRNZWlu6+
gs+FVP3x3uGflnesNy3hh/WpXgdCFJCeJAeuOMTHxsaxHXqjx0U8oEH/KRxuxmK6hf2ejD3cSWau
BoUKb7Yuz/E7/ExnaEq00JKRfL8FekNR9VOTnC+blD5KKwGc0RA+ImnlWled2epMP3qCucglw120
CfI8xrGfdbFmBsYFLIhsWNZvM1JdqjhPbiDbYIOYGVSs6QiPCIaopCTOTrz54hpvfz7/metRgKS1
LIG0QttTqrqj+y/S7bKY8UIWf76/h3AR3bL7t9iS0bwtI87z/6kgJKOsmqQiPcmafvtpLydmUdY0
9auiQHMys9V7Z3jmL8+fzIpOGCO6OBXR5nCB/IWLh40yRWLSS0Ty7jPekSoUIKRQnebkEDOwuwZQ
62ppxvkfjoZSQb9k8UG2kT8gtBqBURVRx1xkar7Qt7UMcqu73kKosKrVXlG9wobE22V3uCNYRrjk
HsymkREPpx327B6a5x9cSj9DiyyOSye15CCOj/Ajtz/qLxrqYGGizOCBlsw818Jiv8nYUX+qXyB9
inw+7H8rTz1gdq8HwwXX2ZvbBlhwRcnZAIgAUJYW+tT3WcvBnpv1jcJXAfM7n6QpUDze1+Ky7Ps5
YfYfeK52IJwBz1t/2cEos7rGSHT/xoLjOe6Xs4YpvZXcImICPgi8Egp/38NIatcEeeonjiytWZch
lnDQ27c7tHCgQNvX81Z/xK36kXNRBT2/WZOQAOIFjzGy851dfOAS4ohcaY0RXZ8WHm1zZAalCWVC
Red/k04SrgOJk2x8zT30wKJhpVRYGfikWfLHlPGfPqMQgxT4pYi67mqY7hVIKLOD8ENPgjqp+P6Y
gpIYwoz8+H6YqPPYr8B9wbijm8yWH2OzJLo6LJL9FWdGhqQtk1r2qvKOStdjYB5C2QPmurBQ7VNH
zpoE+XypJLp37Sn7uQQUC0V5l4G4OAAxBpV/QWyK8lAdIarQIivDf9zXULwwn2qN21LP2fHGzBJn
hj21fHC1I2bsfEu77u8c7NgLJjxhkPBmirwQjZhnQhZYk6CpF/5vc9SlGlDyXVF3Ou2fXyHO8zZn
njT5M8cul6vlcF8yC5BFea47aFS90YGr0mEFSQmr/WcPBR5HotJwAICJV6fzXasA5Fu2OV4nQc1L
O5Ka2c5Wwg4mIM+vsttOnRTnvfCNkHIAKhq907tJsq6EGqKN0fqtwMOn5AzBHK+IlT3BQou8I9+9
4Ghk8YsyDJxgSeWMtv6z4hEpgB/I+yxdpNI7EvfavIwSwBcbe96KZE86AMl5G/r/TlOO10WnlqNE
bsIZXYgwaZJ82iHfpnYdNfm6d0lUoHuTksJWk0//7JjOErd//ANAGTbagXIXNhiqsj0hR2ma5hiO
UIJignC080r+St3e7Rpk5hdBcO/INVHItfuDMO7dL5A+voDGrpB1fZvqNxhU+eiqcZMGsCDXEtuQ
C5MadL/8FSpgvK7kJ7+ubkAu9Gp7Mg0kNChjfaqZD6wuvEvYidmoeZiaqzf/NjDuKJhSRPhLIOCC
xi/i1D3Cp2L8dFqSDyo6mVnhH1zSEQkTUvX6BJhX7O0C0Kj5DyivFC7dZ8NDQk058ONYGWb4O6CC
fcB6hd2YNl7CYuA3xBhtwDUGgHAEXAwpfHWiDWWq91rFLs+iUQAETKDZrHStesrSCR6jAhaLReHM
aSfr2NFtF0lOlnIzkdV0w3Dj7VHYXgrKpvXS9sSjuwtYK917wbFGwYQQE9LfaW3b80LG+dj/aaGx
k0QUL/SNXz2i/tC+3sZGQ+Ky4mdpGGqxZebnRGeGD+x4x/gEbU/U3MmxU2S7NBD8f0r2WpnoxqOZ
DFhqldGWqiklv3dr9AHp1k2RQ1dnXnGXYTmLPx1P98vT8ndFxnflWuriT7wHkP+yOCUTdYef9FDw
v2o6s6wWcAI1r4pCtGAOAsBUiaDjo+pFBeRkF/R+t6BsvHU/L22T4+EGoxmI/EZzOgArmeKx/p3U
zPeiia8LBPdtuVOuVQ8kENx6NvUKl2xMEzz/Wl6cwPjLbvisQRsyTUy3nf8mirpQd+CfictYYEoG
FOlIYTD+xEgeJcaa3WWUusDDWvSVU6eUSPw4KQfuyHELPMEtIObKigF5ElTR4p68Glxw1dBG3Bey
qb4oDezXDajmsvy6O6/2uKHpm7S5Sarpe+ZeSeYjikGMS1vWcHFsIaKcljBSwiYu8uwT71v36XpQ
hj90EOIne58BAHoZd6p1ibQWLtCwdLxyI0I+N5e+gqPcDD3DmqscewCmqSFSBk8yWY+0G3/3hW2E
FTtKUYPPJwy/eow0XOb132mxRtHrCC9dlg9xICFZPzBJQUBwvDRvjmQ1ZB1xOpJACrt1OIN0wTMi
nktRzVylnLZOCKX8f3IJzv25J9obryipPq8YpGeg9dIEJWLqoV42z0adWwshyqM/CCFhyeQFdirs
u11m6ftUplx0pWNDUhlXi/+RDQ7k4zMYzgStj0v2JmAeo1wUuuTMcAcFKZEjfNeNUeYrvpq4wejg
mpc9pQGQDdTlBsc5UtLAKhFl/gWryihgoVs88t9vrY9wh1wZ9RrS0/aBq17ob2rjAizRWID/S4KM
DpBDBQd5ykBVrRqV14VByxejNyUIxueFBzFoYrppkqIiSnpZqL145PLiRAkEl9tXwnzAVVQKCN+O
Rqokru1eUnooz1kw51KaxMoLC++Jg5kzHNlH5jOLe5Il5u92jaZAijJ+KWreThLvK0X6f5OozAnq
8nlqpljtrT1pufDeOFrZKMz6t4Qv4Fvq0ZcseUbU4Ov6xXca6uVVwqcw3/+jw3SS+rjHpVikZjqw
cypGMNEUyUu8NyK/rBAB1eCGhsxxqRn9pXjhvIJFFtrrFE7iM5OMDHQT+swvVM2FVJd5DufFlr5e
drSgDH68zGlah7g0cSoc2px6p6A2hS3GSTDB1gryJ34sqicB9RfDzfjAc5zp2yIMj7q9B4vWVpCk
eWpAybJ13cfTZtWf1Jy9GsJ7gwMZdSfPubyY5GuOc5sDrd3fNGauPU63Sk9MuxcRn6LyJ6H8h/PC
/DFKcb6AUx5vOTlHd9tqcCSXqHNgxAJDY61GX2zA203IGPHM81GhD/M5uPLVkT6bwFo/8n7RmUA9
+DELWNB/RTgToWU0EfeLmFEnJYxVGmx8NqzTVDDpZ7xLaXp347mwNNMPST8eeeZ4W/sOm4cxLMlm
bEy71M+/aJQ/Cab9nW4fFXdp/+8mwzLRXGuWSqcmfag0B6UoJF1EHafn9sQxB+DhDEVIdCkTv0+0
3nBG+8zKVXaa3uR7951L4sU9CoX5KtJEXCmM+a2dBMgEcbf4JKlyBpXURi0xIT8eD9D5wSi9VslG
QIw9FgfQfBsK3O5K1QKAV6tzG2brNcke4xIpLFYCkTpIB1BBnNDNz744Mof8v3LbO25StT8jnLK+
2zqwfQ2XE77ieyUC8nM/PN4pimRbC2jhq70g3EZTf8mdJMurM1sbtH15mkakNhGJrIgKViKPQiyU
1V2nIgU5MiUVNAXbmzbNMeKuu9WEsYJDBS1kx7gnZqy3BwH7lqD18p3wc24QACkWhXaZEihg/GeC
/4EkyKklN5THffRvrbhfpxFYdmW/+3pzfclfCTtFZNLn6ftwfyz24Dwu6I4wcuMhovjwcMU5r3Z+
3CJAF3a7iwzs1xSlLrMAji+Sn32Z4q1VAEckKhfILgTul4w1PSO9ZmkMQliRxZEOPNHkQ7Qpppe9
Nb/qGlgxyy9oiCh6+tEm36iAmc+KqvY30V2SP9qxZiiHROYdyP5X+JqF0M8BoKPwy41cZaiC4JCT
UAWt0ll0+lqHONYoxvV+sWK1wbJ6UEh54/+aq4en7Wua/b3c2qAb4zWQYGdkdiDKhF8Hm1hbqYIo
+PhJ9mYXIapsCq4qVF4PgOX3wdtYxU9gCkHb24fbHUgOD5X1HAIe5j+eIcV+aHcadWWuITyebomd
E+Gc3isEowvMTdnK6yqmzvzzuI8wCB+KRV2zvRFJ1nwdfvXBX90e8KnxWr+TR10Nl0arzlgtfA/n
P/o1MGCagTbV6omOaqw215W4cjSCmc0UFcmEHZ2mKLArgiYbx2Qgme0m22OH+nJikaWkk33GvVtS
pKzPTDDuDE63yYZTwY+Uau4Owt48ogI4mSn3Ntl2scEUQGjUDz3eAY3v6YLlVxF5HsJ+JUVs4VKI
TWJIveDs7RtKa8j0c6rWDlAlR6ez1r2wWJztjZSUsnZ4iFljDZgR3IHSqmPmGP9nbRvKGYeeck6j
Sd5zZKnqiJt41VM6h6J4imRW0Tz1O0os6byiC6tPG5QKlyrknOzxjKR4IwilnNd5+Eup882IBZbL
FNmLFf1yfvughncJJOIzygiicq1X6CIGIxabJHPqwi+vEkHk9GyfMoWzCDtVySpCOfydM79qhbzw
I86cZ62ud0F2rb9KrOSuZ2gA7nk3lDFCOBLf0xtMPpMlTPSC9E2B5oln74/h1R3VNamrvh6xyXIt
0Z6NbF7pHomd1oxO+PM/093M7szfXvvrrwx+xJe3kdsM5c6jJ9DPwKxxuX1QO/Zf8G0DhGZrfAkm
4kv3x04hvKa1eHbWHtptYz6bldq3othJ1YpmKwHWXbNnh8pYjMCYQTECMZ2exhDDO1pOVsPFhP2X
4Gw96JhYeKRIHiXh4SzHMai7GRk789QtPF1qi8/66Q5ilDomepJQwha3eiQfbZHs4tPYNtf8yXEB
XEr6FQfyBYcUe1CZMk0SPg9mwaGwjKMv9ihZzJL9h+BljgEy4RmdBc51066uPRkGV05HZiAHVhq6
vZ9qG6ICpalyqnkCfX2UKAFr1gn+4nn3cqTDEDbyqYjZRBohVwtediyZQylDZELoWQ==
`protect end_protected
