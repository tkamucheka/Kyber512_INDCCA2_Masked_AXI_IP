`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KGg++J83s0yJ7o2/XMVLkRRTRjS0oC9h86tQjl1+xE1m53Uwmm0+K41skiYHo3Urr6lMQ4q2jL5Y
R/1NOu1WGg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jCBx8aLaNWpgdwu0tsffQfmLNKET4Uy44Upxw9AlkO9Ma9Y+tqZHrHroYhGJUxa/dyJZ7Z0HDJ1t
hUhVV6SjuhVMs1NLM1MVw9F3MTSW7MB/qx7j0WAj62FJgoxsCtt6g392p1JAAosX8yACeLKiQ0KF
mnMpugzqSRDI445k7So=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zdO8kU0uCj5Mggk0oLUcYcllNQJVD7vxIj25evesPPwBvXuv6EUsbKmUaCAlFUyG0YQ0mxWxXmzV
V/dRqKxqZ1ZI8+mX4IFaTJSCcYctMZsCl+2EWvQQHakV4QzWuCyca1phNacrRJfur8Ssc/Mhbez3
GLQCRrSfyBYyi3u9J+SAJRcJapyB1syXXhclDtup6m1z2C5S+NX/ql6kVXkcd9P+C5ordunfutgU
6uco8UymF/9QFYiBCWlTkHAgd7DH3dCI1E72N2H/KpX0/0xFBk++NCVuNucOwd9h4/hAyr4L+SI0
6Dzmn6kaBO4lnMAj5P58GIeWO/EtqrPeWg4UJw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FdbUT4bIXyyFULrG0eEn0kqX6tjVoWssNb1FURO5jvyN5IkvkkDKCSLsd4J+2RE35ttJ20+4IZm2
p3H/UGCxkuCYtlZzovVpVf93DlhFUM2iSGd/L3evdLLL8VYETZTScGFdFXqiqe4ggXPHQCSEPD+e
PmMIJTGQka0DD3H+w+9t5Po/+M8b4r1y70l3Py7aYMeCEsZ/yHRmk8szsOjUbwvFEJk8SPXrEERg
EYMIrbryPHXq5E2fCL7hTgHa+bzIdFQOc2/8wn8YMVTmIJCZLBZDXvGSSm16cifWzXKHbPSly8js
RAoD2yYva4rr9cUy8jEyEpUcPGnaJXBDnB7lsQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
eGYl/A3vBqVYodgklvBXVlduDkQKDOe941//b/7D71XaDbW1Cqv7m5eqy+I7bUTyBfnKRV6WeTtg
K2eZlSMADPLNGmIEawb1T81kHA95L4SgxCaMDbzt0t5pO+IQTca0KxjvPFPjj860AZ/Y4IJCgD9Z
vZNfcSeez7bqGB9kVNzxh40hdeBm7XY8a+5R/yPufF2S8KSSaiPSvYwD8yXOBzVoRhqA9q5PWKTd
u6qoeWMnQ1r/hIDsge5oDE06b6+zC7odC460K8KIOtKzeCrfWezkynmD7wBR1fdIwh9FGe2Uq4lO
ZbT2QFx8Ga5NQIwIIZZci/uL4Tw/7+CPKEoddw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
k1GN+kT7KgRIHJs5Cw+hQb7EZrReCsvXgXeCjz4o0RyqpPm8XlxoPCNX4kR8BSaVxBTPm8qGrOj8
IkQcLP4XpLGNjMzOE8knGvgjraCBhhY/bboSihIYbJYXuKW0k/ErxcqbMup3dsmp8N5M+ZYpiEuF
88HraBjchDshDh5xlcY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jzBUDUoUQBD0tzi9B/VXNwpoyjUIKBzxkVyikkxc/QHKpaIlgud+eCQD6psG9RUWZouQN8CQmJEY
0K5qgvfm7GxXMbjLUwnVBRg4Uzfc4OTySfJMu1k9/qGISvYwf4r0rzMMp9aPgp+ElEwTGx3z9N0A
vWNdEjCI2mqdxmP3Q9AYUPTudILppELRMP4SJijczuRIhtAKpxFjTP2gL8zQE0aq1kkWRZfaHW1t
wV7tZ/jCUxkX8uj8DL6Bei6oBC1nTm/FjPhi+htKla8XNUEftaqUre2/0Sxhsxl/FTAzaex9fCj4
AMt2l6o0FpW5JlLhGnTYhWm/bgsyGCPBg6lSjQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967904)
`protect data_block
AYjCjZOGxkX8sIvaj8c8mP6L2C4oBP5/0fUIhhN2eSiP8dQeeJyx6r2X3SbfL8hiKDpCe4bJIUNc
5OicYmz566izAtaghEGQkLHmj07FJT3EEze53GUJjHYibQhPPXhwHI60WKovYjxXjIk0GoY6moMc
nE2lqCde6+UZvWwbm6l/2/OZ1pIZlT/UO0Op7kM86A05r+hu1n/qhtThFCOx9W0vqHTI3f0ZVUlC
dRMkcxE3vxFqscBlez+ENMmtlSIgQyOHN2lh3d7eYaEVmzzPSdvkYJEjkALVxVl5fcfAhIpsgVPw
auGI+/kIhDXfkpZAnEXNgoIpRkDI9SkVo/XiqXVhIk8CD6e7i3EeREcyESrWJ/wUa3Avt14ycwOl
zwjYl85Nap/yk39v9dcGjv51FOe3KGzFBRdchMMO2JN5VpWuMRY5PXZpsola7ech4D+060rmVC12
bAlnSjKsFXQ/cEa+pRyyS5hXHT0q4Eh2zvk7A+kL3nFv4Zi0I2fr4nsh3wcC75hZ1h2M0z8IA4xz
2rFe2uKbzF9uhF4Ts28XaO8Hm8eMiY7FQU/sIdXYJrWLx/c7vQfh5wiCy1Efo0AfJr7d5qDhsrll
KcER5qrHqrT4VzDUNAtoTzB/n1cvHPJsZgh5wBe76qIsBJFw7/X+4cjP+4oh/NQcigAda7pYVVvL
7ZplVK9JeEc+9hGa1f8bZme5FTLplL1hXJFjxgf2EvGhfBwsvnGMDQMYK7hh4vRb1N5SmgVFvMS3
RH7vbaN8Amqy3X4cDE+J08C4RkHDxNtX8ALUZ/fq+zhAUHkf6I98FwEbOAe4nN4YUhiqDBRhoYzD
E3WXKZeG2EqJlrWI/cqTfavy0JVlCWwTlcg2scb38ikX/vH9VcmKWWk35QUxfDQNEjIEqluTUgrS
W5Qy/t5EeMpBAOwRkHDtpPgGk36A18Yut3Qf9/1Lr4O00k/ElRWKy7DwFC+kifJu7dbK8Ba6lyrM
P7w0rfUYqdLSnPAZ6OaIpj/z5mafJSvKcwTy56J1SX+exwDpq/cPPO3cqt3qwVMN6Zn4xMHSjHDm
e3m9aeHV7HyGK1OLmO/Ny8QWG8WAOjs2w86RLQTr9NFsjPudKSgSoe5q2k9vGTKKrni8p/ecsR+z
igRUE6/5zCWpb0XLjwhcS62u/LZ1fdHb/VKqlW00mXC7kVwa8WVCPs6sgOehQfJQKAvJ7WtMTkXp
s7azbnMGMuTqyZX8+n1MzwqKLWo8taTgcrrDVNyI2FCBWdZubrG4jDUnw14qmR5/Xw9kCttx8Dby
f8E9LcPirLxzwBZDD3MPGHrvYLfsfi27ajOFWPS/HFFcTWklrH9v+rcljDqSey/fkf4l6AgZvxr1
rte899GNk+2BIF9vdBC3p3OasbxsShWp1J/01VDRtKymUe3N8GXCdDicz6DWPUn+bHvLFZhGJRg9
ORHGZxAznGw2VjL7VMgDZbOGQz4M60IRAbrsTqmVBX5lfkFYKPhYFtU+YwrpjhfxlZlfzXRWsRox
rETb4HmtHAFxjL+dkmz6djCIMPmA1CMjd4JMkzPdej7+d+x8/+sX7AQWwgJn+Byro+vkA+dtUChI
d5+BS53Ei9o0gU3hry89nSjbk471JL3rqNnpXtNSCgAgaRAOGARu1meW8p1UFh9IgzpZvrXhSOBf
qTLrIsrLSZwJZdQMZ6rALQHL1ZJ/oFejityhSjNnFfESK7/TkiQpcbfEpthXjTjR1H7aU5mU1nbp
ogPAIzMnFIhIeqvrfwmUAHeOXb45MO7LTzSgmW/hCIySFj+IV6sppH+idOhL01U+UnHdlyon33sf
Gu/2MSgWCjKLce65XMF+st2/Po7i26cIIrdQLvB414sssqLrRLB7A8WdLt8ip7kop0Wo13/p15dv
mIT80z9znUHY+MEFxCFNNQIFw7O9nKRrHcGuKj2jz9YMDqsBMijeLALk0Wis3h0hx8U865pPHIrv
0am5+Zvq58+9ATFYZmY3u/2hWGkhXptjbsORamjGtxVeHUCpCp2xZx2Hpkh5q4kkHKyj9IvUEgn6
ifgNEh6zFK42sJjfPCuM0u7BUPq+mNAr2L95JxdU6Bw4r5UMyqWxKUO6F+enXBwDXHxNzy6FncmG
2sHssyhXaYGPoLmKpc4sSElmkJrTgKeblCLAo/VezScvrtLBq3ZCrSBYQE85Vjk1skMPbAcEIhaQ
Y1Pa3yzZ37ua89LCc8Mi+v17dGe2yv9UVOWGkuFgzKKRPEOwNy2BPkk3AHgQOZrWDLUkDVx8gizn
Vj+srTzPaX3SjbSYkw0TQKxCsol58sQyDNETd4hmcnNXTJZzv4SqQ8Dgv+BQ5KqcWqfkgvK/HEJD
/+inYeX9h44WWhhbnDCDzcCh7vqDNE19b3Axv+E3anx8lyeTuQyGEz34+/NGtohusP9qDXkFIzST
q5C4fPmLt1z3eW2npV0nqf881e51Dw88HQWU5oJSJBXP+sXux0MX3aj/3YUq5Wfmwy6jhIFzOx08
c2th4qilnBsScCXicd0YiaMrcsZlC8Aw7mzfzJ5kXLvf7De4z/KZKXw+SIo0ZyDhQzjjkyOJoSyW
ErMbZJjX8qHnt/shYPnqQJPPnN6cpsZNOKZpVEvRXKM9I5NfuVGJF7zJXKyJ6id0IO9h0ArBZ+bo
cr+V56U+TGRjosFG2z6cAzjSoRVRsE9rHbZtSPQsnVPNDQEBXiuZ9iqfj++ypv6MCGMa5WcUue19
riffY44JO20QMTjWKnVnZcjl7WKSzFbFmoQ/Ech6OAerb/Xo9guiJRpaH6s0125QRA1uejuiPDeD
QImeSXOJNVmJtWNo7pSdbUEPIKLX9gFSaO8b7oOSiSgJxF0Dv+J4q9mvDSBviuXhClmBlVvUKGzy
6bHZULgi6eu4+ssnRV7EmxPtsU6WMd5LptabidQrrbxa6OMAyce4nTojRGRok1TF1q2rkCSAjvt0
5uCUP3t+zlDtRaI1wPjIr2wrtJW5b8jkM+VoAW/BZPWgUx7AJ4wS9zlfJOG37eMgTmZv9D7kYvKL
MlvJn1dbPpRG5bzIs7BpUVmCpLljv/XYFlDD0S1JA62LRS/UuHgneL0dxc8peEHIw2C2llEviw5R
xobUu3y47eY7Wj8ba2/rFu+X2JEcnbH2bxYNB3Ls+K4V6coQNwpbxq/TuSQGxYhUkkS7U69tat6f
a6Q4+hgKACcUjSiZCfplG9Rg4TfE8C1IInHVt0ZJPvA3Wq1vuAa1NoaXNG2/CnCuqxSNMsVoD69X
yHIMCDZhfJGNp6snSfhpkyC0YTO9kLTBCJI/mq212oE3L9ZpzUETtnTM7NOIvOFYOWIv9cpxH/vI
3TZ15NkcwvcsHgFnDYIA/8K0wZKdsb81A0RA5SGY1B5G883182NA8cYyTbT5Hks04U5SgZLPPWil
vkABwbD2Dwn2h6XX0j7UJsEml+k4ay8Ht+DYb9A2m4P1K7qoTAE+1vy86WX/fbA6jP8rl6wuzmNH
nEZoaFaRn39iY4VoGHWCFSZnc+FsSq+GwDmUtcsYFzHRn5OGawOfc9b7DDTfPQp1My2Pku0CuA3r
N+TFu9Mwu1PB1WAkuXe4IlB0GO22jZm8WK4LWQu84DvlWp99YRXKysn04dQi8KrwDw4iChCjHDXZ
W6xJ8VbuBpFnIB/4IrAVCDzuHIahr/rYR/Q+JOm225TrjK3c6eR9Z79Qcd5outSMJhjHWqhHE5P5
56dRAX8qW3E+ErOyF0UuAyVONuZDuPAmzJpdghi7vzivedCSsQxXCFzCHwnPy7Fnm6Sc0XtijBca
+I7u4uZY1c4Tvs9FAFpkkCqVuPZkGFqsX2rk287baa1WZ0eJORa0VTghq8gkKPLs0j4JPWVrfAYL
xmNXqrNhG8dqSicASu3VCqaq90bNkzxdef2RvSm7aV7sRNvobSYtL6bpfxrbES64Bs1Mvz23POSh
+6V1je2FrtTmOGwAyvcLEf+snWmZeI+WoRLIz0yXORokuDD8pIxXWypRPki7nm4x0CJHYv/nD4ON
76vtEq7SkqdKO+sQQNm1yvY2r4AbY7rZQgGsh+Ouz9yK3467YGg6NZolvVFR0jyQb94l2TjUim+S
AtKtZKL+ht4tjKGQS+QQTwKCIAnoZOichRYDQAmvoonS15xrMbB1jT8j6OA0+Lkn9JHTqvP8+HNS
MJx4PRrXHscUrG01PtL4fORZb6+CTIWCsUDxRdJXGEFdWnfEK577jlXukdn2pqu4FA//YYx6zkqN
LNoiWk0J93JETWs6ThvbmXecyQs3xuX3ErcIFDCiC7BsknpuBDUdUqou53alSYI7VxgYq4R/IOkM
6vXPz0JkVfT7EN794EJNO+h6LDw/+jeLVTrcVqyeIoqUiA8uWtCHRxj1BLrOCyPUzaC+cr8yCeFo
/nt1U9GGE0ikJgHJqlQUgaljB8HL2fxHEHMf0gwluXjJlLYXPv36pY2YeIndX2KdgxWCiIDSsCH6
1KwsiW0S9PJgEbn9Ur/mKogJXE060lZUGuINEwqr6FKPKRC+3vG0sUfWgRELdHrFOq1PaizxBgln
rvrthUAKDHhIdOrcfxvokiTIRe5qYM8AmEgMtxoatUOoBDDMZxgPQRkqjjfI9So+VUYtsugCC9Sa
23UtDUF7vCfv9EVv6SK5MjmxFI8NNA8Z5sGn9UN9vXtq2v+8rBERl4afAcnqy/uYJ6DMsCr9pJvm
ymKL3Mqa5Tgjz1ZV+lvmhCpP7te4AIDwy6m+IufuqeyuzsgN5ZKuDFvIWvXMwgcCb3d6sua3NCG3
gwDZvyHduMmpG1hoXuALy8b9vNM7Xqb+qJDpOvAAAeLHHdfW+3ELrVdOy59zQclgFeagCW22XqRi
LwsmcetiEA2ATvubog9hheObIDSfPNFlLkhzeXbZx9cliTlUrMEMXwnfRpflETtEcKnA26bGaibU
CTJspX1hj5CAWKQ8jCz1I48YIaL8oEua+1ntknQ53YhHYiXu0ZhInJLfWrzY8pp2lFYzw5W9HTfS
ycj/Ffg0SXZxXg8ZxbWhfRGzAy6TX1LZDHMpziZ+k20++5wr3YhqH8WvP0979qJcp4kwLLkabG8n
iPGWYxK16ho0nXBMEdZXTDJ7HLdfCNebxhooG7K10QyjTYLHta7EQ2972IQuCZIvES38Xk3LZXTo
2L7HbwDeHhhfNbS9ukWfsXON1J/KNddm/dtS17h4QRAgKAdFzMZXtyyylpXFMU3R/tjyaYhMm+72
OkTpET39w7PnABm2YWtz6yyyaEjFzzvZf1Dnp2vXo7AQEm5XdQFOfA+5jhHZWccll9O53DqC/OTH
+megrfG6nCWMKa29hsavbOfmz3mEOTFaJ1340oJxD8xoA43gixBQrjBok4dDv+j0+vuygwkI4JQn
UTQHf0Ppjfoyotxm3ZFdVdPRzH9oio5BPYwlvJZWvxLsz1nLSQXKBELOYZE8jbfhL1lK0Oi8r91r
HE28r9U20z4RY1b4P5G0i2bbYIQlA/7KUL42Hy5YSG0f0vRoFQKKszXSroNaJ8RP1yROAJwbP1sJ
dGzNVOy1YHBMYpMvqdmQZy1EL9FpdYEe6ycbVormQe/pRYddQeJPNEZZI7UublnWLAQYGVWN3uzo
i9lsRoNo9PqcVCwEtPX32T+PmZ2wQ9J9PJipDPww1Pg7bsx1ClwRJ2xjKijuBeTSSQ8822PP7nNk
1xj44KSThNPUZrg+jza+INzbe1UioFaMrhPh5vchVl7ZWcRS2u4agz1Zio1NLk5xoaaZxVWpIl4p
qQhoB1N5Mpa4e3dqQ4b8LJtZ5pz+2KVd/6JE9FyEAgxgSY28kAoX4g3D/XcLJgzZSQmcWhtHbXVl
aD+uUsPSk0a+Kif2uETZzAqVnbgptMTEfLAfhH1m3oxJ7ASURU24mfnHYEyhf405yNo8n/HTEXmb
YzysuzNS6MK+Tco1sQVoXK0KWcYMxeDk9IksMhLphPc6BvpcQGCe67AYwkOBrtCob8Jg1b25G0HY
m8Q4i7eIKkXR6xaKzaMNPNmaJKHKMllRkgW1XbtKeCFTVeaEfvn8Bl9ngcwAYQgRuxGExZ+NAJEV
i3mGvSmGm9sZfXH+xeF99pxQwYLQ0Ktm7M12BkbLhlstlwPB2F++0dT+PeUsCXZvGMotZQK6CgDt
koE7d5PMVcEdjzrT/qTJDedQlWj9legIfn9pdAEnpOS9F8jn6wi/wOzVhg8SLzMbDHYVIoLQSJeb
5Rk+C2wLhPywDrF0h0SZkp0OZOwBEKYBVeNsigUbP4ug+3U6zmitaq4YkhX3KMY4/om3rVAfEdgc
EMblEDtnRjIidI8BRftfKHjBlewtgjXwqstam4LZtdGiYt8nYNiUOyo6FCiPSj3K0hfmfG0jQxfH
hqE5zLirZe3h5XAAO/9yFV6J61XXWznWoFb9ZNayrGvDr3rwTfAG//3E5r1o5hAe7Gu38iYcw4K5
l6zzSaOZe5p9e55rv+1fUWZuKOMK2Cw8J1B8FFJ1ITltcbeIBNW1P0SqBxfjxag1wZfF2rtNJva5
YbFFBbLvgkqDA/Dl8iuuIy2HvHBySqp2yRtxmNJJjd71SWpTpIKk3FRcOTpkAy+vsIHlmTsn0mUI
I74TRHk/NNJnnueE/33439jBGifRTgA613aSHuGK5L7cPDCsOxyKXAVGor+x4sBtXU9EIhbS0/Q0
WgGGc6qf1U5mfPp04SKWqU0IbZJCpobEHq/fMKvOvQqw2sCWkLspDFTG/t9XhMgZLYFzgiA47LTL
BfkX9M5sTL1VpFX5x4vdK9EgWgPHUA87us36LDPR+XrBRTGlavfVpsky02YmNfojmPKldeE7x3la
vxhnaNr18GqH6fkcKYtQ+tVlNbsAKE+RBu/DEDCfwL2NpOS1RGTmEKGlty6kyOLf+LMYohsNw1c1
vBi1Ya6A6HaAscpx70LLGH2BLRZCZ4hAwnjXOoL3O/O2NvV6jHbXaV9N4h4nSE6p3DPxVV1jC04n
yGZLm2udWIgo43q6s570eIasOe5x3rQnpyc+Z4cuTkbY5Tgt2DqMa+Wvzm6wlIhNwfcY3ysND+fU
5BGAURNcZYn5u3c8n1zvRWJGBeGxhljfA6akSnun8dukfrltAXDpHpQ/71WedlGZoveQGOVTu0Tz
f3/wRu/TOqYxD06Vt4He4gAq7fpNIZWtezgq8mNof1VzM32cC+fKFvJ0O9m2RWf9VwAZaF7WHeOJ
w2I5lKqFkWylB/bdneCjsbVpNaEG5CMZBol9zX40Rku7EoVIM4yZ9cHEksfcHEjigdmKbpAmbIPZ
2r1HG9Ja2ybbrFHCcUNHtxTRQiDa3F5eIj3W7qm0a1Wxm+0hDcCNNrTcDA8k6sziPC4i1HXTUVgA
omAHiY5g6ItOkYQRykWhU1QzOpTrQTk5dg1i+58JnjbtjbGOXR4pszpt+/CNu5LhjrVN+bJriYmu
9eVDMzpRA85baGYhl2W0sGlDacmJVbUfJeMommMLDj96Kv5yD8JDGUPP6Mk7WurN30rH57UGaA8M
LHs65zjVvSdtY95g6Bu+IlJHBKVZ8mA1dI8eJtqLBqF853t8+LbnbnZ0LSR8P3bSjSGprmSu3vkX
4Q1gRbFlQG2105ZZkzjYK/O8p38WhrqkiB2X+L/bV3j0H/futt4ePa/8cPixAAW70VXJao/DVVU2
GBds1wqwlxDD//K/CtYo2ZhNAJMSHxYViSrbrRM+hgOShy7MPp/sAjM2xiwdKFVA+DrGiJyvl2RL
4f8LrMq5+G2Hm0qLL9XImrw9dGTjEARYh9r/qjUtd9p0sK4loLar1velp+FBVmc4vI+AErVEegnc
1JF0Vl93vZQC4sTnSp1ugLt08SdpkwxpLFQvdY+GDMfzuiIlt2IHSZqDr0wIb344jvTgqiy1i0dx
7wLSOZX75UsRGDCAGta65Ccpte70ND2zW3q8UJpLVksPXIRHmnPS+SNZew8Zdjs22B0HYgtYGCQ6
pRiRbD3W0epjahn0sM9bIjTK+fwlSD/scyfFO/d2nvwW7MTggcBCsLWiO39FLsH+b89AdBbJDvEn
U3wPWYfAdSZeHDMmKJyXrEfBlEI/x9skAH8q1/bEcTtEWUkEhleLyIWj554pbNHF8VIwGem44xOK
znmsHK07f8EvJDK1qDAFP4gj2UbJKQGo0sWladBJ1khqleXLGMhDUeXhla7VnTVFNl7O1drq3xlF
G1zd0j8oD5zHMoHSpfSphzfF0luVSJBft7617yRALc7XBaz3UWQVauBo8/V4bXKW4MXUe87J19ei
Jr0QE4kzbXL6KlL9kQUwoJRkjyhErbUi5RBeWcLE0XT0ptoG5qzY8lfd3yBqHJkny0L8vNgEtazd
uj8HpctM6Y2cjIx3+wrjbCSxGaUa3dwqjd5BZPq1BocU6My7eKHUxJudJltjh7vAvldPuftj1w+2
pylwX/qVYiZekxLU1nkS1cY0yCP0wPqTcyf1TNQugjQVtP/yq1FEsHf3M55Y5Ud4jItK5CC99STj
T0zYL42+aOqygh05rTyMgACkTOBMhmPRfl4Cx3MuUEija1z9ys3w7gGVtdyZFJ3RLeHO/jt1V2t6
7ULGE1DsvoDLaS7ZOkZVA0+gkkarAIiKQqdemlMLNmed67B85XAKOCPt8B5CmALpbf+ZfgKaRZYf
yNuDFXStO8VJDkSHbnJ9PcLvsQRdvV5ilj+Y30KAbFW0lnYxtI3jJB1c9gFH8p3QEoD6Xi692pQC
i53lS4D1savSmMrSsU2DNrMnwSyL2GURE2bayfJ/7W9Vivlu8si7oHeRTMvF4QUW+8rAPAZmzHyf
tOnLc0HZBNL+2hftkdXNmjmBG6lmLzJqymTZbNlJ7MXYGCaqfd68R3GFFcTy4Alkdo5oMo6yt7MY
3/d6n781WGH7SfchznJ8eP4aS4I+BJXdTpx6QK7JF5wwkB/jRffZrVNQGXHvIWttsUYSW74xueTG
zRDmXLWPZOSPJgYKcJhECBsEKD+697JznCrNx6wF1MfgpU8EhzwaRVKQH2Ihj9dtJwNfFlqHX8KW
3TFpKgnjXeH92AcgHugihp3he2aJGOYaTwUCoSGCWLtUooXDJhJpmUyijK5hBfGh3ZURFI2lSeoI
gU2CXCV0CFBROaBqALNkG6A2RGITjqCXsn2yuqaKoJhxS4S7SPDTnuFHbhmYgYup2X3Dgg+7bEWD
sH/W4oEg/mxNQSJtBPDq2eTUqcTV5imMhGlKHuE+ETFp0rKsFE4rvoNMfQvxVPdbFLRy/XTonlys
0pGoYR6s0jIcjdFwANb94NRCSOH5GEKesPxv8KeiT9mj7ITaDzurMclm1ADF2TjfAeuYQy4OEjGU
/TglkFMGWMcblG3V5kzzMTrjIf1/HAopi6cItPamH981C2kMVYpoyZNAqgZTcn9WD2VX3Gsutq4U
cn3K+lS9hOFcNaBZXplWaxnNdMvjTWUKnviimQ1D9FbEfX1J+WdQe57HU1Srlo+207lG/RxrCrH+
DC6FnUjJRRFeH/pjRkakZFfiYmEKwurP9+nQtKqwlVxjusZ+kjmUWl6zUgx07lJb1YlNjsBJh7uU
0szE4L6628ugeeMuiL02uh2AbWB+oIg6ZWbHS+dvVBY8CKVoq4hjz89Eii7CVDMZNl/ZfZnEDjqr
052n2eG2G/BSYHG5LNiy/UnU37mDLXZTiDX1CX7BVUfFylKTx3ujAClfEAURf3hHb04Wb9/GU2Ui
7k7iIJNPLQ3on/4OVVqc48xT5mUqInb+40S4Jp1ITc/rj/aezFsgXAseuXbGOy6IVNPlTAFbpzDx
daTjkzSOPovcKRD3SGYNf522sR0C3P9eVd3XfruRBNDC2boaZqTEjvAoFXOrnZFZ4KbYJN9n/Fhx
X/Bf9MzU5C4mIbPLN3nzK0QZs6gHOF4+4ZqESPlLCgM4cKNQF/0hw34K5GuMHQsuz03RuTmCzg5w
+noAUBUNs4iVovVQvkphrDSS/VaFNFFE9np+F4rQPIzE5xDukKqNy0NCswe2psDtuupNIyLJOaMz
Yw/bNgh3b2oA/sxql7iWn6ixOIomQKVPSE4xCxtJ6SUCjI7Xu5yG+O3IwV1lV9OhGKeJXfMG5YuA
hX9c9LXtCKLGwpnBptTpTD4cD2qbBS8HGNTP3opxWFgXi+wspEdNVXkSvIQVIQjYFsf7F+QWSC42
hPIOBTsjSIvBQ1ab6/qXbVFDk0C3t4oF7EJLR9/WUBH90MIWb9VHBA7v+HX+UvH6NJBQ0US1lO7Q
goa3U7qBVlOVLzbr6XV7CXG1KvP1QsNs9Uq5UPcSrod0OIHktXkpY/9sWO3wWE9p+ho2S4MagAZr
f0rj91xmV5aWrYqQUeSEFimWZXFwqcifBRKdsKrBNEEzKLKCBN4qjsfZJW2zaswkrbEDzP9MjIM1
Cy69dgbQYTRL312H1fW+vnqSO0+PY2ViDN+CAzApbj2Mi8bBsZPcZOzjBjd5WgFbsd3oJBTRAH15
QGadHiiUVPgMCSpzn2lH4zCAA35ffiHiNOEEiMyi8WfqHdOUNqzHq1QA719+mAjQ2U7fcqowyIq4
M0VWB/4/oy2zj0R8mp436IuEUIpo541dng/yvAUCShqYbJYojvqA5I4nswMEsru7fJT+UrYZA7WR
+lp8gfx0rI1HV8wRZcaiiNrIWV4weMJRyN8LogGit/1cOy51OP7ymRmZBJy66wC5DAiA5hCHCV9G
nY5+qBCqEfNOKKwzlNa+5r7MoPuB2+RDvUCBFSS/L39pAmZ5yrItAuTNSxbsvC6tshmRYWQmcal6
HaXcb6YA492f7yCn+/f05e5OuQEi9cTlTNzZhz8kwWdPep9uxJkMXF7yidTkZWsN4QxSfXieKkQj
nf99gdo71AcSXwwmQo08CYl5fO28yGRTKqpDstSdUeEZBFYCd4il6nZ8BLmM+bh71JCiv0vfH5FC
MefKZerdWEMDIO6JKY8ynC7E4+Yvwr1eJIw57PkK7aWPmuiyQmlYs1b6aJqQNkOFGp833FwTvTsa
D/7ptUgf4ytSWpqLIFYT9wQiUnuTZ+/URoiCA8K4Psyp+8cvj75N0CRTc14YFOByHPaMhIChjm9v
YZQiMWBE3r/ee4ffvbCvTTdNwxRTMjy6CdAqN+YER2iziujq2P3Kd+Vux02jq4aaXslJARwtdBno
F0d2OFWlc8iqvK6iJ8Y8ZSyYf1BtN6ICxcoGePEKadRJTXntYIk/6ALwO/bU1Bxnt0aNskME296P
WB3+1iKofEGF80TLghtG5kurNmey+2eMIiI5Q1479LBjTwTA9ZRLwL9kyfGG6t58Lu/NljPMatCp
gVC2YsyN/HKHV6elgMMzXgg2nWxQOqHWmwBAVmjkKU02mrpVb9SV0z6OzIe0hdUjmv7F+1HkW7os
a+oWayt5H3MTAfpZLXC1iUCdX9uE0a7OxWqBr4o/fJ5CaG6apb+EFQqDPG3VJyuokMC5S37Ycz8P
cM9amXHQYjipyd6WKT4fiUajZKgDrchKzbqg6gJSDIq+XwscspVTfNtkVIpoOLUIZ6kj+ONWc1zX
TBqc7VrgrOvdiad/4QZUpSo2ghwe7gpYst6TByFKFxNlNqpKlKQjtVN8D2QFfm5DZoraiBsN5MIl
K7fjzmIFPt06QVZyjP68DBoB0fl/pTE/7eKfx2/fQTJp//8hBOtuYUOSepdTHfmFNCoJ3r+cwj9v
DsIDt87jYeCm1qwXdBe9bckVXtUQk642HB4LKUmEAiJ9lMPPFSm9anyquOo/de5YV5+frBMVPe7s
H0t4P7zl4FQslB2uiADunLumN2KoA0A55EYUXJeUcaWKRuxxLNkLuHwzjZOxIZdHVIJRzMhGQow5
JMuc18QLlc8m0Y1BPoqPxWCvU1MHVfwVq364OtKOsXyD/vVC9Z1a/s7PFk2KJ80LOQ1GEpCJcmyA
ExXfRfVK7Xui16uUKGoFUEFseITxFT8nGuHeUbRf7iy+1Qh7W9bpuHARsSMmqFgtXzfvjEqQv3tW
aIKdzqqliPpW8IhMypRZ9Hp/X+0tf0106gbUlLMHhGhesjREpiNuWMZuacB3DxqBwXGGTXe3nnPR
UBQxHNRj9Tai+r4pr44FgnyGp3ma/nfZ6wdzJgqGM9Ng34YnoDkQIzCau8Ht4NDMr0D9E+j0uy1o
c6XfsJ7l0XT+27qIzfVGefr3Vxou2jZ9n8MRWtzFB3zYXorvOeB/GzsVq5Yf/zaghBxn002gdNdK
nOn/CIqqKr4I4i/BSxT0h3t2OIPsb9YR9iseieYlwCc8AwsdmiJRFpbs8226fwexiKVEkTLJ2FNL
Z+SfjO74Qgp7/SarUoqFdvQKhS2/nChjc0GBal78cNbLbuipicLQZsAplvuz79gJB3tzZa7JwB0l
zjKnrMGzWe9pXWzV1RUkVeVqMhdmdeBogVZUUwLFYIgb5rsejsai17PoZgUqACvUe8EaShn1nbGY
wH8jRwGxJL8ViARg2Ua4K1ncKN7ox0hXs9PTMojhVHvs7APQjJDDxq9wjk3la9HzA1NmMx09tOgs
V32DTSe18EUgGLK2GBkZ04WfR/Gj+BpbOOq5EeW4Z2s7cGDwylGYVQ8M88Vvyuk2amxEFjsM72Qp
HgIKuHRUq8IbnO+bScPMRKzABXLUkRRF0RXnBdOdTH6AOqu7jxNefp/eH346qUGaAG02SJaOs0BF
CBGM0bgqdvA4LVb5m8b1G4iYT54Q4QGFUBZ3EHrgw2LOy73I9f2v6Nu/6y8Un7BNRlZ/q0BIsXvG
79FOff1BPtJxRqUIzMI3hGgm+7mBPhF4wjx50cxvXr+Ch+hETh1GzrvPnLcFHm8fQHrVPOUWB9Vb
ArVIgNQjDNSpPzzSAzoOJw688iJ1uXH/UV5BZB0zSzrDVoOugLRLXcFfRRwLWvwowtJFXuogOswf
ZeFnJfnjLBH/7kB4aaonML746SPMXueOXrJ34/WblkF06hgYQ9EJ8pdpsqj0/jgXrru0PfklMa0K
ZkjEKxlC5fY7HCOUF+A4EO46dEtXZpTk4ZkA+j18e7EKqbWQJMT1aV3tmig2JV5Cf4K1gjNVemy2
WTBWjg8LguCd1q6YHJqfuwGzwAYTLyDQa7nUUQ27w8ulaxPwMJonrInp6XjESY9M6EB7/NYC4RiS
tEMgMxVZDc/u+U/4qGCT9Q2Bot0nTcERN76ygtJTdXIKOu1yCCfi5tTeMjgyqkdznQEjO0ADqQxR
oEJO0+W9/M2g1+YjzaEdKxp+ActenbQgQOhEI2B5i58XmLKAtkCyrPSQDeyKku+rzjYLDsyLIDdY
fUpInEDX9kWwQZrCOGda5JxPWMuVjrMupv2yPcAe4h3FyDr5RAqLpkWGmR8K7Kbz2RrLcGvblFk7
m4uIaK/dv9EBo3hyjRdPPXzVtoXoHHGcMNWotUkcrYQu9dnY9Ckl/WS3zIFduA29ollCzX+tUmJo
AeTZuML2IsrWHYDkjI3AqHMkflU7P+i1uIovtVFE02XdHSSqMI2Z7blID+k+Rlt2AC04AlW/7GRK
aRJo26Gxh7ACVo5qC5u9sR2rWWWd1ICTKEz7aa/S/K2oV1C7NB9xPwUEZKHh/mXZzZz4ROJufR4d
XCeeALTnQmXllYSzFdOeziWKcvxY6uOWqq/yjJAujflQN5sk52rqbGaKwB/SuZr4N2PUAKuUHmRS
R8Zu1RK1QHyfvfeSo/+ezut//kEE8Hiop8u/VTuWg6UCCVjqShVmEt2U96fr7jq7i2Iz0+LrXtmk
VCaat5QGy8IIVvDJi7v2unOU9T2HZh7Q/TE8waYAmuCL4/cCEs/LjYZY9Sabm+g/93gC6jdAmMox
znvZOzJM8if/x+cCWI0O3+wRpHQRZUlof1UZbOfdPA71wNvOM6zUeC00hcQPSDjfK5qbbfbQxzbD
wkhhPoLzIiFsQ0seUMG3GKM0Ug9KcLGX7/5w0onROrwXUYXJfosy+RYQIJdbDBmVlmCHKZHLMeTS
A1AGFHJH1MC9BanP0BCjLZKke7kM8Ag/lvThnuJ5m37D+RVU5+wp4bHlI1XAEadSGlfOb6IZswJG
YkyyEjIbhJhbWFS0vgQJ667q9LDd9dGjydd9J+yC9YlOahUmadWiJCYIcNOUcLbyWwsOjIMhJic2
DN+gwekaRK/XT3Qs/D3UO2ifdofTQgEccb58S/EYpJhnc9Ja+se+KiWsmf8AbGEib1ZjsViZS1I0
bXuLBvluW1oXO3vKu6erqwE5DqhhlHBbNiNMIsjsWbNWZc2tdHgreA4MHyL4DUJvl4yF4QW+rlTm
JhRJuvR5I93UwImy94MAZldts9ydcwy1UzKMf8eHPIChFmf1NtGwihBOIxz0QjlN/Z1Rm/z+nvm3
Ub8l6uJQcg75PVz2+e05y/bgbpdYNPQk48f5GNBfD0W8J5b9zURlYOXz+4/GGwY7b44cWun2fq/R
q7mcG9uylGFOlZNBvyJOv1e3iD8MS3MNRgRDQS0j68eIY98DAeElTc8HohmLsz7SuZyOSwO/ierq
ZAjaUq12RPBcic1eLZvpDJujekHJWmYXLpYWbxHiPS+hkOuz5kiySQrZAIJNhQb9payViYJKc2GP
tnToaAo1q003pCW0KTUcICfstDnOKtxVAGBgYXVUj+xvmgA5QeBPVUprWVrajQbXIZU6wHC2IaxB
flNVsLDOlD0EKBZO1ziPK4qIb0RUY5G2dvZk+CSuEGOtEnqisB9qizSSLH++GmQxSsUsMCb7o2bK
ZwSV0KUkb32pHqfWf85ytVmw3JMNWhAk4B5S5UEaAOs7hPMsk4UC1QF4qhQkB3oUU1mcnJHBf8Ar
3A9jQSXfoxaDAHhSTkA30nvAXFh/461X47zFjmeMuPcMMZZ3DcOv8aegNRenbeVUglxYbxCzvPpQ
v5ErMRl9aiusQwj9ezN5MeoLIru5YsZjk5PQLUONf1N7qADro3wNZvVdVhNCiaqT5oZoM3ix3XE/
5Zbs3Ua1XWSCUIbrKolRlUlulNwwk1TMJW4CI4bQNuyB6DWIqrNlT2u6V+Qonyy8qLbMNlbF5Dd5
GaLvYRnLnYsXzhKbqs0sn62s6lNc6KDwxFdyFLJcesFxIU8SylsTPQKeWqjywPv0i5pNfZ23pwaQ
/kX9aYHG/BWmQWYZZYBFPfdq7kyMH3AuZrNqm7WzArP1kgSMErasSkueI3Od9XMZhxUHMOGw3ZZz
Mt3TLkuu5fYDrbC2J/LjTfnqEdNB05RT60du/qpuxkHVyBkqxplHYZLYqN7wQ0CcE30pPcfqcIH1
gQzzuDHmufdSFubKibpQnZpdbLYozidtjq3RiVLKlB9BZoHOtvkYIsv+obAfbIWBE6LgDH9reDRX
X029hdGRM9iIywoL/7oJcqReT6rzMaGUv2SEpGYvAFpa9KUNfYnASrSsG5D9vk3P6IDbCRXa86sy
D1q07uso+0ckv3vSUI/eoOfNgBLzLLhR8ur+/LjDODcL+gFkyMi+JBn+GbNwK7yVxfMDLCSESyVB
uLRPuqwTPH5X586PkrNafArbcx5a8zSJqWLaPTgGaZsB9GsN7dxfTErsgmdBqLs4s0CiHtSFcQMB
8ET+wja/AdD98gd9qFSv8wDjmfDczbRjLu7uQEzX2Jl2RG5154V5dOil96MVNEO2LUjfZrwhAIJL
ky4Tz0dyoo3LHp6oJ+CZSUKbn4alJLMkNuJt5IigcOGPPaFavmC2NTUvfSDSLkxQjdeffBpuzCx1
hhRgIIopeg6G8q07wuY4TxcFt5WNH6RwPYyXuSzJdIxBVt+Nti6q+EJ+8VhBRcGnmuV3JYRygn38
sNs/Y113b7A9GdEuCJ/7EsqpVkTWTzHbpHT1MMqSIRyT1oiTCgX2ik4sywJcmU9fxIHupAFVi+ID
tsCrnGAlumhBQ9SwgUIrowIhuEO4lpsphfEf0bfT8a4qWbQ/dubpmqXU06BAuIIwyR84DMNCm636
eDa2cudFaiQciaRYHwbrLNm1hd9GIkWRr4xv9AYwOtu2GaTwxwKqmOS0KE0oaT/k+kGkuMXX8abZ
EwcAOErMHR316BakK/2BqI/F9lIDOiR7RCvvQo9ay1jYD32VR/QNB+Kw86ngAcTGkvZ31vHAIz58
+TNbi3OhCDIWga2h3SBi/ILmeuwXipA/3/avIBgpJdmZBntAV4j8EKsQVEHFYYk/kvw5A4Lqmw8f
LnNo7pyZE6od7S7dI+6QePGpAiy31q4z42upOynqOaUSKVXgo35zPIpMAcAq1423AqGddIWOR8hD
wKzMr+ELBlgVoYr7+tQPypovmrz32GgUBf046U53FdGUV0tSOGJGVuaHiX1ePEIL6aSUVlvhl0ob
4E7pbdQ6LWnnWWkV9AUuG3MDBOw00aU0oEfsygQ7B5zi41/JpnUxuNXKyDwuiJZ7Ou3J9hx82j6Q
0jSB41/FhouKG2BXLwpsg+dQxrlI/YfFdvZ48hvIkkKt/Q1FZF+tgSqHwZPmZAbP1ewwWGd9g4OU
MnIHAmz8aMw12PRyka/QLdobymVTwvGuUknIp09a7rDBZh1f6UD4Z66ujA0CIaIQiFaluexCXSw+
sCblDAe4ApLU2ZjPqCnyJ5e4Gh5fgy7h0A69aA9C2svnbVdW82k8bBlm+/fR9JcsaCg+GOCQ8cyc
YKxRGofJBaMJsz4EiMxNeLO1onYKc5a/DamJDjYNd24/AVfWSItRi0eBSS1ZZiyHGhcQxTZ5w3MB
vM2lJu9xsUUjANK9Y7wYxPihR3sv/a/w15buxdQHRCoiFaaXpw5R6mmF1lbx+PW6hyJSC2DyUXxC
y4azagRFP5/kj07RlARaZ5c2ueKIPQZRFYVysa0ZRbctSQxA37A/+PZ5wy6Gx1H4pUcprtO27RQZ
9Pt/sRzeyZPZXk9f0HiuQlOHf5cPI//eOUM2b1wk7PA1od+w4rTJqQzosF2FZfm3RRzpe0iSAEiU
CMN2yW+QnqEF2YgQrMw878Byrb6/0ZsoUeqTERdv1YZiSC6Dd2375UqCRkRFyk2x71pTIknsWrTC
K3qLtN3NvoC7SSnVFXwBrhf0kXRd5cywlSDS5qXBICjV3DXknSqfIB+7rtXLFQRKtvwyRMvQBFCW
qsyES8aKC1TkMLsX3VyRqJ6dr/IwxtMzm+dCbujdtqB1AnNJbpGThfC1vdeBYdR6RGDU5qmxQ/+l
QQezQfgBQMrMClSjjTIsAJwkmBBQmJU0QZuyNDEAHGE5KNkHc1GN/fYNs75+mO21fnv939KWbQ79
T1hPOIb1t+bXVitiL7JStpQGd9+umTFS68GIRNR+zf4rzwBd5fkA1qQ248hBa9si3KgjiHnbLFF2
Ur48xq1Bl8Y6sN6WXRdVI1ZlXr5b5gjv63VKGidGJA5siINogKDMQQvtNzchDrKVSqZV2wWw9jZI
Pg9bbDEwHU0PLcUrdg4KQFjTbsFMjR2OKHmLbeK8xrSV+Ip173sHRnadhbNg1Ty5r/X1ZoZ9+Wki
AeBUhymiEDFYvmmNRzse0oG4ts28o4c4aFDiNHHp0N9kIOcmEkDQCTviidWoNosuzI7kPpfi8zTK
nZLdrSsuXzgP5FAHWBUrRJV4HYJOQXgGmyz/K3Dc4jPiWZoTpcgtaYtUvUgGPbwkdIIlX/DVFMEb
4gzA2Ilq02PFxrY3GhixRkkAMglV6zY1/uGKcOBymYgCcpz2WGWCVftt7/a2iAHOJyIJzplD+k/b
xa5s8+nrLIsJoptgLo5PsXFLmyDteQw2iSFZoBr5ine6qgaPD85xrXFpm+7T5yrU+xLMCXPjrYxs
0eqBYnsKBikDFcA8K+Wi5KhfH7Pp/Fu9KIBdnjmbL2PuufjUs6AQvrsPSUfY5/i5E/ScLG30mKbK
UKOtvihbVYKiSajGm1s08OsbHraLEwAviqYlVThYtKT9KHbRLUwYOBC0XbwyHzg5gso6nuyS4X99
oB11ghlhJBFSW6Vejh62vtu3Ccj+Yl43+GzYAn2somgAde+WQTuQKxOh7+nhme4dwrilSnSzWeyB
HztH5C0JjX4tchZ3Z++B7IFV7NsqBV305OGOdBXxg9E5rXmEasi8r6qNQb6I1uKqlV/PiIwMBb4v
cK4KtOJHaW5Xr7Imcj9acUJ+8T2RYp2ii2TML3TfZK5DzLp6LHMefYQ3VdFU5it6mNMeCbxvrIe6
xlDUUEV3dreAD2D8IJPxwOr49Nl1/WF8aF/dkkhHWHTrD2AWsczz+KeUNri41QDdkFtHtbh+sMNC
0Vt/MXvlNEXtWev0EDAa3jM6KhTflclcKU5tVhxTsSKgt2HTMygXRjoXY5Qp1pdhQu1N5CUWFbVt
xcfEkNXdyLMjc+VGO0eVBp0nyer1gyCg5N0YZymBYR00bEhEE6KiwkVexOa/zejK8WKMBIUdY+Py
zJO+5YGWBkirBrwg5slteBJ+u4V577F2EwqGnNwSiPS1dMhYDap12DIK9kkyc7D6fB3QVbpFUw8f
thms44vrIViwfmc1E4U2GNiqI/lu6TTj6vBI/WDccDqljt3zcsSnxKzAyWeCeibfP62dEpYZRNoG
67bzLPu/gJ+uOf85nIqDvs5JXqex1NCdO/3b1IAUHKLHAnTZ/HRsrx7x7T52TyCQd2R5xF70T+85
qZs8fxNwO8uBpJLltwalOssWuDeRycUQbSkkvIhfdnq9fWgofNXKxAh0S4I/QCxeSU0jF9m6wsVa
GDGAhiMs9kQX9pDGAxmwS/bYpbvm6l242uvk3/3niq2o9EzYNR0yn2c9IvzNmdAjsV8ew/JIKNvP
mZS4Wy+9B0bbGY88omLLKtiFpuKlbj8Mo1eFSZlRfvlZ3Dmzlc4kNfZalM3pFSSAdlDqHvUVR6Ls
S2fvpRvyEg2qUBTF1R5YXqrjCfCbaPwP/MUuVPJQexM7wcOl55B5iIUFZBEb/hpnoGj+dHJFwT25
LN0F3rc8p5J0e8gRwdbZD0wy13FU3t/EWmR6lQ9qBE10MmlaAzGhHu1x4XPxJb6J1VeN9a/bVSjz
0knmqs2fkeCU6AuGhJg/OF3BOpq9v1bJ96yMjHaPj74exu/yhSo26xv8mP5zMePsUxfbIbWFDSwX
rfa6mXZbLjuTTWsSvwcDkHHTpk5ItpHyXQFBCskf40SPiW/3aOsy5JNjiqPXoXyymKIKqnwISYo5
YHIOWkKR/MfJxU1+BsxTF8NkbWLdKaWSLsI0oFpopF/sbbTLsKKsiok6T1KGk2ql6YfyWRLnY6fp
B1qWFKS45yJVenuhLyG5JZv5puT82IghviIbLkzkvBzCivPcvGD2T7n5F3v2YxlonCR9wbCxkuQJ
swF3Q5705sw/J0h0iNiJUMWxqMkS+88Zt4R33PuSEdHNh8gNRog0KU2ngnrMtwp3ItQE7Nl/Aurm
4OFpId6GFecTFqP0lZSQ3JIjHr3ai+FcmXJbnAvoDzyW7WbaPlgYPDKsJCkxYdTj45K0HGf6JCMH
IPXCz9ArDGcohunVM9yGQ6p1H0R4AvBdWLWR+d/3PNlNhTxQ/Gzm+JCNp+NqRcgoLH3s72kIjSAN
mHCgdyrGsaWL5fRaj9HFNyBfHib5HDqK6jFue55NgQrOTM6DHoX+weru1Ak0pxXZf80aPhfs1rts
7DBCLMVgFkx6FyPcf0cfLpcsURqO3PkS7fYw/56SJxP+fl9SIZBtpr8pBVaxRezQKSGnmWHke3kP
Dce+/mYZGkiL2jlWuc2Gspi2CCjo0NKi/+aMWOBOlgw0QG5DeSSMlmDgomvuCZR6PIyFZHAXsZ7f
hkkH59GHB9xQvxfqiW89jGw+tqqW5V8mG4WKz0FLCFd3RHgcURfQw9yIUn3ppgmji82lC4G2H3Tb
kSp7kfWFowpXonqZ1h6f3NfkBzF5YK2D9KK442s/eoDA8QdXQyKUkde22GCJyCaGxtZNuMjaVIKb
wTU7SLFrzV5Ei0ka0FrGEraBxcBsWHA9LVG0vMNTGhlvYYNTJMBYIAdgMSTJ0d1MNLLBIQt4MTxa
hkjpGYb1nJJtzcK8leWHqU4mWc3VLH/yzcWjOwsD8RYncR/MbwcpJE75M5yy6N+ezar3O7SqSbY6
ueMotOf7NyYJtfY4Y94O6W5jh1b1vVjNIF7QxF98LswFF1yaH1jKdU5XMPSymccFzDS6aPzict4n
rTb28O+/oidAJv/6ytTdvNEe9QMcwKEv9g9SRiTnDYCY7fV7o2xEEnD580vkb/GkZx29JA5GIyzA
StDTQDYi/u5+Fu6FhBNc4/aG1I4GOsjYSHpUcppk3ZS+YK2nESMoOUiogN4AEfehl6WATn6LSGBc
Fh2Tzv2mu6nX1pg68XlCiLPTgAN4/wXAthgBKQ1+6M4/MUavOsGNpVkmuYps5BLvacaMkzg9KRBH
Xcc8Lo+2yZz6uYwMjOmSF//2oTEjgz0hw6DWsC5+wu0m41cFrvuy3Ye1zM6/wSK45U38jzj0Iomw
IMlF2FPXsnrggNVBZ+WQV3/WwXsvSiXErCWIZBZQsdpuFe4N6+I4g2YpjzIiRqjWhSKSt+NDoNuD
nuSqw/Py1//2WHD/+ZbNVekolx/wlNHHAIkiLP+EOA1cob+Ai7Okb7I8XFE725wUAFzoVuPMeqc1
8iPDpyoV7G1TBE/6DPADO/hPPGTCFn9IVT8vynXljGUXR/aSNThHQs/V5SEANGZ0EtVvPQGjrTLy
hNZRJgWof6MAsJ0QZB/ec69Wr49Y1Ggzr9SmnnIjs8zx4ksE92Y+uTuWkj4ppEXsGpO4BkZeoC3k
VlrRPrW1wLOALVQYokunr/4FGorsh/afSxN9Hy7QShYrj3P3MYY62DdwGFbkPe0esMck+DNx3fOl
DxsGatnAV4/juqrwbdZl0D4stREdXzCzv42lypP2xGisegj0kKJZG4l+qVXhbWEJkQQ/gfE3eqwo
0Iz3CiAOBrEbsCs8NCSZN9U2kg7KOks3x6b0zBXXU0RtjpN09fWOIOzPUG5vz2+1gTgA0n/LtRVP
SvU+401mdS3tOVnsb9tgBg9nGPGy9xDcLlFa/wjtNWtaRQlbuGltWtmsBlr5ng8mszEArqDirueR
x1bLue00g24FTOjtGlBnwCdos4bSyoXJJq4MBWZ+pnoCqpJOPQT2FPkEPVXxUE+xZtbxa1GXf6h4
eSCsDku6qkRPr1aPUHCzQGfM7MxHUoCSNsJvUVaXUq0WOohXnf5Mwuoi1cpVjgpB1uB6fOMQ1MTd
iMNjHpdkvnHjWV5uv/pm7+ZJAVTXrCxFenX1xr+tnNuPMjJiheCyDM/w64FkHaj1cF7654xJgtun
bGu6NO2fY8p/4wWwr/Ok+W+LWygYvKmqafT7f/ILcclcl/YpQv0gVUBOKreS/cuIUphp8aZ0Fyzx
OJKOnEEOFnSRkBXvDR9HtpvOuKo1260RNyeXYAdFZQmTSZXYuSTk55iPTM7Q+fOpTAt2x6lWYt7q
wvAKQ5A2kx6z4k8HZoBGSoEYLYMgG93LLhuK6x7j5Pt2gm+IXhg9FLwhU9/kdTTd+Pa+/j9LrZAX
bbGiBplrYm7Q7wI8CgrX5Hsdc1ek7cwuvFhhigSzLtHUhTFuLaZXA341nPmbZQSK9XwI25cu7oFH
0xq/SLr3hjT6lIMLar87edVM+GLyRjgxiDyqvKsToGoB1XEDtIYL2XnJLG43G9XWhUU02XB1Ds/W
uBv3F3hVpp5fXng6iykcB3PhMV1oPpdkzOW6Ziuw89uR0YgqqUalauUjBog7ijX4Z+WfOcuRT1vv
wN3NWP9kMZPI3NZHkhSbXj+hm++gjLbTz1NNOVGIC+KIEu1Aajqx7fLu50vFqqqJfJ+3p5IvhS3F
fkFo1OLiAKzcVrUv6HB5err3NgiEU9b6IExB/uyYmRRL7GKiUWgXkT/iperqXh1z1prX6MVW8I6q
761S0dOc8pXHxkCkvKbMFq7GP12okPQIR+b2RoM5LO297W2HfwYIHTEPi4qm6l0ve41remeowqpz
wj+RQGgafqrElwbbUqK7r4xUtNx6tE53WA7TGrL98v6wRG6QXVtzYWrEvzDoXukpqpuUAtP50A+J
pGEFB4V10ngaTnvuQGYXgOX+I/JPZJsk7vJK5ukMdYPlgGuSY/ZTz1/FSJ8tcbBLk9jStseLxrUe
6Dtx6DGWm3Y4d8+KzJiw7bBdhCJkMguB5mbnern3EGvDkO2/R0BjlvVSkHQ60HgzH3ZokGDVDVMo
tL7lmZ1hopQ92L3VAKAIF/KsREjCgUez2qp3eITI8tWi0FGHkbP8h/VRql3wFLWZSUVQjolgOy/H
+bBRuTW0uqQHNpW7PaOmqDOEW7rPETY72/7QiwXtkUSRtVNihMj7T14ux8I98+har9IUjWqxfIFI
mMHeE5Ty7Y5u1U5Qc3LNqtKT3N0cspgUI154Or8uRycpCn0PTFzHgV5Qy+QAKVSc7lSV9z2X/9im
Av1lquLSoXzGsDLD5ZdJMuAP+n7JkKxhuxR/QcLAHloic6XJpo7kwuZwM3TYJhZrZkF2KAO4croP
FQji6If3V0h7WCvT6HBz6jzj6ehDMDtd6KbA4d7S9LVpzOJmyQ29XFhd/5dCO/aPyX3WUoXYZokv
/g1pSvh9d6y2b/pMnfZuVhIN0xZmTw/jGK3hVQQyx+DgJP0/QrqA2RxIHSvPu8JIJu9PocFjmfeC
uQGslFDiHK0J9aEWFw/V6f7aVJAjzOYlSGJ0s1Qoz256VVH5J+f7Ucu8JIDCAPrH8EtMEq/WRCZU
BlB5FetXhBV7B4wL7ZKd675yDe7KESnRHSNnV0so4T9rh9wHKbPH2XPb+tuFekGaEnkhJF8MbSXf
5JnLHD9ZgAcpM2WgU0ZWwcQE5EZFk+TpahAF5yxUc0wWehzssa1O/pFdyX807qWSHKmLnOiPZQqb
8iD/UBbNWnwLE7q4f4zYeJnJIt+WG78672lYp5T2UCFa626uiFmHBUwu4LiipLvY37SoDVW2BcjA
As6a+qVERRbtRcQBT7yxFUlBNjb57uMpFDWLkEqnQLowdjRpEvUhze5/B7vc8ExAeWYW0+oDEpMs
U7sAw8wc10f+J/4TORLkCxMbLkViBaTYhCS2YxTE5AcB+Lg+D8o1LBkJHpEuY+fpb3FNGnLs7NeI
hTen2WiG6Kz0AnhMu1gZJTxVdXe4d11U1WZQ/IFZmo65so+WQNA9DAA6FNN91SYTwM0g8+NqCobA
coSAghHzxutGsPDP0x4Tpx09d4fsDjRILUmpcvYFvpsVicrLVQvQftfKDka0rPYz8zSgjcQnQOxt
nnSTh9dNrqMGVwrGfhY8o59EoeFHN2V4oRoh4g/WfDvCtUOSEz9LH5wOgcJkOlqiLwnZTS3U4630
lDoY4aKoODgdTjbEQZaWJmHLtFalJ2zry+idhZLIzb6tZCJF2hWJ81YbgnXDlnHYXtAbom6ikuQj
iSGFCXRU6lLTsarh70Rs7n2hJR7+Oin12py0MmhCce1e9epcHQhwP9QcEQrdxq+n6NcVQfAXZvNA
Ls7C4cZhKqdHA/3btiihdP7+Nge/sJLsuEzOAJ1TjuTZukpB+bFtkyhIrGzJlYHmq/yniB0lkTMA
y5FTRSOgtAIJsrVxVuOG7doDO1ARsjBlmcrMbvWB0DSAjgJG2Bxfg1bKl5FJ583YcG1hSwjN64g1
O+T+jDDo53jLRdsyYW4xidAL4Bg6vsWed2H+wOrIj9QVA48pwUEoxY4ILf9OIZaxq8QhT+Fw0kAV
dXClmP7QsFseqEL6sp6ACiFpPPqMYts8RmrOin8+5na08PFTf+F/Ql0130DJJp69npvk+VwvZ5mb
3RlajhCsfzwIaxpDAWWRyxH9YhTJjtJqtjdaFMzRTgfgGmGGegKw0Om7BKVRuHaEL777djywkvZ6
qfnloAnnT5eFuLoUY4HopCQ2Xl25EMe9fVntNfX1f9VdkoWhRaaqo8SfuvZaKFKqWczZRgsK6oKC
m0siQSoDb1d3O/0c2VRaXce30TepYRwC7J4VXAlX+vmN8pIxzNjpwuC+x/Rzdd+G5QtXZS1CWh7g
cpehZXhbFxXcDHzfusq3kcO8IGWpWOQUOWJ817gWfXJXUHCojE/mB6wAM6DjwH5JZMSh1O5ODTRQ
n5aChBRO8oo43DYdVM4xunDpeg7rlkTb2Qn4ZjpPmZP3TyLSNy37aStvGg+AyAdn4fPMPr7PW7dq
2wgKMdQQJA7f9jZIQZgkqHzvTMH9TnpOqf06OUiDJ/lrdfIH3sVYEhmFRD97mbf9VhLVSETqMBne
bWvMV3wbxUq8XkSnZMlghyR9gEPv23Px0G/jMc55uHZknCWmq6C8IbZKgz7/al+dAiVsrxM2KqqM
k1IQpe182qGQLB+8Yn2B5t6EtD3O4TmNnFGIgtGOPN2bs2oyutHGu3bDzc0LR/PiNVS6di7U5JLs
TZlfAaS8DwvsdQ1iWMCEqZjOPphUXEZZDHcdlDVJsarf4iVoBAQmyFxpm/txzdMGouQIFaqeV4Fq
z5ctlHrD7irZlzWHJXLrFUJpr3LLIQ01OeAPL6Rp8tdF8PMvwYU79KsmBp66GHMNu1ZxeSJWHbz2
SEAmiAziOknLpwkEIDDzbeWW+Ix+AY6DwqqZ5TQoR+pDUoyN23DfLGEUgbjEsF1DV+OaqgRHZcOf
qiLYELFw43YMscla+hvNbHKWnys2+3FGk8xaZn0MIVIwicvikkEjyCoKtwZkeiVnVMbNw5Wfkj2W
Vlxkp+Q+XbvY32OTYrCddsf0Q3Izooz3Rj/ACVX6n79d89bL2kw4mcN+BGeHDloPHU1IF2Wny8Xq
KPj26v7eXJKrSlhtk8QeD2SOv3RYEHvkRQQHkhE69v8WS6e4oOnzoMy/xlWV134hWTWCgDa1Nqzv
TazbUeO68AvjdtDLrYoOgPES7O0nHhxB86odcV5plncmNHd2l6uhfzwX5bO/Pkmr7erbWptI3w1e
3LriXQ8mIjwUd7T5r5TmBaQEazT7mPzoAIXinRfwFECdNbUVoMZ9I15Jj55hA4EVYXhzfKTPK5uc
ecA+zpe3sWqCik7sKGGZOyXQ8Mo/KncxugQOElNfYSWTTC9cJFu34qMfoGeCCMhlbTgYQUMDrq7I
3EYKjvhcZFHOWlsdix06GVlkPFaOC+j1qkKDUGk6f7A4Mvfe5Gnz6VXBCouWVnoo5/jPS/9zHpG0
Ynow/kd4r3lEk9Q0h64gUPOUwMJd9nOvu9aVbciOeZwmEKVsdB+rY9r8De1WiXa4kpAR6APNWVjD
hxUwVD7ZU6jwMmOQNbtbaUv7L4SitYXViycue/SlKT5dSUR4XbliVHJVhbfj7A7V+P/7UlpoStqL
TXFqj9NjH+ZndPHS2AOfeRQ3uJa4Tj5E40fCAgt16H24J41Az2keiXRbO0oW49G6LJ7P3/PbpMAz
+IktgKrygAqyH+LSLj/GT3IqkZufJuduzYURQWB4YL1xB6nHwA3CI9bX/qhvx7UwHAXgkuWI6BJd
zDRb95KmPVqLZJbXm09Z30gKytNmYy4aZ3SdnEalUCb2denVsaIz4GesDFM94ad6FPuBcRpC5kVM
rZBF7FkuMBMAxbBQv1uKCcrQBK93CGJKQZCaNzyDTlNQ13NHqqoQjrTIZeS+Qm+41u9HSTW1Z+iQ
vTCy280/TyOC+mTf2vQXhEVv3vsr8kP3xpx4Vg3yJnSvbejBJKJluyTaY4avsBS7lsJD2BZfRTjE
pLy82g8SzLdnehdxQtQIApNz2YlMPbNm+buQpTFfhQhRxk4fpDymtN/xdwwPXVl+MONECkbHjyOS
BNpCH/YFRVlBeLnN8oO7oYBnBg44qooEqjH0hExo/0Yppe7hQzFr7zX/qCi95R/2db9RrZjBNHyb
s6araUpKDuTN3hXe4CEq6x9pHj2a/SnbhNzge7hz4aQTOnw8BLWOzxWPDIfhxlJwgLke0Sp2mYsy
2wIfdX517DnQOaC8Pi+yH27kiGG4DGVToBf87tyAw5RXswHqQBhDmyuZP4twMGOmPfd19tvb5KbF
/NZu/s6at7Ah38tuQ3OVRy+nrimUw/AbnlRCrYk9E761vTkY72XoMUy1JITRPaVRio5F8Ko+6u+s
Uw3u25ydiIpBcimVdoHywt342zRCvacvCbCg3GU5vB/mcO/c3u2Gws4jxS6SZB3xWm6WKzf6A+9S
dX5Ur8qHllzY/laO9gX4zNv3dziw2+s7CyaqN7WCPVuZiX+JhoXZpkWNtU/7akcywpdC9a7YkImX
Nj0+opabso0XhZ3VNYIbSYcxtAjX4H66tmXdFQ/9TnkVej6VPIjaMJDPVMVFTU76SIjaf1e4wVDF
JOz+SaRyF+Ztf43aeke0mN/LO2o1+o7Vp4ElrN/bMI/QKfyWTFhHCHY/h52e7UFUqrAyZ+NQ9gia
VO3GzrX5SKbTXkKUnfqID5DHOFJcACBQbGVilEmKAORAFRTEM7DoTiQfRQ02f890p8COkt34qPVl
Pb3Drsla0tTb7IuEqMinCSYsfUxDwxB55FGvXYyzGcFZujNo8LAJyGDot3ocIN4Li3NQFuk8ZP4K
xopR8t7d0jJ4w2erJ0Stj4FvwwmVelIuz2WeUKZ7XP2ZIa7M1RIMOegjhYm1nfF08hcmndT6lZWO
utI1JmiNXjfqrqs/KHUN9eyRk/Mt466ruhyBI1v/BQ8HT1MTcHR4WfxsCQ09STkKEoj5j0NoP/6F
PmGXwFRObauTt3jcERfAwBIhw0Qy65yl47KQ/4F7DEJ94o1XEqsykXeQ55FfejY6LvJMFifb+HIL
C/D34uD0/Az5xcirWZdb/Rm8Eg9TLisZ/33LN6726w89j0JeqZ07t3GDzSbHulhOes+4RPb1zmAi
0YxMw9Hb+CvujkF2y/Rwg/JcX5bwCUFWTozL2GGtak/i8S8IuwJYWOnJYbGhVYUULTmLCjxJSOqu
f6ZDoHanWJi2DUONmJ/NryQTYsrlyJZhpMCoPp3h6Ba1VrbifSAjgpD5YA68KtJf/wnQE0XblxjH
Icu+99FLpkyy9D+kK6gSHg843t9aqAf2f6bJWZDbtXnBfQkNWx1b40dALQmbDw1muLNK4dotIvp8
XAE++afLATE7b35IA4UeWowHFX+e9Niv7kp11cEB1bGVFsxPi+OzohsDtpaZQoEH9ijm/DYqqDpu
gU9hReoN5mEsfZNGupmJQj6pdrIlxmN0KtXVdxopvCB4toIf2Hbdg9tfLgr+X81s1Gv7fLLu+EBi
PPIw6tT2UbylFPhNSpGq8CMzUThhFxIPCzIHLRssmdV7RiAN4h9nkcLLCs/HIFTDpQGlNF6IId9g
rWZCdUzOZphpfNzvmw/+tYYKarvsynACnPzo6oMS7dRexa4SINd8YG2ajriY/BiHtFmvYrqDzMfV
cfCOtR9v9TpBbyqPoUb0O1c3toahsiJUosmmEUOXCkIxoFfxRpe9ZJeVe+uIWRLktM3pGyDupUq9
1TZ9YuA6iuUNsUkqXSd61EWqgj4BYMuMh+i22fRHjgmSOFbeUIA5BEnRHykaEGkqVortvfw1MVY8
iBQOUyW2CV7jjZXByUi+ugeuQneD+s2fKeqX5xlJ3Opnuwq+FUpITh+66Ivs5rKvuhf2S6a+bTEi
Vi4kwCf4nt7ctxRjBk7+diJxxwx3rTyunj8+IGwN3ikWJAOaEp9kFt+DuAVqmZ3SsYZPtKLIvpqX
eY6Rs3+NPC/N/TLg5VwdUj8g61QiYHCtRz2HSUB/sw6pNRs7KW91Mk6qNerdN6JjXB+43k+0QetR
Vb/hbzAq1L0eCbEebr/l4Wb5cMmBXHS8kWcWfilYkn/aFqKRo3OxAhPk4/d6Hh5w6Dwkk3pHwRba
c3p4kxv7hUj8rYyQmtT94Ud1uBQmDxgpN5w7u+idt0RMrLd0ppB26qNFWmmUYA4ckvTeugIIbhK4
1Leqh6QDMZa/k6DI+/PapsPxgB14hDMoiX8CarMRdcywQQ5H0Jvab4Wwyc84wYj5n9mSr6tpKG4x
cL4ocyQtd4IHsX/Y87U9ar9xiK9b4mAPJ5E/8EfYm6pWGpfI7U68nqjSkFFqRiNGyb2S9DD6CwbY
o4LxUnWZW6t56AfO6UuYWqgpqldOAovv9NnRao4j/FvqMTBFJ+u71oiDOPbTjXjH2fcRHAdVjdz3
oNj3zCABJZrAAXF0auFh7VOnm9c+wspfamvrs1F5Mt5wY2Dw6SOKJDDVlqWru5eleh6kLD2/zoGy
NbcfFpjyXvDYuy/5tpb6aolJTOxCi77UJiV9a9oa3kaK4VD/3R8Cwe4tSpqbRxrxGd5fjFhQuu12
XE4kA9UlVr/rfg0soM/y3oVu4dOQyZ/cKnebMBa/5kdtTIHwxF88t6DB2S99z0tPQ1xn9/AEH0Yp
CIZJeoB1MhT1II3hDYtNmz0CSaGJ3dA+9NSiOxk6GzFUjYyJD/INU6fePoPdtnSrJASfa6Zlxex4
Pnle4fTBy/m1sR+0HgB/Ik/5agQfxHl+344MzWi2EhLq9uuOULziN2wnH7ao0ADaFmI5VGu+BGIt
6HdeXleMRtaiVmV4aqTc6TX9rE5NyVEjhyng03EJGNdp5B+oZ/jiy+Z27GYOglqraFpSHQbcgeWJ
vJ+5G3Rp68eXEc6eunJ4JYgoFraXmtGQGihkJfxvQBly46UZN3y+RqrM+TeVJkZR/nrZX6ap8jiu
qwXB8iE2YIYYqAxJqm3WqYQMSr+QvXTnKup7CZFwHVhj1cP/FqvtA6sePb0obrU+f8y8GCG8vz+X
YAUSF+ZqTAm+gVjzFyyPvj522En7P8IiEvErxdzZ8tGgGI55fm8FbTwoJ/d0Mj5YfIUSDk7kN0u+
YRpfb4rB0HzDN5Vg0gA7SbGJGfde9W6Y3BDfAodCh5PIeflJ3AE/McGOd24bIhYZ8uRxFhoWe5co
Eahgp6Eli3hnujM4tPgCF4WwNonCg1Ubfk5bV2DYRfLXPOdyE+/TUCsTKYTzW1B/JBTAVZ2Bs3KV
+Rl7CoabkUzTHoNyQiDeKXAJ+obEGILr7wYj7xZoDBnk9VH+pT2o2+CBBEdMxYT0xl7gSzPgLxNA
gymvywNIPQnqX6eOPS/sUmrrt8ETgZ8ideleb875ZgfImLP5ra82ieKkjog/kIIXLB7JHwrUjZce
dFtfIQfRqNLC8e/k6UDFQr+CvTC6VzG5ViJg0Z5LybkZqAkOEzSbmMDNiTp+1VLmjMb7C5cTDzqN
SHz2ACiqqccERDjgYFpp/oYNcDj/8E9SN+hT1hr0mPOBX+F9sPm3K1HAkfXa3EGaiGaizIv5HaF4
W/xMYi9nSb3FRN8AaByja+S8lWzQoFERYEZ0UeYiv4Vnu+/KFwgIP0DraD34+MSi8oVwsm8a1VTf
75z0yPkY4kB2OS6et6f9K2xfkLHUe8+nY0oFoJ4A2S2XeTmzufWqgWiivACw1mouqLctBWH1GxDm
Zc3DVv3LouQ+ObLExJAmYArW86gtE23nvDmJ+fHMiEHfLC6OeaKGQnIB1WIPsTrUen3kGVqSD5fY
CQ4+QugvN2iwCdnlEUltv9QSGxKzRwj+wW0k6GTPFNnp8OtAAUA4kdnhhFf+x6C4A0qd8l8Mli8L
q38mYHw3wxCIPoa8Y8we8l/VesH8gQ50TWChF4ZBTY1CkVO7tS1LPUEvU09en8MS8xS4FLskn3zJ
SXPiFZnHdoWmmy6+zADVHgEVbW+XxM9CsXMxGXOAJ+oM3USgZ96usbM9t/eu4zgDxxlHDCYg4wEQ
oKYuHZn8Q5EWg8oQaXe9161x1hwE83xOfgbLEDMOhb2xTIti2wvl0+1rqiaiWbNKBiQNFxFxDE6v
GmaZVWwHMvUpJs0f5qO2zuAY8nhRaru3lCf2NhRlRN1EMLGunD5tMe8JEG+YeZLRfKNcwT2ChZn8
dRTSIj8aJWA1qNdQI8hZimUUwL3iOpN2kZiDvv0+GBmKDkC4v+RQS2SW17em5j0d99W8sDsjU6uu
QWyy+jpjM3qKP/Ia4xkuAacCRLFBmElGri/TYkeID81d7vcLFSvzxJ6zg8RpryzeMR89aC5Pd7V1
H07COrtbNNjeTrDAximXaL2I3IhRnPH1CuNuEnT8HUvQ1uhs4QXA0jgWusfkVP4Wl2SF0VjLmkVN
si8oy672kYaR5VkKUiNoIiG1c7LCsCMDZfVes1TXjDlspScQfGNK9eqxNNYlIwa6njGCdue5D9Pv
zM0jpHYEnV7FDgVF9+CvmQ2KAj+C4UI+HUA9j4fEw++tr4YvOM1V1WN40LsMy+bYNLLDul4oNvXh
hhMKC+4fXC5lKr+0WRJrexOFyA1zjJSV/g/q1XSlo/KmMr4I3IIjunZYC2xX7F2jWFC+uYSTgfMr
y3lV4EHD1BaNNHFWUDjk8wOLqm/9cjZ4KziGBj62bpv6DZ09DiorGfR11vmFJaJ6sD0zURf+M0t8
tiCHDfEFUfj9LliI1MJp2VgsWJGKSt5WXfsyh/wu9Dc2YPHZO4qHSkgEdGJd1Z4wBEdqfGnP/mnD
vsU1l94RCyqDZXIQhe3hquUdw0b+Ii2DmUP3XgJCeXztRMTfU6I27p8DaDHu5fPtK5+7X8GQkKiE
k0S/WwFMRk+vDkOkd/PprL1kvqLPq+Eiz6S6tXVaPD2PMKnu16i7gNJW1YNbNY9fkm+EPaa9Ho9r
XZnJbmT4kSHMR+zbE5mILfLhczINWJPdIcuA+3m4Mlc+uXoxZQSUThT8KhDqgUkySEmstB9WokMs
6w6visB+LSI3TfSB7+CmcZsWnxiLst+wh1hXwYKw9EmHek58jXO45KTGqPcuX+4sD3seN3P96Fof
FBM/dwr/Ge652qG/js/d0F0Yt4fsqhT80enF4bF8E3vaCEkzo6Cj3wOGF9pXqVvVWShbw4bgmWm2
sFCokPv7cyT0ucKZ0rqGaH7/56sBgQ3sT8CjP9tWYX5xlzz2qwbLj+ivyuAo/HXtdw+Zbd6ZKXyK
nEgfylk8tLqQymmY2sTBnRdTt2tP8McBlPrBBjScw01E3+dKIuEnGFrB4+dy67T3NFRG1V83Z5dA
wVwmzRiqWuXHDfedOQoStB7cEQ6VqerasgDVjNH1aDHQeJeUzyIpbj5CSQuzeRRZDgk7vXr2X1bJ
PywZMAtRrgFm0r2JUFyFqNgGKbzAsgLTnA7odl+ql2cP9i5wRd24Rz5KlhrJj/rgBHq1ME6TCbEE
ONQX+vdYsRVRMzMMFaKi8uELIUUEGpvR4Oly4NviyD/tjOMh2Bg9AJWV+2l1JrsllbxUPC4qOV8z
xoj9nYFyyzxbN4QMP9sF1FgcCvDgYPfCmdxatriLM2uWkodc5IVEYtgEPUrTPv4v0vDJJATz/UJZ
PmzvVttNsGXXwJhxS8A5Mzz5QSr3oA2FYFtIOnxIKExUFdDvtdyYU+Bkr3Ws2ZlIFE4RsMpnigkB
x8lHmBHa/pSOCJVltx10K9wnFvPwTVpyz9SjcAoCHBRzRFMicEPyZqtCgweEtQgR81Q9B3m+1Dgo
qQaztjUaLZ+fymNQv5Lr4hA1Kxwvu7RbzDh2G04eAv3QPADGAtLCWfT/K/iQPeP91ipbTE4Z+CkT
NeGH/S+mNW7fyf1Rf63bol/Dy4dCBfXYzYQlFUgsrtq/qXnEGXnQXqMg77hfKVL2dPR7qi+g9zrY
Cg5V3dV+DTDvruOXX0BQ3BNZSmry2UEGzGQuu6co+mQ+Ly3LY6bWE+pj3IlijdOwzu3urgKmn9bU
cZXU84a/NkgROmJ2PJOG2KpvySY82TwSD/zuIOcSYFv6u4XnkMpxUDV8Y8HJqDMdNbN+BRWC2N2t
V334K+F9PW2/gB/VGm7n+pWx6TZu6ymUZD5S7xBDrcM/h+n4e+96o+dZX2iom7i70o14vY+TxjSQ
u8Ri6nau+KeLRVh722o7aYkehdhohaxwKUolgGQ9UX/vniOB2Fd/eXeOvAjn8xehn93qJlJvtN+6
SUVzblGk68lQspaupgFEzSgzwHoveCfQFRqYtk6KsRgd3Ce6q9mvf1Va2NEKLE4rjvJ3fYoR0tIs
1P/uimTeqnXotsWzxfjrHBZCwPnSEDuowKNQQIcLIJnOQj7bJX6bx67AwEKmVXIy3Bx4qYuNoOq0
2sh/6AE+tXEkGPaDIBFE6mpmkgS43icSqPXmLqiwX3FYZ4Y7yGS7NVwedfPcFZXzyFhSeldMOTOH
Wgqu6QFU8PiuoUYUlebrfyr+OatI1Haqd3qGVJGTIo+4KNnG8WWste6Xj+17QlZN2C1U4JYV1myy
Wva9/U/QprvVQ8rAUzUJ8zFjHv7HVmbS/AnGCDnVvLJ1MkFrxqZi0p54GS2jWUXRU3gUkwrfH7K4
wXogagDfTNJj97Kck0QZSDL5wXq17VyzSJQQ1Sm8CyFBJ1jqcwZ5ODeZC3tGE92DbSWxtGYk9SGL
dfoZTfCKKSxc7E0hhGTI7o0mAlm1ukJWO1LnSt2yypWqjHEqODUoUyo20WViIWGHHz47tBYADQiI
0CqeLjlMT4b4+/l9hWtxFma5xeYwtumh/wwwu3ooY2p/UpqCSUzcv4l372hLgR5136HmGkhQXsHf
iAGvEDt51lfc1eEeFjdfjY4zgSgtCOHZ18jjY/jzcG2Ef9pwXFVSPaXy+KcVgN2hgp5GTEMuxO2e
kzBZFJ0ubx8J+f2P3EbuUuBV45NHmvzrO0ziqe3mUWonUnxK1qDKTpLBAGNNoD/yOtunKvxRlm0l
uWdmvEjqb+1RVQlhyIUgtf7up+7z1EV2At+Rk5XgKA+DgjevQx6iXGTgP9aDzwAE3+4gdNSJp8h1
FIjNTP5HDNWtIPdUsSEvxDqWMuGTzBe+2JS/VmMpfaDmHnQjmYfCZBo2+juYQV9MJa9G/rpXGJA4
7aazOloI3HQaJAdtaIP+0OCHSU4PghT1302ESbUoA3PycxF6qgHYXdWDsp9COa6WhkZ8raKh5esy
Eu6y1Ah/gem4q2FnqxRRbraRT9UFdA0FVzCbxV+dT+Cd8/sWkrytpDWk22PmC9OInPu4oeMtJ4KL
yR4B/F+gi1swrQACjEuTZG87IiPw1sZfQkTuqzjV+VBltL/R12/XFv2+Mf9qZYZQP7Yo44q2FQ3c
w3Pupap1Jdv4pHwaqq7drCOPYHWstxhHrvhbLbBhytO1sAVJiFnJho0d+QSEDq/v7OUmc/EOuJYS
BdRbwjivCEjLf36tYKvD4Dorby/AgHEjTVhlcRmY7FUo6NHebuPyDj3oVjAb6ya6podUJl8DomD5
SS2Pb7FGjInPaiC0/oylDd/eGlCaQ5jEEJ4mqGU/FXCfdDSDoJ9V13UZGVGvEUtO8tBifnfeHT2P
JTAH9XPu62by9aJvutBJ9VU+ropKtoLweMtTzv0tu6diOjZUXryXO3zqJ0SUgnI6uwKk6xjVB8HS
CYP/GcTIQPw13MAcwLgcZkZeyqdUptPGWwmTyjUGmTOYj36l0y3J/eUihbZFZqsipOT/Ml9lie3U
TDypp8fEXPrMrZHiM4cjyUBVddKh3p/GNfAuMlae2scMtzdDK6obVfarjdH2uU1Z6axs1mG4xpBL
e/jk3XAYrV5Wgqf8rgQIQmuYgbcYTWlWqMrOPUh2NHsMf8FFYMVlsUkvHm2QE+aD4OAJPF41bBQc
a5omOm+osFwId4KsA+qj0ddkFKs8n9rfi5NuUGggVqyR2n8/Ezc7OBrJycA7F0oDKVCizl9ToZOW
AWGe0PBCvgxL/lGp99ZI2815GgcspJg/lua6K31RfGljc+VhmvQAyrXacwiTW9FW2HVtbj1/vOO3
THnYryUbkj1KcLjitIqFQ+/Es47fR0/mqHKmxV7Vzd4uNTBWHbsOBCjp4DrQ6dIL74BhwcyGbPjM
KikDLKJe6XN3rWYgYeZBiRR+YwyebmyCRKtdHVJu56UIPyzGvwNep0p1ayEvkq7FkXgasziWLUaY
IUQjB7UOvss/2HRsuBAa/PKyPfQXcDO+XNATR8enqQqI6ra4OS33okYoPp0KcK6/5X5JsABNZk7r
d9PPhyjW3xu3wdbOd5P7/aU9ARBehm+QjtTMl4dK62/kpU+PO0a0TVEt6TmMBXi9ULx477a4zt36
ejeBR6gltU1fh7A4ZX5A8jNZNppMgMgzn+Owbkp4PaFiK/iPfUXAl+PsmDLeJbpREBkigTQ9u+6n
fo4LvqRfMGioyDVs7Lk1yyJXCm7w/PQ7mCLolndMAyRMxbNXNzo4PXX6u9Unhszh9Ta+W4/H1hdO
mNXaCqrCcd3ghMy+/RmbKn/OTAXTn8Zjkx9mbF7l6LRqnA112eCHq3eznDTtdOUmLjSZvncG8s9P
f+ylvI3IKGXNRAgIiaJxcbwjiqw8etO+rPija7bAfOgh6hS07RyhKolb/ree5G0P3WKaxT69q4sG
xGizb24zlpucmSkd11i6bZbACgoxvQm62OjcNthjxe6YLoJuaaimY8mHNlb7qFZtp5H9ylXHJEfl
FnoP2G0spzGHk8mIVZeynlIz9B7IQE/aLnTkw4jfy670tEyoksxztmfELvJLZF1v5GU/aEDP5WkP
DpBVVaQQpChPtfCNBrhg9WjTnzNZYq7NEF1huXmr/kbiBI9aUu/s7YAN3jAYwx9DrQUbXIkwV8wK
ipDZ2KXIeNK1/QMlMtlDz/0qZNMgjiG+XnoYhkgM+/8dfwkOwHgdSuyGkwYDI2mj7vNyBoXVZxys
/pLYhE8IRLUrLPPTdky04zLyYva0DK8HV3iaBCpiKC73qIoWDYcUtSL3bbylSLxcM9oEZCDeyZBB
DUw6TpCS3bjiInK76tIskQpF2bzjyxomSGbZ5J9xyFrkB9MokpIsaH2k+CZqMyzWy88HfeLSlTv0
x6KbK8J7uKagqVMwURYhGwMCaYzorOcG7SsE2r30gksonHmpB0Q3DB76tUFiL4rvWIQgb9jogRlo
WqIBhd8kIgy24GfmQG9LKD+1cE0kfrptUDHu0hqJPinTcKBTH18ykoRpKFai2WTrbcPgUV+98aFI
CLB39yQgHSIQuL6l1HqZPe4sxBtx06FeIxWifrvrO2m14HUQ5hzpYnmRLHJt2JvMJiXGBbJ9XcAk
oNlv1+RVf1/Q52E/FbpgXCK/HTzVbIqC3/WEW8kXKhibN4ckgpm00lxTtVHEPjI+JBVkFaBZOu+y
kR3f28lpaRwIHrhxdpfy3BW6CxpK97p3Pz9TZPIRkZlc+HIjGpjorz4ySbD8lJUbKAi+xN+nHsUn
RTS40BtfGqRw2263rRdgvCsbiJWyfb5SB62DQR6FXs4iWhEZHH/xS7XRl/gYUf4K6qt0Ii11nhdD
YYJ/JwkvJU1v8vkv5G8IvhTznnBy1iboUVrMiUH/3TRVGTpKUQnoQy7Lgxwvr2swCc98XwPTTURI
kVMTEx3BmZAbc0IT+jfV2wPtMPc1TwuM7mgEDJpy7EikQ6Kv94e0xXQcokYEYVzwbfyzfuGLCELr
AyJWVIaAjSSUhPJNpe4tip4I0KkWisLqPR5texA7tFyq2LHk6wiyymxCAz0ClKK2wK9Y81ZQUg0n
R0JR2EGlvTxWPmzepx+9wldaxI0M95/90ME0A1wAGHfdhxQcCUIj6F1Flsk15UP9BauK47+hQnZ5
EdSPCtq06NRn4adQ6Uqzog8DhyX1UmQaQ8+bAHKnsm9EyyEFBYvp8K0buRkh0gh/3OjiHidVIOvY
MKK88MdIEQy25MF6GweHZMm1P2RVgTXI7iosQpzQ3bXE1TcAqArojEgMzNdWooimHWj0emhpkzCP
rs7jicmJO9piDsMCmr9uxoDYiJexnFdcG+7TSer3EUqAvKCiblc6EWBXijcMTtGa1w1sRa0YhPrb
Y6CtDIqGr6eru7cnY4+JJWh7UFS8IlN/22nG5VbJNOfPh7K1utuWrud3tyM35A5MgrKspDvI6piy
S/uaV4aRYVxj8mMYJlKUqukW69Wkmq6/gxykEim5vHQs/Lcrt5vebt7k2LN5JmFGNCy/ZcJH/5gc
iv9NodFA+bEQoxFiIT2OnB+2iyivMiPCJ+P8Av/yWHNns5Qz/pAsml3li3YIy8xEvzojf+GnD7Cu
r5D2e5S1lYFXsnxmiDCNRwF1Ie2H3ipD06Qom5qI1+5XLxAwXevcMXzucjRjgUtqeIhidIHIViM0
PhsWTjRiBIYIYAROl/xPGVvgz1bCfLLoFndKCj1SYCOjPO3JEOphZalrSr+dH1OeZ12GOFpC+lgL
iIrZjwxsOQGh7767YB2EjBV09vtSk0+GwIS3UUzML8INRkT97jre6c15FNCZTYJDIxoAFedGZniN
ZuoWEqzX1T+kr5sp1pEKQyzKYYqJ5vX0EOBd28m/Qh9ECj6A83aYiOOEQPRz/Q7kJyVlSqcr03mE
u+b02/YDwqBs5emX2Vw35cdQJjywo4BBCjmufklCI03HzWx6cU+JuEmNo002Zu9lVehxCe7OOx5S
3yknpwjao07JLw8Gnz6GC/qeJGwUrjs6CVTsSaSAKFKvN2lJub5/y9pETL4iIbB/52KDYNy2VApt
7yTg1nX3pGAds/Tiwot5WhjXb47KXPfHF2sGnJOvysadnAgo/94oa7O2qpJHWRkV49G87qUf8Vqn
lOXhszbqsTfaCwJE7ckvxu/fkrUKuKwPl/pdtWrzHyYdg+d4vR/EKeFgwgHrL97rtOeqsUKNOuCD
VCi+zs217ip0WF2wdr4X8V0ZhkuWKfSWXSr/+p2L+UgOBnJqC27jEnGOxSP9hzLVElIpXA7VYHzD
77tm7AeGImWpkYeYzzhQmQ7x+YJAPNvVh/Z+GqBKqYrRfLt6a9ez7V4Phgjmef3K59pqVl/SU69M
9orIrSeZrQaWI8uAg5KoWJKsx4WH9gp2H0TtGQSS/AGbn78hi9E3lOtirJTJU4ERbA9SqSKNJ83w
5eKiTdZ5OUyEXxrG1cpZni+BiR999zjwb4QWSKbgYv7+LM6qAo3SmrJtPuUxIu66XSekOMGKBirw
e6SigF8dIuSFyyiVjm0OHuXwd90yXMtohJz3KFq6ZXlEFb/D1FxqZk+dwj1r3+FILsP40evtnPKf
dqvLS0WEybd3ZAO3/0uyzVmB9bcBVD7Io+HOvjan40XWsuREn9faZPhRUv6c6e/CJ08AjO0lFbAH
l8+ySw7pg8oe/K1lTkyhZXoT8/a0TWAd9UoB7cuO3Hbiy3sy63oXAc/hPmxMpsOwWnM12b/FHa7M
rvCC5KY/tmJpd/mjwYskcde2uV965YS2M5jW6hm+CeVIB2DYe+D9hDJAkHl0Dd/EhOS5L2QgvjtL
x4FeaysOu/hKGpSKh5vVRF7ebfI/hr912Ab0zC7haj5oDkn1Pj4261InLGrsDEAcFDmbM24YX8lF
WTwhjstjxUmV3iR/Q405BTvXJRH0dOVvCDHBhs3S/DTfTJTOyZPNEcz+xj01onO0OaA5wAlzktqA
pfa6OYs+tnX0bLL5A84E1uC6VkhrZRkmTbjHkY5I9qyClwrjV8dCUgsXShsjhRGfMN6V/onS/p0D
B0Sn5jHDNcGVZYmbTsRjf/C9E23Di17aGPjz7oQKTd050YeYvYr7nOH93RQ0Wb5tkHggB9WQ6Fug
1nWbcKdaZvgWGq5Xmng6dMtqIQ3kp9vMcbiaa0MML22qIDCC49nnPM1/wE3gp2TjR3R/aqflhWzR
LSNgRm9BkhJSDm1z2sROMPJlEyHPspy0+EUFo1h8VIDJHvJNQN42s5f/6htfiu9qp9bNON4yFt5k
X/+Ow/q0jMqVrCNA3J2kzSXdCF/ib6hPcbskxBMfkCtEsrwKOU8AT0skAU49dmtQRzFSUfiyJqlN
sqfcXmld4MSfGOSazm658+LHU53Wiv4fwN5hH7zqZRsJuO8v96ID5c6ZuT+Km4Tv1bHez+peQAQU
T2QpFhQOvBtKIhhfp69M6PpHP0isl6SExigWTZHBcp4vzN49KmS/Vfm43dc84/F+nyarNbCCXva9
k7O2yGLixmZH+9xenMcN+0vzJmmuvh9O9lpWUsihZzpK7cme5kGD95ORNXAoe95pDi402pkNNU24
+d2Tl2ahhyjy4Dk6f/WI78opw+wWtnFuamU7b16Fb2qrUanJ2o0Q/E+WfYfGAG8ZfRWbkb9aa9am
q06aMQv+WeMFtqIP91sQupFJNa4wciIJxKWS/h4XKyDnjwh6fqYViumVo0rgI0xufenlx/PmcEDw
F1k22Xjz8vr5nMzqUNPifKE+mOGCe1SMvGxUeKKuJsxm54BjOPd/2BhVqSquJgaf4Q8vEb9pPDBa
IvDlxvDbvXNoc/2LYZba6kN0r3WuYrVPGyIMozv24cgua5f+YBb0AU6/us0xpY10bPkCernLDHbI
SOAVbqJDI/fR1qHtk9jHwpUm9qIjcY7Fm5H7piT9zIMy1chBf+0D2icq+QjYtVSaELluOiOpsvsv
u4hnhQhOUd5HR6SKcJ9+x1eXRMrayP7T2QhbWN7qZHjr6PqtSqvKZzHwJ4KNRkpsl8bAsxoOib4D
zcIAUBqrXCoVQFF2hLvCUvysbgD/WCZfkTLp+pfhMgSq+ATNy4QNrgV/N4o/W9HVFSoopowKnq0C
KiyUj5mVFYU0MCc4ZQglck6Nk2QoNOARjjwTLwZ2uJt/0QXFPhAVMZ4JjYNGwU/0PilT86pvemQD
qafBNnmbIWsn7B26z+oKGvCtrTXWyR4gEk0s+x3ABx/C8DNBy4jsO5xje3bCNOpy4EdtcN1iEP+Y
AJGgRNr+/SETM5XrlaUZfMZ3O+PrjyfNI9SLeAPNecdXFtp5sadz7xPy0M93wA0HAm1EsZhq2oZr
zaVAnjLS/P6IWRCozfAqtjYF0GU6Pjgw+GHY/I4TIOUdAFJWFLbkafmeZ94i9BPp+Rk13ksN7cTy
6zMemjUDD3IIDCyS18XSdvSXy7AhCn6kCb1DYbASu6l4zkNTrIAv9Sm8VfPCaBhwPGTZnHiMAkoz
/iId1i9VMhQ7qb8e1h7bfhbhyyyOQ5i7l6RMBsWrXySqqF0/GwOujeHgQ8i5VACpZKSOwutq9y45
cTJFSluaDPVxvGaMsHD29Zz+FhK1rAJGHK43i2bgE9DIK5PilhTxSw1npCZBUUd25k9F10eotPNr
bF5ryV02JWq2D71ybYBuwKLblRSNri9zdNY/cIi/l+Jv97Ewv14nbXycwNzlZGQ+QzLAESIT109d
il1cF/5NyMEX0mqy0dhAkAKrnyTJIMGssQZaSrh8WteYlxVBV2PynbUcYxGNw7omuCxqz9Wr19Kf
pJ/aHfdVSG0L+crIzEJmXQlNYva8g4w8UQTsgcZtYK3oE/nDiTw8sxe4oVDiV/5x/I02hslNgekC
OY1m1I5lpycPDOmp2G68RFnCOaBg53wDMoMqpQOKkLlUGxHi+H80viD6l8iDkmeIQitD6drHLeK1
USu9Wa2IDA2m/h2bP6cT+foGal0B+5G3Of1HCh5TJhJ13uAcTosaBIcYmujiDm37pv9TyIWoVOng
oCLMDL0MIPDyBFuXCEWjHgtoNFDpxiv6xQQ/gR+fEBlfGOBejeZi/IBZM67BhqzzkVL8/4/BV3EI
Nuw2L1DnF3mTTCYoOkZPP1CqfnWIdOgjQyXRn02lhazoae4f6576NQrYZ+GyajEr1yLHEzL1mLin
cVrBhgHxzlozt9mo3sJhFXOT9laOkMJc0DgShK6CaEYHqcrYgF26bgj903lYzboOenl2Ki29fZSB
wjxa4vOEgHsRZKIDWRKApaocWoTDRv2jHJaTkC44onoWbuBd/0bxNiHgmquxX5UcevMU1cgpLX12
FAm3hjv0YT6hbqRiT+maXUWA/NcjICG6/Mnb0jkoY6Rk5TZnHRa+ki+tY3wb5dvD9HIRJlYvP+Vi
SSa+3NW/nzDEEsvWvbVUcg37Ba8sbEaG7PmSiyfCcmtVsUlq4PmqJP9P6srSLc3Dp1raGd9jGJQr
t/VbCmay6R6bPFr/hWzRADGr22o5dHDkEnjere9cXruAcuZ03KdtwqAQWH/5e/trQf1Fgn2vhNcP
LzVutSlK6OpK9FLkuWg+HuD68jmFLST3Xbpp8fjmtNgKSsciNSufXQTeifVnSiMeudDZlZveJIqC
fu3tmbVG0pjzGlZoFUdUKVXlINypoUleyg4xxv/qHtwgvmleJswUOqMInP9ieBBVyUDiXpwMiLVH
X2QGojwhzO1ASBoPaqtKH3pMTHoBGr74wwT8ehKp8O6HOPvpZPNhFSSPrkcz5AUwRlUqJx8iISum
kly7wE+xhOpMGNR9+xtQiWMSNI2eD0D0sz/I3vYNx8uc39JE6HfLwIlHtgVTPpC5dSQmF+kfdio9
a6tTv0X7Tk/8K825deejbMbYlVIs2hVEKGAbPGu8iMVHomDQNWd3PX8+Lza7hToAvjW5QM6refE7
hRkn+6DOJTBOyHcYr9Jxi9B5pYwzu6OJFHPZ06izgkDUdPJNN07db1oEe9PTSPz0gvntuOGJjUCs
5pw1p/xzo05NpkY1+z7HWbYKdITJv6YgafqPByqip4aHBYxIwHb4rLRu63Nt8pAGCyo8JZI/aM/i
7DOtSxCz3se/9URyk5uQhcdTny65UKOnLsTaKNocG28t3UxJuazCu4WtvncaprSJFBj3Ynnt8YSX
wLV934jXA6TW+Clgbro+CSR1U7OAeEcQ/V9p/DMB9vUT65BiY7EXS+PoNKzJEC5/DAUSVhwPERHd
OveVgewfKN0RYs8XC7IA9Il6TbyiuUrOt/bLOFyI3nI4Ei5GUN6S/CkLmlM/OTyGn9c9Mj9ZNajV
W32KpRBJ0VmcF3dDF8wfSuuCh2Hwrph0V7hFUcua1YPs5ed+etWkhdTTrja6ZZvD0/1ogZFHidYn
o+vTlXFvsKYWoFnajNGrjlrKv6NhXe8wFaHopbrmGVYNKhJnQW3wsybgNdWiKmcO9OS6NuKbMrLx
/j2fztbLbrHWBVikQqKiBNl0A94t3YMIWhTUohDSlYXsqOdScWgmn1xXQe7wzKs3W50TJqtirOW4
Ttm1kUajzBESaMeGLoEtVpi7Z/MkjFwPJXD/IyBFX+EtnJbkEaJK88S5eBzdDc8GfGQzs2uWNaNw
S1vx8yL/gfieBbZxLcH1bhmV6v0WM9L2lDDJIwG+JaKLGnDuHMWh/d+mO2xzUVWACeEnOfP8oKtn
W5xyYdUzkOWLn23+YmK1qrq0lXogycIUIqCXaIqEp+TYCet6g08x5BMxKsgya3+gNoL1YpHyi/T7
yRWX1ilAT2IDQuCXmIPUCAtfi7iZO2+64EaX2/7GpVro/9qpZ9AG51zVTSDBiMMWmgIgtXq8zYo5
DO1WSMl/pP9ZqjpRN2wJvUcpfLxIvJxmwIfdRsyCx/zoZ5FPa2a/r5tT9DfSpH83rVMa68+6jQtJ
oOxkjE8c15Ya8JWSEShiZCJEti3AaWWBATIZ2w2yvuFpfCdF7PxleiDoREbIiuHyqXs+jAcKwr7Z
T+7KfbYkaMWv6y2LjGIzbNcNmHh+muOLC7oMOE43v4gYGTyvyZIvjaTe0t1M0AtyE4tmh3AzT6bd
5jUSdv8I1flEdQTu/y4ww4jq0G15NCRuzKLOC6iS8wi2J2TOh/rwxkQEPbe1OvHIQBBLQ8B4FF0J
r+8jMI5UhWEiqgAWtt3/aUt9pdD7WCHYsjQwIHWhfbJRCvKMFB9TEYaPrmc/phUVA4VkVUndzF79
imo/Pw0noklKA8p16RfJW4GIJeUQwOj9lHG80XXbwhBA+cONVXLFvLqXNXTFfFmIkYyp1XQUdBSd
OCZtw7MZCSToDkSLH57Sd3/Tjx0C/4+NY6TXcc00YUgD5DPug1M8lSVNju0PNLzoPPSRnp3RMUHz
DQ6Lw+SeeQmlgYfWKV38SCCDtaGD6V0MEWJIwWA8ekVbfg/ITULBdW7hnn3HSM7oUZluvxmH5e9X
IH0PXuKDRFnB58no8PMYXkRRv7Dxw6hgSXbHqChF6oAD1Wi7J/WLJGvnR/GE5PwXepAKHBcdf1a+
5yg374HLDt5SvuKj5fIXTYc8+LnM0V/4GPdSwbBvKYWBk6G8UylMs2XnQ++cap34eCe3ZH/UARXK
bOfXQt2TdKGGWjnJHeIjR/m5+uTx72KbLyVa5hFzER2CqTvBC83fLWsm84eOHLsj93slq1u27VU/
o0v3lvYy0eOtyyHcSW5Kjud+rKvpDznC0U4wH4Gb91BBLdloiRxzK7tymqpcaWpdXBa500xm6GyJ
KQ6/vM5hsI5cuj5UvyvjvZ/v88rzidjPdgZn8Y5qErGeL42X9rcAKKzJnvf/vXjSwHrjoRlYhkGO
gRDWQ3v605NhF+2rqH7aJu/H24ixw14Wsvc6wX9+GyuPaWroTfT1mNa4ZJBRpFFugUC/R/mr4R3k
6V/r5yZUpLU6XePEYfukOO6q+X+7KVUFhU4yBCDXj0LHKBi7QYhcBf6itK38NEjwf3huKXtnjuQb
ihHPy8qJ+sIadjYrY5t3cgQ60f0g+TLb2mXNS4FtFeJ/qr03Rx5qIpXrpQOkB90QTzF0FGMYMMqb
+wzvWEbNOw0RSMdklo4OIY+4ErDvwJBzr8KGE1fpyPZx46RXU4Qbt1mvXv3NWLYoQhfNWuNjuGJ3
yHRNZAh40M5A7nnj7Et5LsWb4+DPvR0Im38M9jDe/heBfG/4lauGCnd1SQohIIA9DMey19mclt9v
SYsVYqZ9h02meLzevrRJd15sIHtXtYMMPFeXCWCyh/0wxBzvbgSjeshUYYgkMpeM1NgcYBGixXcl
O65rC4PIgPK1jS4pemRGakiU5bS6axW70oHjbZEZnObTYxlQkLCVa6I02a6o1uTrqHFPQjqJVpFe
q2eB+XSl1pXFRLuHcRYgN7cJEFrpliIjXzZmzXf/XVo4zdb+COBMnn9xgN/GGBB1e46JGx4jKm7Z
LWYSj84G4fsx47u6EPV9fziJ7NJtyYjiR2h0QAO/NaxXluy1REQ15HLCB7kRNjay7oNkEbUJ1OaC
aMObWLlDYZp/4+q5S8CbvXnldHOsT9aEwRZv+DGLJ8Tf0iNqiMP4Li0ewiE+VN0dBp+BB12JtclU
qrx+T5nCei9HEY4SrFNRiLFDdH+LBg6p0msdS47k2mzd2ZXpiL6fKLhL4sK3LBpwpcRMsNtW/+6S
EYarYDkY/dM4WHJgaZak/bMW/V+D0ZCIMJom+ALcTxc1oIXr5WK0cWhTg3FI+ASUmc/NjQF+YhkW
f6XXodSM/A5gClpFn+M7/ThA0tOM32wrpd0nR1fd2GapB8CrodARUSmVA09hOMBzBvL/DicQBHOd
H2/OWSfAn0ldbmvvqgEifgWompU0Gi1CVq46BXCJV5+Iqe7/DAQ5cfIv4qoVxFX/KXAxINiOzQNh
CaiF/bLrQCMj8t6sgy6K4VygfqZ1qVRZ8bKk1J8dlENCWipYXpG+zjc/HHoOHZ110gMCc+JatxTf
COyA5s2QH0tqpr66ykp4iTcI4wsyDXPh9PTJ06S1SE+vaUaRPUEMpX1bitdoqUQoPEl36RJS8vQs
7r7ZPP8QZRupleOYq8xuD6HmW+jk6notJbRsfwdRLNY9NFrU8OSsLRD1yMF4OStzmxyy3k2VcOg7
OIsRtW2vRIV9fz71XFeyVKMVz08kMOJFmeU+ACGQloHm1OE8yRNeKgX7bF1LfP4vHFX+jGrgpjXb
tt9+uaawPSLMZEm3Jx+SG/k5fs+uyw7lLkqjBhO6XbMAaeyl/8CqvkWtPSkKhxf20/dYLfTlI+qB
xKUqsgLsurzbV3N5qXacn7ues6VF2MDUbfHvC6jaqFxjRKDDgn+RsUAKKrFFaC4J305G7hWynIOR
IqEHsmFNMBi0xZWJTnMOTtkOeu/zBnebGQcnalOY8yu7wDz2OrgacruLyvuPRu8kdYwLYA0dKTeM
sdAznXG59Iuzc5LDxbEyQE4UoG/ApkL75fiLMPGFINKKQs4E2JQBCgD61ehK3+DfGcNCt/AG7ZNu
fhltmZ2LJPkFRUib5J3yoVmczy1jfl3AM8dgqbFMFSAs2qS8Auq4mLIJsAMwOsSkhgd8bNU4pDfy
e88rq5TxogUALZyirdwXreMXlky3VpnNteQNctdFEU3W3+1wnMSpIgKNGGUKw9B/+0czRnZpixCc
lyr045BNgZsDHqGLo020K7DHXVhlluQJKEw95imfkpPTtR0cnTUSKDmWMB636LIyzYZE/g+rpPtF
N4gXOyg8G78FZiMa2kSrksUr4hPeIDBqzOq2ipndQ52LQXbIJe1gLTMLqFqekILibqs0sh/Lw/3/
cBR22ySZlSfs2uBaBC6iCGT46YwzGp0bxpMn6d7q5lFfC6qtKFXyTmgHF6LxHMeUBaaZD8yLP0g+
OJTkmY2nywZAlSB3j6UkJVDTgbG0YTsd0i4tNIz3i1K9Q2vftVn/LXn0wEbThZEF7jr3bXilfFC9
/xh8yusJRHmSAOn292D0LCUlEs1lAdBmqfnzjAni9GYuPLQ5Z5Qdip8Gg+v0wU6fjiLEWLDY6ayY
dUiQ5H5aX5rrFfHlULx23KjnHnN/ASB9t6tO1x3SXYYVuvScpSz2Ni9KMwzHwe2GdssGkcOP8uxa
vZCOazD0ytbUQYgWbzRQZv9Ay3QxHXzkX/BZBiAQyS57EF0BiN1j2LCu2Qm1XPTmehxymppHK7FJ
WtGWrIedJ+41vUHeskoqrpQTpnRLPAHUvPY+8cxli1P6IdPL/14oWutk2VbzMJQTgiRKZcwn2Mu1
l0WDkffENlfbWMgKxRp7JPnuOMl9jBJCYLqbscp+Ffl4M3L2oLGvJEoh7C0JcHeReviH9WiXPQg3
c1Xi7CcHHNIYHsnt1l2nYUO8hrBwYDVOdv8Rbk/37V1b0LFSdpVI59N2ET0JngpSumCkrr8k863t
6FqYPuIbbBJD19v4btAUh2Q6GInBRMItKQpSGC+vKD1BbexgDLAOQF95KWLJeFH6p1SQ93v1zCHU
Ne6oFg51yxs6jLrsELpZHyPJnFLnjhCp2M7r4bfBFOkJMsYDBkXdWJy0raRqLwSWO3IgVA/6Uu8q
RWsgpioH4J2UdgklVv8VGttqhRmDF0vXSsAXHbJZ2/m6StFk1yBOqg/cct04v35BznOSwBV7uOQl
K/6qr1gT409psPFWHTvQ+QiFnTagj6ie1tCFPJBxVDqboCHxjxrT3fl3RaSUV7K8cDuFxg6Lp4gi
5Rr8M1fMD+/odsbofhJBhZZUe7FUz6wdCG2AB9d212n3B1/SEPxBCUKZAQQbBCn6DGHPy55Aefeb
fIooi98rj0buXiWvU6dQDGCrO4Fm8rP0Tdkl1XokodWkm7uaSqMzvS71zBkWUrSv8cK62aD2rJGM
lyLVE89fOnVbAs+e1h9h+IqnEhZcFOEhv4EX2RHZnKHDqHPXIMAvOBfuC/fk1YXpFpQoUgQkdnqF
xG/AxSpZ5s0Vt2j9PCphWMtnhbj+cvN5bSgR7SMYHiTbr+8LWhLL4K4hwkJFRha4qk+cQW4CuWEn
M4zbGACWGJ09XCkDxslyQU+dOfXL+fOGGyVE65daO95mihVYhRAmZJPxEMEzSbARnuZtjtqASd4P
+6Z3IbNobZ/mXzxea8FWum72jhkHYgMleqFOCXDkOxgl8pOu7CbqiTLx314Z8/+7hNcYL1uAT0WN
T3oTvbATSEnd35uOQrsBF/qmQPztIcShp9b/RE/H3KXnNdKYXbTWhWfnrhlVyOoaFhOwTrBjCFyX
wqCq7F7bajXBibDAwN3GTaLzL4LRqMDmBaeVTzFORNmo3YNTMllkrE5C/UHzr5Dqf0Zxgl7+UA3f
cUliw5cKIO5WS/DkbWvxzcx/faEZpJRwYr1yYVulVN87OTt5odUlZnr2kIm5l1S0nBWeGfVwsMrO
IseyYQ5efSBod0B3XS0EsanbGY7Cz97xNvanUO5zIqCfTEwMOEtLttxgveqMMVx9Mv5PsyRhT6zO
Srp1Kff8Ooodhghz88p/Rd0ajCokQj38UhxhBm3Bd9Jr7A7x+Ld+7/Y+SndCRaJZBdeZMDi3fML1
k+tbGnPGs17aKaxhpJtyDpoGi1HmRDsJQludrKTJf3o6B+O/Z684UoqcwZPHrjTwMyCDc9Fkj4Cv
tKD9OtMZ9/7/BBavzfuFd5k2rbJsJigh283/zEcIVX4EUqSo37S/ZQU3OlckkH/5MpY7p+6vuoIf
XokQIfg9233AU1N5BH0dRY0IM/BMAqhDJCrzm78Zt732j6IZAHWtDz7ovKu/7hyehdAn2tK/gLsz
fLukj/2Et62h/2QKNIMvBElYOPk13PnCsWmU4cV3YFLJfEPZfEFTLm5YB01Lr0hDzwsfJenfBayn
samXxAp+PyOMkRER0GvWxz/daEDzXy7/bRpJwlVXKDyEBBrfT7igQOVziKo8jaH1SkLVqJl+J5To
tiadRJkJic3mhyOpyJuV8t8XYi+zTHPF2teQ/zyq6xPzjD9Jdv9RFOtPRRY+xG0+f2GI2IPpwksT
qQEupKXx+H+Jnl67nVj59n9WB+/vA/rsGcxi4Rkoj3VBueZ6bXVWOsCkI+WESoKSV1wjeV3Fa2IF
YnigNG8kjcNYLgiBFCehUpycua6B6OcuJOh+bmdI7JUoan5vERf/gM/gIh03mGMsMi2+tcMZHQr7
xMEsAWGpmFxHc7P5vbAZF1x96CwkGT0hoXWjtQwIuTSvKghc+KAb0ilQ5q18RZGxO0GGRu2c1Pg7
ETeCYUV6cl3GzQehvBzCgbZGhV43zQZalnjuCoAhp6ODS1Oc7rbK/ifOjsO4i22nI4l8OR1njw2v
jHzlf4dMHU46bTWUAQhxao1KW5/pcUxVjhl/+/b2Ttprkbp36GmeJFNODBYZNGJOQKJR4Wv2xTfU
BaJUv1xyuXqUUJRHb+xufVtHjq0bAQ+ET+uhbFEOVIvSgNrKALGYdwiCtRL+YuJgIdaCD8FxzCOI
jCzIPQT9p7xUTwlBCJCvtUtbWNpLnfnn4FwVP5hm10JlAPz6uoVUlbCHt1ZE0fCFvZpunyu+eke1
p7Bpfq3n5ydDarleQefZ7ipzP8EcAm3AdF2Am+0h5mdIUiaHX3cOxteIN5GYRi1R+VA5iII25kcc
zb2nUOCWynhlLhz3oCAsQwhYROVxhB+gZdORvdnHtrKuXNrt784s/TSzX7XWDAZ0qPjGDUAFbVRX
2R/ZsyTA2h5czztkEkPMONC8LsB9sd2Y68RbDDuxgo1RcwTt6vkRkI6z7S0NtGn2JXZYh6DgnKmf
NfYp6p98VoGxMiq3rlj0kBOcuF8jdO+L6J9KnaWD/IiDE8nhgjxHdB283V8WR2OuYQgX46dJoe4F
zneCKL7jQUMUV76kcYF6Di/Qt4uByR9LA1styc+clwP4Xi982RYaKtllG060Qf3NSfHA36xC/IDm
NyiQ60Ya34ol4WZ40QhtIMhURqvrYKVHuYWqwLT4qEdfE9MM1rkAdq7c2oZHsCeal027PkccpvZg
CJzL8wWpCIl1pEb47VeSN+GDWKP8IuttCugHLaWUAV2F2VuXkVCYJs+qHV07g9roeBqaIQ0orGAu
AZfra3Jct+M/Dq07Cp4ANMvacQuv/KTWFDo1NAVcS/67RfLFV8CnzCUOED7Y1I08qHskuBfYkWfp
9a0JQeyQaz4GObIFCw4gGjKB35amAeEqkUsr8QpUFygd8aLMJcmmb3k+lC8OBeiKJp7Dp4cqZmGE
Dy2sCC0xq6E17fMu3D+lmM4nL1EYrbBt+tAt/uCFjCLvd/zYiFHXr6peJLXK6y76nmR5lxpyChx8
ENX42UPWt4SLzPt1f1Fv74P1HgueJQxJvbSw9cvC1RqiThIDy/JTCIH0XLKEJgyyK95egqxvGL6j
NUVBZRebSOnKOo0nIHBGPzNEgW2MCyKG6DEDp7Wwu/SxE8lE/vUDPQ2xB1iKvpKXT4p9LG4QV4B9
Trde9SH8lAfXosLcrxFpXQuO3RRH4MoL/viHMh74oRz/RMsk/8aDtRknfz1lqbvciYvaG+cugR16
4QWcInqpbmswvk4YERsdtJeBaekoWrCE3okObE5HGBibYEdK5PkCYsNcreaG+x5RQB3bI2MbHtGF
V65EzaeSn0yxfqSp4ItK3cAkjInDK6Empgepjnp1x6tjITbqiGlEiQC5uw30pheY/iA8GhbaMsP9
GMA2ezAkSlok1bTQvvbGERG1mnvcWpoc9ItvDGnkkWKMVINtS1qxcOUrsZtVE+DuK83gm+Old6tN
xe6ZaYLe6a0DhWU3L4Tfx7ieWdkJb8v9SyTexoeNfUkUO+s1rJfTK/M1x2V2C+UoYdnwSk8CV9yj
59FvxHEtvWfwdS6rXvjWLpwd5xlNsolse6XcwnSzM0r2iiivODQYau9FP0wa7SIXvReIBb5/zZ0j
T67zkC0jJseZ6AKjJAXf5vASzT0mYURcaleJ7G9QiJ62RBb+QbKRxKA6fnAY1bIfHzjZBTxI+IEj
MSDO3HQwQE2Cd/5KRH4UNFqS1rjAMEQQSDSb1nG7So39AwHikcKqwgofzYn/rpKB+zIrWxKuJu6V
X4huTJx+SMvSO7cOcPhCz1zNghQ/oka1CFueIxFDymHfuQlBPe4xETnbwxsxGclUO8PQ0xijuVQ3
7NKLj8yon4t1c5gmrfXKT5ok10qTNXqZoMVlZlCKkLIUGwbzBwYNDRdgJzPwFtVhDKlbE2371/ST
LlWgIMp7ZSvN9epYm1nQVEgFRfkIU4R22OfbjyumyB09ai8LFZMkvKQjDw+SPXfFYg7YgdmBnRZq
rLmJ4wy9MkVcDbIET+IdjD4WG56EXFM5rmUXXL4IfHcsAMqg9DT5yVX86WV/X6M5O2DGMb+vLJgS
KougdxcXsljnkFkXsLMcN7sGE1IH16nWZ+MOi2yUF5dnGJOZNP6FyCyLstCSq8wDur2w6sWyzCJW
l/4F0iUKSPsysS60VxNa/jRnx6gD8SbrHk4qAeleH9U5vWL7qa3JJJqIuXebxnZ5+YBhZWNPQGub
2/5pdSyO3jWU3yt2VS3Hcghh12H9/Ti0zcS5i0kVN3KWaX2MxuudFeZI9trflbvwRn1AYldbdkAA
gcOEEjelsFbhn29Bg8hBX3F3MTw5Iy3ybFJQm9zJ2JvD92meDf6PEOUZ12pk6BCNNO+5Ew0aqX8D
tTe4SrYuYakaDcybEdhBD5q2ZOz+wyrepx1DcTGE/LKjBNkTkE/1mDf6iq4UsJwEZJMfI/ZJKOCf
i3pLHCYEwDEKP8/qFFPyaM/l1RyOWZ+hqFBk2r+tG1+8VErAAkT/3BSKUf6S9t+kYHPfkFAvrQSR
Iq1H28e/3NrLerqKHSEB1DUVLug7gWWk5fPe7e7WcWvXVuD81Dl+A+jvgnRnPl4TCKHdov/+U4rD
YthIQtT3sSu6SRBwrst2dsZxzuYtep8NZhkDHciho9tt7vI23+Z1clXrE3CIvhlLAoMY8YAvFgiW
Gg4na/SKddzkFn6HhpMhesQvDqFsjGkSih1dz3P36OElPIb3jm28biRoybE6o2gYvx5889Uz/g/0
m6hZXXseLl++53fBTOsWvr2IuAdBcKOtNpcFgBCerqRKzvJU3/s1ZoMmiDhIp7psSFiWBGCcQRDx
NZLwOd1M+JaaItiEZStrracZFyuxoyf12/DCatveumROEY9oQ5b6qEsLwuZwbnu7mOeG9VOoXqJP
L8uwAxRuFpS6Uc8vyqGCdx+agEStFhyj4zh7gENl2uqVoJRrV9Bqy9vuu2F1ubM2KLiq6yciUdBV
+eubzYUAHRE6p6s0CIBWYoCJsUdc3PBnYkeDJSdb8mT7vg9WOuFEAKjBF992AcOoBSdJ70dbxHHy
gqdfu4aZQTMostQHhFN7bZiRpaJj4VVn7iSzSFt2H3A6B7yvzxGqffUnubhN4sYEQhurT/baN4vZ
PkgNHWSWzBvesFodc9nYx5ZKxTcy7OH4/vS3uFkxnN3uTxI3y3bHFzaCHoMlZ0kclvhLC6nMiRzV
esDd6ssVrMmKcRvbChQlV+LoLemZmRQsnSaBUtBI2CHpbO9o5WP+NVbM5JD9tKY11Zbvw0DStcng
b4NZPLYOxQ7XA/m43hbqDHKUcorC9jxFPHbXGgYJ1s7pCikCIR3fpv0Rih1QSLEnycn5HjlE71nJ
2w015GMcJwtR9lte3RNyj5mIwTElM/pwYIc16qTo5bznmP5OO42dZQasdPP/gzRDXQQ4tjDLKVnV
TEZMRc0hGt/9SnBT5+AT4cuHAfJDI5IDFLq5ylQRjvGOfPeG6b6n+B+Gz4JfWZqjNbMnTpWiG2YX
IDHSBxhxFfpYd9lm4MTwfnvmszKqXDQmQfrwrJJBF3ABP6jo4PRR9foXUXirAT7Nk77/k48yvZZs
m6xRqZO4MLtMBGZIbbA9fRlEjcRWO9ZSwaJFZVn24taPJ2Gz1dwT247tcqTSwhfMW56gsqj38C2s
GuynOBWwCUYr/NBoKwVWLcBWBXogguwJ26E83t5aY+fyoMsfaUNByQ2Ddr0CB2srMFnDfD7Owyqq
gQfW4jKv7st6scs1ITDzkHFWrgvaj6cjm9/wbceD8TtDNTRHoQJMZNPPTkAuyqKo0gTzLZsOfWDv
v6xyWCNxgo8iGWgD0WFOP4HYhGiHwikPTdkdSOPplOa15wFKoa8GYiQGJrdjcDM2Z7GqEYNKx8Ja
cAN7hlwUZG/5+PahgQpRnshExt7J/DNXmfGW9ZcNL8/mSd0NRRe6sLgTVVOA2LMsVAN9e1MSRp1q
qpsfMARiYXvOBa1CsOBn8IRJ7a9pOwJf2qF2VGf0QBfhJBsIfT1CcCVU3xCoppDODZiXgJ/IhdoD
gn26sQ91x0vFgLtCGWukIcYnxv9R0r4lT4Sn8dUbkzUVuVzsYsw7km+JPcS8PWymUgQIqBsqE+Cu
SC5o/D+wy1VSQ7WwR9rnkTi6AGiLm0ogyAKSXpHe9aSx0liI2kaAVHRYdhc+cAOvqIugJTiPzOMI
LdcFyael8cKIPb3yKtHHrSB7e3YjOTcjx3KRAF3xNDkQcYMakqyo9xdH3o/oFy6W2ZY/pO8nUEUj
E0jHKuPIQseEhXT0t9Wregx2GfhDSE7gk6r9x8srcQNAJGkZf7Wejz4BVfzkmbu/IvdhEo7c253v
mnE7wvWgtEDCLER08MPfnB7gIGU079jCGTPny3dn2ib/hGt99n7WXlqVeNJh2S+jFwFj39jHz+gT
38l0kGtGsbdkyPLqhDYyKy1kw2GDijqWY7GnGpwa+ExTbmdka805N5RdIxbSb7pJDCND4BjFxcyd
pmYgzNDwz3xdGwwHkj+JE1wjopAI/8GrFcZw7X5C0k0DQnFrDwj75e9wissTOBoTVxI6ABU/RLiW
nEoTwGUA1koFbdKnnVX6PE9zJmxZ3qZayznrgLmVfkDsR1zdqPtyH/rUJ2eAQ56VCcZYmzlFYIm5
jg/IgG1FYxkaw/alV69XUgjfRLSfAPZyd5HCH8az9Tqo6YtAXaQ4d5VXpb2LdGEWOFkoaag+SFaS
SAidGL01Ez5UrYWfodwJESWV0my5oCRXlr7LJR3X6jDnD4GDs8rrxtj2jcDvzTDPI7ntt+5PqVWt
QIXqTSoH7stdTfUUWKHTClgNDZ4g01eTLJcl2IL/vYr5hv9l/jDu7i/44oi2tlO7LFrq08YjZ6r/
O8cARCTW/U+Ewqa2cOlsfcHJ/LZtn5J0fyPvth2dgu/tOPQXdRQD1BX90i1MhLqf+1oItaPUkaeX
vpCyc0/UtO4mXvnfEHUtTTEs22AK/Ya/ilYpyilCVec4CVapxgTvKhDf2uNatEaRpCIoQXzs6wen
7gefqrOl9ptn94a5Yh4AHeinSYnjwr0s2hnyBlrumkKxrdWUQCZMLzVNnHWKTQRei63YfSgDheQf
jMyuvl69lBOHoyT18BDi+xTgSGQdblzabm8+CA75W2UsvxDfmOGB0xF1lkB2NsOeY2w0neajAjLJ
gU5ZTvgqMeWM3eUyILgSPfWB0/oPEmUgIqdj5UNsEq9LavgJHSr3HnEXpcCI3UtgXKcVJrA0OCnt
n0Ai4+IGl09yTD6jeM3uAq9QbXxwBDfflieATHtroblTIWOWHG+/H/wZzKzali7Gkj45Anh485bw
hkOyoTg8Svb9od80oQvvxwOTXQioC/Sc5+oRLHgfAirGk8keHlz72yEq/itj/Xx337yKAOa8FPAM
MIyorBCnIbd2odbxreVSqOwLTuhhP0r3VOibew+oZpGYWXHTUO1gVfBpbGHsl1Eoewo4VYXPB11u
cOL6VrN6B8RXokoDpsZ66vvAqgpcWdw/wBfCjL1iuWJU/cnOVLvWZ76WNxpfBIQu7T/dBo79wGfm
ppRpWhxIC3C90LcluI8WL4ChnNdGGEV043D3jm0xSNQ7T57sSdEjIpKmKZJDT1gw2Y+geYVVtqgs
Z5wWpsfAArScUWz2t6Dbh/Qvee0dxfDJITv8WFOvocny1zRC5sAWKpxjMRu+QLdHpd6M5UDfTpOB
hQ72JpuoQHLdavo4sUT02PRjgOnOvt5uUeQz3JgV1Z13oAWjfBxLXFEzL19G+8wmIbAtfVMFBJ2I
vozIqY2hJEBEDZprEryHrmVum1e96egyATolUQw3Q1T8mTB6xQ2J09bl1FWHXZcMeZDLJbIt2bf5
sfBfqFLT9zhoAEM6T+LKTB0rpyw3muv0nMCxTRKrLRIsTYYszUjXvfcgtlfVw9oMvHLyPI40V5Ok
DrT7DQztYWCSj6ktsuFOnt4BecEKxWqUOFoUhqBT9y0VsQ8pBwg2iB6EYhKN4J7ilf5ICRXp/9by
Hp6jjQ1olZj5kiHzVraW8hv9pfd3Eac+Er/xoyV6kvfc0KQxwU+Xpg4lqhLVUYFrS1TMuMv2SnHN
oyaG87zCqCQnJlxcxooJ5MkQX4B1aBOTzonXB6sjat+1eRyLMzo+ToeJ+nhV3JxHz6Wpc+pyRaQ5
nqummWvOP9Mls8kqkkNHROwwnO20uDcCXHkIfszvnYKZ6WYkq4kn7p1kNDNrJN7KAlB/0BDO3dK9
EsW6kLgH1f0g8WDGozxPzOxkdsbtzp1b3UJ7wcp0My1v0VQScaZa+k4ohLehsAAS8+FV795m4s9N
R2SpqtMoEnPupm4Y2R5onfUwjcfpo2UeGSV34HpaY9mu1+2ZmlAM0dwtCiEZEYMHRpyLb4gd0K7X
gMvrlE4SLQ8je7GnnxRqH2SgeJ6QcjQWx4KZfAyOeEEmkdQBr69BEUGqGEkhg7SrVx/VaN94oCuf
VVH1Tk6eOFgp7+qW+6LdcO50gHsOMrwqNcSOuy/rG5ucOa4ZiDlM/Y2ldyXQF0pr8OhsAtNBlNeI
FKkCjpMIV/lMEJxLjdGFrPVYCHnb4csrnOe96FtZq+RxMZc8xtDuE1WDDEnsvUkn/oJgV5ZPIC/2
yAd3G/zz8tKb1aZtv4o55FUmFWazwvx/c+aa/g6Z0Jm6GZYX2BoSv61Du8wzAAXeVHfmy3o0du2p
Xmj1iQNaOuDw386d8CgXa1oPautj/BhChx0o+MUHC11lRpLXUV+X22t6giqPq3FlnQUZUBrKe680
g8HsKYePytvV4XLEuWhaBiK1i7ErCqpsBz1c5qweHSEZC/eMZFfuhWJtf17k9yHPKsPSIYhdl7Uo
Lxqavoc8TgCrVqooEDw4Wu+xy01sAg8G/UAenwGAU94TQaCR/WZfp+YAs//03BaW0LSOJABy9fj5
PNt38rAtY1YDrGm19Br1jY2vOzaqFquC0IKLBmoJ7fusjgxXQLh6POhIvv7ldVBu4peQO0CE6mCQ
lDml9manUdm7JPJGA40TJCgLb70YHq6tsbG0YFpxjnKj2HxdlCvGfBTsMnCxT07d3ht9TMeVHpGg
zvvsKCGJozdzrcq5glMNiTfZ5+TVYZ6yY4v4AQHw9oUzLrVc2pgxHJLWsK6Dp61BMZ+OgZilyQq5
gN1WolClus5MBmaMG9cB6VkD6vCEEmY1CrDmNyyhR62Sqzw5kUvjl5MkRFM4khktpaPZAHdE75h1
YRnFmjWHrA9n69kPazWT/iuM/dru1xhhwYvFzQdzGMYr4CEGvJ0Hs2jqE6I/y+cy1IXXb168+vGJ
Ooxi2qEoM301oCjJ3244D8urZngGkHRN3+ylqU4Ee7zfGFhpTJJZalwkYUWdzvLHE5sf8gPR1vSG
F9CNJxaaUNTbX6eo2XEI+vKtL+lAEBXMKcYzYkAh2jP5BVZmigckkrRxfjbL97bS1K6/1PIEjdrU
gjMSSv8QEtlN+R8E6L85Ql6DrMcbWJqGFjFGQGLmVEUYysExLplrcU3M7HbnaTOAkeeLRTD59qZA
ycBkmXDgCCLvWoSt7oZvu66eDpS72O/fl6nrku/xqJpNAZl7sDhp3Zn4ZGifQRsfBlYpxgaZFPS/
ffANbhc2jHjEA361UbIeAqHUWjrX0h4thm6GiiLO5xm1OdQUNCgifUZOn3eVRxZ8hTqYMhbLPCoQ
XYORWnbUaT7FpEVfh99lDFHu7pf9aqpegsPcfOZHrgVxY0Y4C8YeWBOqRHQZ4J67nHMrAmlZ1yW/
EF+zVPtrzmrIECo8VweQSNYGZg3ApukVdP6SX8BtnRN8h/2VshiUFp1P7cGyVuiiFj5sTCUIFuSI
SxaLMPVcIQ0737EDUwmLSXYyHQfIcVzep8knvJTjn0NPalQks3DxOkpIHUoenlG5k62Bri/g7fVy
Nq0nEdN/iYWIW3V3W+gWGNyvjJsx010ErNwvcBae/Ff7M4F1dTMLUJUzb7M3cUwgXfL/Jb3guwGx
1zkqC+K0LNwZnVfeBYwi7xsgATdrGUwNEOGcSS65fuPIqO3bbwHjmsXbA5rXzPN9JLk10CSU+lRf
4loeyn2jPOhgOdze9cZG/sO3ExnTjD0JbMV07wPp8SVR5X52Kz/S+uPbc88JN+d+Vsh/46/oHGNR
ew8HomXKPQ5FuSeyMGBkvvOH7MYwje/iSpJuDvJZGaJnmDVedIGdBH2C97fif9W+1nKI8LDe6y0v
mGKovtSDolPMvEGYAU4CWVfPrvUhyWk32QHG8VQzM7ym+w1zPo3WnAMA0T2SKqh25kn3GpHZG3Ns
OOqM/9O5rog7/eNvAwrpSFuwT63yf5uBXoJKjtiKxXkOXjV7ffSmeTjauM/kGo2gwkLY4xnpf9wB
F4TInvCoq6ILYQ6hA7Lhz6WqaURanXBI75WGkAZpUwHuk7lrwrDzvsrxwaW9sotpc5zH5UEWFMcb
/raiThfKq4+LjHxgLN+KoEQy2xGonsuhenJOhyn7n+DQrsVozXywv2xC8N/AA9oqB3ouXcsH3hSX
pmIRHxnKUwFAMEYmP3HYCQCkjpSpC9kycOTdtfZ+nf96I/2adcxvblwsH1rKKpO2+Y2hhuEShz1L
3IZHdBcoIxQMLWWe4MCqViOudokHHOxL9H3+rHjPeRl20K6p9+0l9GYQMN/LJVu041Xt3k6Prkt1
mNsnC2DPW8N3O6W2Lemgwb3HOpi23YatzMC9brbjV4DcV3tVLIwOQK3OW4jLpBRMTueOLq/ZPyXZ
FNCullZ047tv2DzTv0qL2/kIJkMl4NFMmJNksFq03W1LCAVOwjxw6FC0bYCUKhIMI0Qz3kXi66Hm
8O7qNoaSnvejBjnspZqIKLAdvNR1WRtIsldHBr7g687rxK2JcTDrU0fokqJCkbkVgpgxqOgFMOJY
KORU+FAgXPZLqF2lt51BLwMTPA3AOpEWtDzoHigyHdVTB8Z2HJzjb6o2cmJ0AcQnmS/Lp3kVkZf1
7BUzPwAELNIQrt0iFLvdAk/bssL6Va2vaz7t5MLCyM3Avt5S6vNTnWfcLUC5R5XJmzq33rigrivb
IWcQv2cGzl/ZC7ZInItctGybjr6bohVDLES4HyRrLkXzuMruAMlr8ehotHbpgZEPZtPCTGMjE3MB
3Gj3h6QQRYxVoUaB4OYfjPbsPsVoG4t8XX3b6p6U6KC6F18afHAvYvCKnTGMGGCUJhgRElS0veX8
PVtoRXiOTkNoClXfikgQIN2Z4Hr7toG9t1yUdWXcq7zbQrobJoqqExIpegNc2a93PfawVqVYtMus
8kB5SsKK89PAAtsX6zKlzNMJT6eF7ZAf5U8wq6xVl03BZw5Pu11EO9RARXsY9alOGMy6HlpPql12
ehK8UjOwQ9SsUvG+fRGK7Th0ocuC5E7is62/bZ4H6fl9gSRIYC3IvlaijbMMeutrYSQTi2nKSlS+
43pioAQEdMBz8GY451U4ZIdgY+aX7JXSlIVm9cBHyHs0DYmj7yZukf19i+YOyRzah/L7A9286tb4
ITR+BPkn1xid3wo1LSRkxOohlXBce1KYDoHzkpe0mUeLjVvEm58OD8XdJ3AV/0qg+JrroYYtDm48
SVb0ijGCNCTJ33O6PnUzQmdkPElC5Pm8l4HPygCzKQQSX0huNOzB/4YSgOx2t+VpEp5DIpyRLWfk
CguT3+W6NFyfud3EJlp2cL3+v9PxfDFUW/kOe76JHkNs6VFl2OVqExoJra/drJG7f7qjkgD51Np4
drZtbWzkheRLIs3s6Q6maKBlkwtFEdC3GtW2cBVdghQJhyD5aVgIVs5N1+ku5A1mVNjM5xFwOoCt
NXQKsAxX4y7NAqDonCYdAzs9KI6W5c6RyD1ov80zdvTBDDCcc2iR2Npnew9i8lMy9PEndiISARze
z0KDz3LCv8V75XIpJ7uF+dNq0SlhkY/JRGo0z3AtktQhQdIbyOkblTHdzIq9abEzaUSQWChRN1DS
TnzFttZ9Ac7M+djFDojQDup0E8LK0suySfJiVzgPiusJXM9lmplfJvuvG5xeNA4avF1tuU7wZ2/I
aTz0S2QvmeCoVAAtPCWhwD6cfvjcChNIvAMsyYwQ+ioD+AT1guPz/c1GmN0qg6QPqyIIbvdodKzC
vnIw6IQsWxSwjzX6oEb/cStfyhHrUneRiGFiXGrHE0y+JiGhxqV3GfVHCkxQkVHl9XvC0j33q0mN
ek9+SzSWqG7BGmYQV72I9Vp0FLrpPQUk3Ap//T0AiUbvShXnq+74CrnyLhkkQxz6yvYhZAmtKWgQ
FbbS+nYG/wYxornA2KxSpt5I4rN0nXtGu0z4Yxa1iH9IkiejmkPhtHrObolFnfDsBEWTVehATicB
Ic0zeqeid7Ww6eiPNHfq8SIkaUu/AbYWYoy/kB9TbhBi0lqTxwgpGuHwhPHhzRiQ33633s79BAp/
Yvvc8t1i52iV7F84MvyBYbIvwONqa+j+USLQGIRNU+9zNCxwUxOqhhch+BjXaOdBrksojfdufq0O
ljdQHaNCpiAXtG+JaKMoFVoKKAdB3ES2Zzsrq1GlNFLMN/RW7NKyh6N60W1IMpJ96UIpDTZ94FRo
sq6iTwOtijK7SzaTpiyKsmxdrjmDf8XTmXcTnOZnEIu7dNZKJXUg85YU5OfKGQ5bpIl5c1G40Px1
M5tH6bfBBnNdOVH9TaPosz9AwQQ7JbGq1faOxW9cFcWGy6Tjs+2v0+rXJdM/3JYhjKFdlWYy0nRO
47V3FU4Wjh8bucSYnRxI3zT8ExKpg/tpS1FTYdK52ZXL9tqu50zRpLyWzWrrcXtWeqemEoD1BhmH
VxVLBLIFNEHlnSpBrUBru+PnHSyeUAAb1V5/IlNrq+2/zG4kooRzsdKjRfuA0i4SxuHeYHV3nabd
Dhk58r8+PT5rkcVgEqrFKqBEkxWqHNE+KfVMMJXKNlkRPjdXojhwoSIuSbmwgRkzqUfxbloGpKYG
fUp/o4M2WfKqhTsf2Gr/mLyydls/gDLXLGpoeWz10YhKDYTSa9mBjRIhZs6yx3vtdcObvoDdEcob
x4zonw6eyUBJSfcxrPl5NNtcgXFJJ+skKu7db/93yfk96t3PMbq9EgfkWLrKXzT5mk7y6qRve40Z
SEDw9BaT3GWl9Fz9fGgN20yt5mOo6aPLw/6k1nRV8LfMml5lGQhSWkRb6oagqb6oHLgcSuZnOYyT
9Fchj1VzOVmTfAtUYJsehjWcX9mu22AuuSf5gaQnCCGhvES5cVfV24prKKnJRDTFV2+3ucJE96nr
xi/tCEYM024CTAUidFRfTCiPW0dwqcfpcPKpOS0ZuTqoHB45pdF7MNbtdgaCmf4gmPf8fPAwv56Z
LyvVvM6pJzA5jiYAQIzZw8oDYknB6PG843vQslzwa7wKi2ly22QdAB+Ri/HeUKqsX27vq+2Mazi7
dQnVwALW/O541UZ0U2/XHUdW0pG6bX5hCo+IJckPjloKEDlM+7YIdSB3ktbRFoFLOdettvHxSBac
WIY52BjQq4wzfOH+4y4R/0j+JVeKTlfYrr3/HLGzHQOhmcGqCCzWm2KC5qejIJ0ZMJjy1e80NOL9
bYs+006oZMtAgc1KciHj63wi61F4N+z4ogCNhFCOomXOqvEeVbHpE0MMvXko1e+H6NjzInulW5xf
txoQh9IjKnOZYkdf31wJ40J03XLvccJun4fTDd7Sj2U6mQ2AF4xwjfnm/+VaYVBQxB+sEfDyqfAT
RQ7q+PkwsVE0KEGuUhhvC1JHbVkRnlV9B1Okj6gnaklzXrhc/leIRVp8MX6cqvqg9kXVuK+FGwa2
huBWL5CBfwXVmKenPLl8UbfndtrLg3mDD27SqB5gOBKx3Np6YxjS4RY0+DT1Vvlay+Fi+B0ipkMt
74CZuuAQ+3sC9TgblMJT9/J62D61hPy9g4QrxVntHz/7B/M+EwUn5Jxu49LrvITcqLAbrtmljmc5
s7zGVQrQjEKTPPzhtRtd2kwfO/fuh2Q/UIn4xyLg4zFwFVc95imgbWRU2zGF2hvxDmCUnliJFN6l
1zhbsBXo75ijxeDDo0+FPgEk9qVWdly0qZ66ka1LmGPAe/Izq9TCXn8OkZxXi+USR86Gs4tlxeGh
FVVsZDZ4lf1C+2dnn763Y+Oa6FTE/nA91aXc8CKFTDSDRAHal5NB7c4lTvZc0pUbaO2osJkeEhYD
2qjGu+dWgHAkFEMNLypvmCPXgzgYJCpptAdcX4ZTW/ExqdXhbChho9AqHPDWgyLvsdYaUSoHxf3t
5G94/gex8HasWfrH2Aj4CuYyJzzncxl6j0dK2mwIShXYgWTSyVzY1oTtEJBRImN8+YNYNaqSltBR
mKLyBdNa6aByF1rlHkJw2fECQ4i6oY1wdW2+qU4XL1LnNhKKIIH7Pr1c+U/NtBBeLDhdcPbRf6ug
h8am9zflGYjszWgw56ySMGYGu68Q/FEVILprfksMRDjAzV3TTXDzYuP5KEWeirq672qhOAA+ZskG
hlS+P6E6mZnIBw03wKZsL4UgCkff6P0DJtWdWcjIsMLgdljqSxx+x9r8rKSYfMB0kqdJ4k7CE6RB
eDbl+nL1/slGBvVh5gs6Z9z+WfDoU8RU4j96VOye29skA9Hwyil0J2vqtky0J2hAVs2m+mo0N6y9
V8PD3QovBxA5r8G6ue+LeYjwLZhC0JPzVTKHL3Rlt0RtJFFqVEw13NgY0uWMemvJyw7VX27VOX8G
jFt6I0FSl+lo13s5+RlsHf1KgRnxp646T/rTspOE6ZGSpKss7Lox6H6P25VWb+HS5PuRWBKoPsUH
6A1MrSEmWluJRZFYbUpR3qjUV7vNY+EMzALKvAMMUltMQc25og6CCDjWu2rU/emaZNpvEbrHZ2xs
wRXpmDm/HYJfa0Y61ChobbVykaXKYCySSVWxY3FslQK+oWsWbtpPIro+xSSgpF6cqdRDKWl+PK68
zP3iHEy8dvGNkNgNKuv3vMp4PnxPTlT6aFM8g97T7f0FPscSsbyh85Q8we3Z16DpHGifrA43SFq2
XgQft0P4A5iYeT5UFyQur67g6M6pitLtyMACZGUSzpldB99pUH0Ymx8kOelaljLP7pwHqRcC3qx1
8T59Vo/GQUk8vaFgpP/SV4D5n8p/RrylxGks0bv7NDegRIrOVPsNiOqjojpsVkzcVa/qF2mJsVWm
RBYlKp86UWg3UkhI+xXVdMVxm6bRtBl3mXrzEUwbkBYNv4JXFQc3t65Ahvdn6iCnhtkfl6l52dSN
hWvcWMI8qkzfpnASkE5S7pWQ3epQ41gM5hAo2aukSR7lVhFxPSF5uLPyql1iQ4FMsErPXKhNTIlG
TUko4n2Gm+C9oeXaeKaf1PAIYoKfiIEFAcDqIkjzL61RJFUYk1HROVXLtBoBYoWpJ0jjyn+7D/1z
ckh3xHGJ5pa/H7eUMCkP8OsRqwTugVL7xs/pR9omOlOnMhan4A5V79+stOqGGzD2rLe/HuVzWQha
XxjTbfX3G6V//78KRsHHVb6rmJAUXoAgkqp94CTfuJXUPgh4H6gVAbJAE77p9Qj3RgqcJCyH7ESV
lhQ2NUAKA7szjt5AhpP9RDD3W1Sp7JJzO+eu9Qc5wToOIB8V//A2byE51drMKS9MkNp3gnRTOe4r
uj9oxTkZIaC8vJXGh1LLwVNAnYmtERfyUcDgD5esT1LccndeYZM06yJsstq187CCbr3Xa7JScFrJ
PYiCCdSoGwaNdhHJUXwNp1fmnC3LvkhgY1yFpAVxnuPhdzNDFmkYYqy5tePA/LUNsySTy8g5MLTR
/R6HtA/mTxdwu0IjrvxXiQgwBxp6YKZHt0BdTqO4qGa8E7Gb6r6D1wNScHNiYN0BZcqJGwpvu4xh
BYZcGPcNriPyK+FpARPzeyKaqSQTkeW013CQOG+m8YbhWsyqk+C3TG8sbnN9sKhKv9nLc7V6NFVQ
fX++uJEazIeYGUQrjRQHSabDliLDAcKalx4Y+FecEqHKemSLn8ojiC1uH0K1Vs9kozNFyWuF6sMW
pWtCNVbb+vu5WfedNnal34PDrDdV+rnIMhf4N8MlA6sIHLC1Oe/w8NXC+r04Xpl0SglfNHPuHuza
zjDIUcSBWSDt90KUvc+AaMBQjNEP9GtMUeZSCwaUBlrlmZMTTw3rn7+/Shlx/QnM+woUcldvoDae
1ZJGO97YMNusc3oEvXeMXpHY5s5deeKQQD45DqUoHTQff91zATDQDwOXZ8h38f4jQDWDNH63mFBm
Q+HcdhSatpfVxGfMIMxlglIauZbRdDqYdzoRQEoQBxXlde0KEraOiYhNHNlKZU9+s9j0Rzxvm0ve
AnL+lGNtH0IQGd1rF361JgwglWhv08eytZREeh2r0SQoLPnoKTCf8wXfvG0YuhbrPCFudyJY6/31
yzoaXl5cBfbH0MvEpnuDVzhYvJCm3/n8RVp91hf9WM3VVFxBf6kpOI9KBJ8btvHvMLcDaKz4uoyH
ri15ABg2y4BgnqfxFluiTynmZMELVvk8Bxz8d1geed+v9pePc/o1gdyDBMqATM218f7KnxeIBaX9
2Vzpmi9WSCZZYRR5O/0IriSvWBGx3BrVeHGA0CGc++Bk8l9zMViggrhletxIHyUSwFQeOgviG0Fy
r8eIdD5cojpNk0QT8SVv2JDIVqeBde8RBOyNBn33UQhIB8pTWwqUEgiKAevBnqBgRv2kzxuDRmil
8rQDgu/DxsHBRPZoDiAu8ZmEcpBqVUZMfbVX0ivB4DhEWsTXzpT2YVinucCvuLAel4xYJjltCLTu
YRUI8za4nXG2ZhgNPIchy/GgSm6Fscv0wYpDNrbQL+Nm3wCTGimUBJbRFRki7gQVR9B/M74ypX60
VZi2Zd8+QMX8jnr7T14OM+BUrmpoO6W/cZhn/6WgLltAOBXJpQra35/sAUjj9ap/UVQ2VVdaCN1m
cOmuWongSI2meiQIU8n3D9n/OqN9yA+SAL6PByQOfDE8c0LXptFQNazjp0gaJxVk3ihj4IqPTJ7j
y5v0EeKNE50xTpPIEoxWfOn3z0byOTg0Ppylvml6jRYvHckr+x6HU0zJXWN9czn5r04gypGUpKTB
5R02HWaypaIeoz2Gka2tJp2tI+SSIJQfbnS222FOVS/1p6thsF2lkfENwArBJpGvzD+BmtFPMABy
KTFvH9LvqG/nWi7PxCrPcj18Uf90dijECn8F7xibb/cYowSxd9dEPlTUXVnHyUPK1V+aCNxz26cV
s0g6amqWBS/SoK1N7fvV9oM7HIgOFC0gLOGgefQz2FI7CSVLD3g3pd3BjZpshstqficYjA7cN6p3
yH9EE+bo5v5LTHftvZ93ZVc0qE3g8VntF29+Do+2Yht43D9nQNBZA8pAdTKFeZGyp1Hg3yoylotx
X7S/bURuv4YIf6CgIPxxhLQ5o2BNoMKE0OjnXvMKozXlb/Q/LDghlSpF1xXuOpK+7RqClcyymm8h
w/+a0BgwAnEDAPQPy0AFuRkue3wr3Dzg7Cfp//P4+bEJNGA/3TIIeLzyAEtWRtPjXipl0BBRzQUe
7Dh/Rw9iaiK7G8wIVHl1fg9YPWdDPyXrdp1/+jIYIxqkWTplSbSj13ATgIfmMUD9dBHvvUvK0/lW
8S6LpZCRQdbBQav2orjX198v6O7DyS7Nr16Mse6vo7+8J0DIC63avd7E3aerEhusYy0QPXuG7Egi
0hToIT00xHsghB8fQilqqsyMw0yVVnUg/alIYf8/9NfsLvHwDKrBF2Gs8JlMHhQE1ahCVk2KLvP+
ILIz0L4chvctkiK+01KX3q52W2EefHbzKBpscDRxEKC7Nzt1iLwwqSeP9eU1d6OZeBOJ7KEKZ5MO
COkbIn+0FTf1R29IMQ1AdBqtbjwzUj9z9LUWiFtseZXdErA8AiwlS2b2HnRRvLq1fkugaeaATMXQ
XC4BHdKz41LMskRAp5511QGy1SEc3JKXPDMlirOsBV/v2VpdwzN+1OMvc8ytLARdj6WYTgAfTwzq
RNu5FcHQI0Dfug0EPN3Agezu2mFFSIn5QPs/yp7JUJ02+QBguSF/kPHIS2n66mpDxu15oc/nrSIB
SxmQdqZKuhJgZmkBfdZlEaQtbvjcd8rgQVAhQhGwZFb+D6/1pMwpmKRs+jK0iXjlkschwulzFgfm
Yhcv7R3N3v+KIjgVX8kvbgFSOKLvB6eskhz40zbP1OK14rQfhhL+t4ytcBajPhVIXsfGttPnM3gD
uwmLXlm+d492qChqCO4aGZm6l8G/lt/iFdkyLj6rQ0VKW3EcrvIQ4KTjcfbZSBDh9opP//qETx9+
/C+vQdGtrwB9vIccTYtgWKU7JbC1LeM6kH5baKI/M3QTeYYZObJrs8sdf5TXXq7RARgjyboINF2s
R1AXRsmrPb5nCjUg7p8aG+KYk1NFM4E/mEJiHkHqOo/JDzxLXzRFEOBimcJOw9bQBGRFPNe/aXk2
Tmyd25kEUWVY1iLkJI8vgL3dxFj2pduwK+LmB3xHnbTHq3fz8UyaDhhYUzXSY5ticmIfoxexYy+5
yrDeZmB8iGxlgSfuZ+zNEbb/bkXUHPtBFVn86UUQ3220Qgan7TnKV2D+wI07mXHeO/XQmVYvOvid
LkKH6Pf3kreKh4Yk8/cpHx8iPDR9sb45ezw0+rPwKSo4l/GS29Cb/xiU3n38d/rCZnRLs4rx50iK
CQq+8vRjrKJQZ1JTDMximadeZBhjmEg7qkaNf/Nh64XSUYpy2KvzvvZCwBGk5NbYHefByk1ZXOB1
EVmCYF63ce9PwU2kJhiz1HQpxwL9fM01jOk2CDAlz3pgrZ72qh4R/lBOj13+oc7baDgbId0HOEA0
nKxWO4XyPQQOOgN5ChV2VuzK8dQTwyFvW//o4cQRX8FQfgqjr41a1bmNFylBsM6l3jKAP6U36vMr
+F7UsyCIuFa3Gxmg7wG/AG1I4W/T8SKoEzf2F/Dwm7Ppg04MoguqhMRwOfi619fvli14lESM7rXf
fQJXYI4FYf/bKRERzYhOLufXmHmy2ElE4LShYdCBBhL/Jsj6OMOX1+iYgTfafwgdB+IWhLHhaSav
jkVHPUVDI0aPriiuByQyvEW2Bg9kaLnP1MqFOSv/TWS8AvEj6aYHWgTHgEC6L2O3UnUsY1l9Tgdd
vyFeTjap+V0ypxyPsRUJjHnU3RNTQobC4Y3ydfCCPi9oLvS1ok3hmrhokw0mADnknENh4BS/wGgU
RJ7M0twnYs46xB0Bppsy01TT+9D5cU5lXvmjKdRegJ39Hpfg3YxJ6xAFNY5QBqcd6csT+tiTk0BW
CwaXBcKDOqbsniY8fw49cv4w6c66LJY/qxvXDHlSsusX17wDmb96XpLqRnkf/NmASETw/5xiw0VW
foyfriYwH32841HgFYh+8NxK5exrVaODpGhtEHDBJP/BEDkxUowbLzKXMvvHhjwfrQf8nvucw0XP
VBHf+zc0R7tEOdjrv9JneHdSaKyGkk8fJsbkjydjG32kt/hVNVEn+YvRLWhMkom7ypXTH1nwgHCh
ovUxqTvfhw36g6J6t5cq14f6BVdsUdrOjT5UAi6ZW2LMhzSXjVC6nN6ioBtHh31kW1M8MeH/Xbxa
MTMINiAZNLUFfFveCgADWlbSgPZS8t6UoXKroY/HNj0tGB7M+KCLDBWQlj9BQNhjh/6RJ8WkQSMR
CGr3AUpyS0whSTSi9WTLfL7BJm7u/6ogYTvKSIFXRpvee/PzWMgjIn2j/mHdSlJPpylACh7BIxK0
3BBrJ2s8KgeeL04c8Ooz84f6zKPWojHJpcO3BnScGIGQBFT5LUXpZWcXDkKnj6Ezs8UNqqoc/YS3
CFEHdcF2HeoPqBXJ+Uvj+QtAVUjrRQrRAJ6i0pcf418CvkQQZX9VyW0o5RO1Ku/B3+Pmz1rZ++hh
w5myxfnc10Xco4HWSVMBzf4ch0EbBbftuNMk3fLLjs9gNUc/fWIoIhiaM3yOsevJw8SKtHdkwvhA
BpSRp1GNTd5I7Nwg0fubX6sFNwKB0C474rTPyKly46vb0HsoVj5v2VWEaeHcrbUvOoOYfC4nf83J
9UWruLyUhDCKPVitDP9e9SJGofeKyQYEUvuplTs9lTbtrjj5RcloCLJe6p2aiQkVEWxKyDQdNIHo
nhHWd4RcFfUxqN/ki0H/GXDdTwE9vBixh+Q0G94EXuU9QYG00uFF+lxpqrm97CHzAnNf/CzFJvH9
ecTJ9ldLRDkuXNKmT3FyOSD6Wdcs08hZTEyCEjiLZyRo0FoaI/O51oJxVtgGZtKtyq+TPWK+ELb8
D4NMujCjU+VAT+tJVO/Wi0qixXqY7z1U2tOcQzuJQTdZdXjcRspeXZOWU6GSRsQNOsZh2Pf+gpB9
Mh5p1nX4b7gBxdNUOnYArV3ikIckPSin16DP7znXIKOqXLrKK/l3Up1kTusRX/sJmSP3ApNREkEm
WwPpRsNBNAcFNdhKD8L1g1Q18NVmqZyPYrr46YThiYbvU0MkB+wvsI4s+mLUUwCdXLyrNufjeOoo
GOJ2gBGJdBz09E5fPotgnXqT2PQEfAEp1FgAxXVNQtbBS24G7Rsqu2jtQZc3wBrxvw1+z7leOwjZ
0V8KDbPkyNl0nofvEtOXO4Gf2dAut3HuHvSou6qW9Ww6G2a0nt/ZZZ6aeOwP1miR3D2OMn4MJIgQ
052LXrdr/ImnKREAKLlE6JsA+tSQBQIlNTXpim4qR7rktKRaD3KgnNQaMXR+dFbRp7xXyFsWDq5a
QTmsEvJyvLWpjvfSfmYDZkw1CA2nQ+JS9wM059m+78N2A9bojsNyGb5aaRlbOudPTI1kPcX4W34u
eNb+gaP+M9+pRBgNZIBf2egUEPPzLEmh3L6wDpdQ0/+dBtt5p4MvBL1HlgeVGoq4L7jb5QU6d7Sl
K4nADnNY6TZmSWMDbTn1p7q4fwR2K6JH52Wk8QgAOo/TO7kvukbQg7F4veyf8dDX4dVT33xeC0+9
AjSnoJ38QM/0hZB7bUD5SUs6jRE4DlYmUFN9y+GoKAquNbQr1BouOSdsgfFVWbbfvopskKHlhP4z
iiyfA3eqmPvP2Vjmf9Inybfct1cLvojSW/uiMdlaDCzq2O1YIGvfdxbBgjuUvZWz+tqa9en/kKKO
yCFSxwCzTzMiKUf8chleJjMFiz1xl6GWjlF31nxxPHMrlJVP3ofcvIb7SKQtluH6882EvEb+SCdO
9yby8BrapJxiDoScLH8mK3Do9xzqBgsMiDF5BGTPA6yyTRqnJ9ENmN29c5ThqPtnkZn+9fHwv8Ad
1+m+QkVRDsNALXIVN5Twv1K0dW1x9ijr8PfGO0j8vmjr6vSN4uTZFf6lBFIxnu8zMTH38XRuaPl+
bm4ujLfBiDn5fSz2ZGIq+uBMjqRSvoAwf9YY+1mSvauH5+zOncBrz/K3c5msvGruux9V8nYWHA1l
SnKsTtO0txwb0rpHX51xuwcuXBygvK2iV/OEjnlcs2kuVWdo1iccpR7Hb4p1WJu3w52iZi6LjYjD
GsVcmSoboPpyfZbbwqI787hG4DMCpeQD6raEz4ucMORnGagigZS/7AyT81HubcJiKES0xybpro5Q
mCawAv8o/ffK4XYl1aFMvoRhFQiJN9do0Hn0u3/yVzxoxmLmbzClCdp+aMcVCdSEjYeC/dQUbkgB
/ycsVZG+kyrOzXHg2/ey1LNqs8+w434Pp4Xuu+ZYxSRe3Wzmhlk4B9uGmzGRhjFrGuSvb4HmNn2/
DJ/ItKPWMbcTEhn/rFFdte0jUUePUuGXw/gQG0sjvRSvALmD+6QtWzWmucADYX0k/dlG6cJlc2RN
4x1SzyQkU/bLP035wlvImeGhwlirT5r5Xm7CU8m9k7sfAoxRyQVH9arx3liJx3XrKiIOmwNddbqv
03jDkphuem/a1T/JrK6VXnsUf6ij8IasMMOFwhkOjPKGu0sc4e1uKmKmq5/oEy1LqKnHWtlXq1Xf
KGBGSxvnUVCL//YZcDHUuGG3IyFV/YGuGzFFb1/jQyaTNnybzzxDqL5HHurBYR3aKhWPoiGBOj2i
dJ+cWmeKqtjXSg1GobEgGq48BgeRqQ4cy3V1Ll2NbWF82hzDu0oRXashgowPRbe0UKVV9x6XWuRF
2yUrMemyJKznCvD0j2dbF4rMNWE5SeqgOg1vfYZkd6qr4q8+f/M67n4xEssY08gYUkDFKVYlcZnk
cfRA7koexJM+eghiZQgiOBkUXVuXi9N2uPfyaLxoPooZvolWf4jhFzq9kmQr3WZMgrAFoULM5CtQ
17zIajcFDc26uCLAL9rfQ//ZH4PI6+bsRD6QMzdSuHxsY85Qcb6geJc3b94sJL8QkBfBMVNCGgho
wIrKsVL94UpDMsVLJkRtWjfx4siu+dDeKSmU7ERw5d94zUukST8tU6fk8oWMyD8Np2AYC13lfW0k
7a6+iBBG3/Q8XDFlcv3OtbbOIMsixmHBMDKO5D6BNXq8viX5iEH6/rR0SyvaHUGS+F0BokhNzXbt
RLKJRiYjbwbVFY/daUhz3c4mTMDKm28VQDy00VxoSuw9SAAb0n9WFopaC7QO8TLYY8Wh7FUkrawC
6sTWZLY0cxbdzsTmYAHvxSw5O+07llMZkPeVd67lWBiDyVk2pnXxLFppD/ieSn7WeyK+HzUla8FT
fqgxyTNJ2Y4mHzA5ye6VI6EUEqqysVL1J1ErkjUnkeojXC0K+1Uzpy3vWnfehVrYYVdg2pdGEUsY
Y0o18pdrroPW3dCxKgdi09Ru1S4FzvXb2P7mXGTyEBEa1Y54S0ofQPZfHCCyplwYWu/M+zVdubUz
g9Kl7oAaLCCe2Ti2bHtkfrCSViCy4m5BLkoPCPEfXpRvAf0rufo7jsNxJce1E1ZPY7LbzdwT9gm7
bTOD4WykGA0C7qhLIzVmSqU2qUj6PbUYO+pI87y0Ii6hkFYsAFpG46lFzOXP2RhScL8wMWgE4Wsb
UFM29wmvvoYkrDzNaCwtgD8V7hUimdoOqdWH9SAoQ/Xj+oqY+gtEmlbFnICnHFrt+rbUHRU3RXjo
em5Uisk8yD0EM+V005m+9tXef/7m6oSgP+cdTJJNAeJFE2cqD/kjXqzKuaYIyONsxl9z2IXvG1TZ
Lhbxkj7py3gi4DEvrP9wjFZ57uUfEsm+4gyuBgi/KrX+Z7ZIfupylUmvHAPGZoH2EbCW5/nOLVnL
8S+pqcYsMeaD2dqrGcs1FLJVzG6Vihfz/4CjJH3/7d5p9E4ydwTNaXvN1+PZuWpDZbD51IgHgT+r
WyHEqAKUF10ffy5CROgvpFYqn10S+G4Hy78fCdMVbcv2INXtt21Zlo9F1Iix2FMj5ELDNetmOsAU
PFEkfHl6ow8ItlwwQrGK4rHwh3TMdk+yLGIvJT17T4jtITIVm+Re+RFVil1FVaiLsSih8KYa8vg7
hcjGkxorgTFBuHKEjjR1JPj3KugEdo0DY7YEch1EeYe1FtV2MXHBzZ9PX164Xy7f8fg1gouEGf/k
1b0BjSQlGXKfYETV8ZdnNtUoGGh25EfIT8MvCJqoSJCSvNvTFcuPi2UIU8BrCDV5qXYrc0qIOssq
PZvX4tp3hLTPL0sMv8Ucy65bUfIDyJ/JHcmBFhiQbQZtSRTQV2gVA17dEl7dyBVHv1E2TUBjRhwq
rcb98D81BEq0CiK5j1hJZiic2143KUwu4AGyBtVSx9dJ+tde28T5GG9LrdGF/779YiCyqj/iOxqx
BuxF9jkifVEcbn3ziQG7hW0AnaSc9BTXxt9jS5oi+f72tIpPAYztwys3IoPGOpc4mmVBMZOwoP0h
R1Wp88SEMyiUkHvBvgu8X51Gx7jf0DZIFsGkzlMGwrI20eXpsalcz2qOS9ZOtDfIuynHZs4lUld8
hYHKfTQKacMJEqAPfWEic7CUHMtPWsPAV89l8a/cIeRvMpc0VGAUywEnDbE6LbZA7gBu3xL5yXSh
SvR2HMYejFZX+1lXeW/6cnUPZaoQu32lOgnAQgr2DqjgPrqQn0wo0pNNMsd72hIL75A8fH3zy92q
gF5Ag0UasfPkKGUyHeHEtSIDaGNxO0qfVzBjHIUZ940JQfwTG5G48rjgXAFOSVEreIltKGYlWGpk
Zn0Z8VulRf9nlDi/1UF6gCQ0ru/oLNJvSQRVpJXWIGqzlNJjmLqkkZ3rid3jz3Mx8aWy17gesqoK
dc6XlM+SgUa7TSmw0QnYGZ0s7z2LjSiWaYdIY3toVirp1KFPAHT4RWmlHaV+rz4Il2jo1/Q+wCz5
1RX9N2Y1n5RpAiRngZYX74xKOdMoQqJ4h8CgjOcL/IsV5S6LTezD1KadS4b+wBR/meX1Wyraj/gh
BCBzy1m5KRMsC2cyznY/dr/hzzRBYi6Fc77Hr1v1zL78CddH2eRqLEfptMhGhP+bhWYxRPVgjwcH
gP2p6IptHRpolmzsGr9BkC3DHKFL1UGs5DLkVJmpGr2LwxcedN8107ny7ujH4uX/qp2rLoWggfoY
chV2zBd2DFd9D+W5+fV24DX1mTo8s4CJ6I/QFP4+tjqelqxKivarM62kNZ9aI7s4Lu77jvwaydFi
NgiEAlOUhZzRaDIGXgXEeUJhsuwsYcDKWqEt881tlyFEPBZWortKtna/Q5Dpyh1tGsNZF8AyCGtt
hsE68XMufPJQOJ47yq9CHxxr/c8ZD8NC+G2cObd12DsbJ8bHc51jUphRuaa70UR+76l4sRtWtfDk
itUaFqAuvY+vluWAZ9GHL80ZQ+rikn6orDV6PO1r7ZrAc2VFjWGreM9HsTj3lylFW6XlyF4hLjGu
0IvWqOQBwJhlnriXitkGJZwM89z5g8OnFQ+nLHIlmIPWSX1z86HvYjYabLdL/KXDb17Z9tCIzuNC
R7K5/kr+EtMS83QTLTqBRTD9ZLQ1VwHbJ7lwSBoFuMXSVYpcMitUs4TVAQPhgW6mdFDt0ZcqAy0S
+j5P9CeZfKeC269EPNlnWu9HLlIUERfdg4dzUeVk3eFV7qkeDXFFAS9UhldkasBu7qfqf6dH8PJm
qWVt+D7mIvgVYIdEpI5gLefX9eku+gVBrQKLT47IO2FiqQ93MRayJIr7AGqxGiuQjrFMXeMIvla2
GPW/TyiXfo1mirlLMMLwyk2cvXi+30/xIXkMCjBoRlzzEUBx0rPuWgbHKkHLibqeSd7RLqlKSLjC
uHTfq5oMyPp+H7hwJrlW7EpX1fClGRoZUbvT+yiXwefNQiRQwN+nQjcJKQiwFfq8rfHHWJJ6mt4t
/5YCARocLk9UATRagbYcI7ypgPZa2cu8cSRHJXnb0xdkjkEvQv7jrnnulYgllB0I3FOt4A7vs47U
Hy95xT28jpHLXFoky8ak/OUJWZu6NiJErCkTsql4WiswavM0vYvPL9aiqxHc6Y4spfvxWrlnLl/6
lbTDLSf6TjZYcqhM3k22w2UIh4zmsbY5UFQlpn2VpjNro7ohCjgtdKPXmJ6/HyYjcU7inWAP0PMP
obszEUYgkjr+wmISiu+NbNwop1ZpQQAcQrfrpZNM0MpvoFFt/OU8T3WkN1/yD33gDWw8F+0Rx3/j
nDoCbVYKrSSfzYxyq7t6lG6YUGAsy2t5DShCpKpSP4/EwwbQaEJ7d+J7WOngrQMD6gZbDUq5Ol0v
3b749CtgQhTEa+198P5yIPxmEzd5kBI8EHAyHkiwkdgUEvKaLhAOgVNJ7Ee8yevqsaVAMYuXtALP
gy5Bk/w0qVhW0a+pVHfZoHSEMBxI8CjkHZBHiW5YE6HWA5hN4EhRPAk/g8l720+dyXym55qm/wpe
hyL2zqDLzYBgr2BkXTGr+36UUz83Zt9yUPvevd/tXQHMxOt6c/xGOC1vS3HjsSbqdbx8OIl76cnS
IH1clFQhBgA5rzLrUQxIZI4jwmfFaqPOT4gyrXLBzqjt9BHcT89Yx+FU12UYPw7DkmgPpGfhSLuX
LQT5u6asRD+C6dYD/9ZUSa/8CRvyPXRvOs0HAyZIZYKOuxzLh1NVImLUR3g3u+OcCzexRNKvMJmQ
iCVqrjUtHzJz1hsThBwCmHDawZoKS7Pngq9y0DUN7LptnMrCznOLbirFD1nfhZjUXx2mdFKFVmfX
jATY8giZufkc0yoW0kVBBRNaQHImWcFWGHO9UjucL1veDR9sMAdbXEKe8dRGfNFZKA/wBQYcgpvW
jBgxVNig8ETpkekSkv49w9Klvn4YcQGfUor7aLFE2dBynpMQ56JaIaQCgYoP88RGvvTEn3EWGOxa
glTp1+HoX97/6hgzbNcaKIdwnzKegOzbBUKOv0uZdFWQKXO7CxffmawrgTqzEk5NnRLfqRgrCmoI
trZbz37CFCnlTRB7O9pEhaG9KfZOyrSLhGBKtuiMJEX7PK4K5J1tTicmWiR/+M4TycbSLWSUmowD
asb4sYyccMEzWiFSyjeUisvk7kT+wEIPULjTJkvUsf032KzqbZce3EEzEy7fOOyelPAgUMBdX/94
g8iFxPmtXRdNNbiAzF1xF2UTibwvbxDC0NVWE37MJaWgnEDVWhRSoOd2XbGrRwE6GhWMg2HHiYt4
SsWo/mv+MaY6B2hBL1u+er9VSyXVCvu/gQzsYqHHwQL9cmlefxJEcL0iV2l+N5sza6O2yXBPT5S+
s9m5z8mhdevmaxFlQIYrAh3PkhYPrbfUNujV3ayrK5DZra0mgwvh8I1XedscSqt4Ur5/ULDMVm0e
icr1imrhOqVnzoJHzp4daFX0/N/+OtrLQe96TfQ8Y8xzc/Lj3WxuePCQapIS0FnF26r5L9gjB1Ws
HYwK6W3ytiW6o3rD6QXiRpnxhmGcx6e7TWFoGKgPOccnLEW45+0argVJVoeJZMjopdVxHI2lr0zj
tyTnG+uUHyAyMHRl1Cd959QZau4VO92Aers0iZVVf87f9j1kXyEyQqHTDJzJBdUiTyfthepbwOxy
dcet4LbkDHkj6B67lscD0u1LLXEGtol9HmVEco7n7nfeJahO2qEIlPBKcz6vcE1oYwKwhXcy6gUT
P0ToAOWEVVBCGR94CNqIuYaEZXRY/g9JQ6BWlvOCa+sinTg7ogEaxwF3xvnEXpZqJ9s9gAZ/n34c
0VdXfNcMSo9Wrfkqe2p20HYkHtREPBmGFRafdvTbd9OT/XAUUx7IYSA+GLRpJvFtpmVQfW3CEaoQ
YyPIViSuaY8YMyqgaAA0E1SdOOBHRt6xrGrQb5ZUjS00zhe1lsOh8NL7BHk2sEz1Z3b/pLFn+pFW
gNXlffw0DbrSspcjEvNrbCJmAsRe+nkmDJ6YP0+jIp4odGSP/BjKob5TrTYtadKBlABisENtLChY
gxYUF7ViNUGNPV9ctOHolzTI2qx6WeBYXKLlKf1yCxrqRkPLNyXGIcQiRBpWUVam27tJCu9gpyFY
5bq2jw4REzeGWkdN157TiQgVh+T2HQoJ845taN1fQ+jCMNGYMdax4xtfCfbmou1ibhsTBZBJBQD8
7jiFkmZbyhO4RhDLRUjhMdZNR4/IPUrIy3ldSj9wH46Wxraad2Es6JmZSAQ7JVZ+KQP7x9NM+s/+
wkC9MS078/Uk54nTkSrbmsp9f6HJ9+8qZtxGQ9wcTIJnmAMt1DdNmV2B9oWURnlTEjQNhJjFYfZU
z2IFzpyg6eJ8r4FHGJS5jWKzreHvEVKbcP1EQ55DSaqLrAUBfjzcwfTl0K7rpg9M8r+AYCXRWYX4
tREvZ5FATZC98MxuFpqLoZrlmytLoqNe3OQNz9R5k4rm4oLoPOgmNfDc8w5sMYe19P4W4hkeX/0N
5g9HjaNP12pv3+pLrjLhXbA09lcbv5nj98vsMkOkRYPMPmKyQJtD3Aua0bZISTIR89Lv3Ap75A7V
IrsmogMJuMj/aH6fC1mm2R1nsIbzAlqwvJmg2953WCN0JEJEWWMyXKkoX2XioKMKDtgr2naE9aCm
FdnzffqLGG3HSJ/YNDaT/Pbpmvb2iVBcxTifZW9q/9WljuLB+sZj0fIojJLRGMMJnsHjBTozvftR
3rOxXyuneBN4pGpg3seMvvX2tIhIAhlNCmuGsVnTHcfuynWdvzsToRlZHruKZ79wG6CkehE1w4yX
+tF+WvDM9HjQiqVSa9Y2N/MQy6/iG1ANpUfzG3D3+IB75FbelCRtNL+ZHNCyAAmFB2rWixpvIcjd
8eVh4sT8p67+uHRNCmp/p+EL6wq5Gl0aNa6cl9b7c4aLFpyxZ7ZmpUWchI9QbfnjQalciZNvwo7v
wdug9knolbbOH82pjAAYcHdZ2D4UrUDgyabnXi/DNQlZ5X5O3WcXsr4VpxRBtbTOj6gS1CnktrUJ
YDNHWa1qLhqDKkz2XaEbceRhkgoDcJ1Yln5tbRP5FqD1+h0FYWgmHDVt8oOH4Lv6CnpbZTNLkTyB
FY03i78O6Nf+iJmwmd0chVAU2C1IJrFI9z+OdGnzYC6J5V2YXcj7a0MJurpw1CbmbgxvToECefBQ
nlaumgPbJA+qsoYHyzJT/+XDr5u+aYbbt4PfziHzKcfdpGxpGsJF3UVpy3IvAxbL7AzbPop/rTIy
1bbfqicPGDomdxGiDCL6xPCoTMMJkRxSl1hguYr2f2XOWtHRXgPjtdmYyZ6uMn4MKlq5wA80QgMt
QoQAgnRFBo+eYaKDKiaGVEHXdgneqpM7hQeObHFQqC4quVPTlIvUyTAjSIIzQg/ankwtJVD/slnE
uIFb7czmmqi4D1Md58Tts5wnencneKrsbbsNRHf12chCqJq6j5we3qvozkVqmB6jBZDdcAKNnW2B
6oEcPgKD+YkAcnGddzKzWxnAjOdZsiU6Foju8UNdNTUXjj+/MzooxnrAd3UMHKYlfD28tQWLt3DA
UuclhuPOjGIFvsFJmqrOnutE+bz/VXGk4p17H9JI3P4bTaCaW8dUMfXt5z4NiXAksUoFCFgn9yg1
tVIzLF92T6rLZFtG1qMPCTnLlZUB1IcoXvDF2W4JOtl3ymtiIk2ycnwceQmFgVSvFyrS2S2qRuVI
6D6k/7pPLh2bl/DTN5gPxZqIQWkYPKHy0SSF0LDQLKmXZEGZ47gIh848AwmSTqKUms5T/EpxYgUC
zTCKACsJ7/gRqQc3sUXSUYj7j4LYiLZtjkF9Sy0uHKdX1d/pswK3bx4+RDsCT3LbbMauh1lt8jNh
rJ7ETxI7n/wtzfP/q6k0/0SQIvHod0hAY/3rhsA846+9Rl7h3STrmt9yKmvHFWLHeAn5+TNbuvxj
lFaSVNBAYgIGrDPNXnjSGb07QvA4gMIf/KpacZjfjDiryK2kcCRbOOv08OrYPACKSlLmLpRiZUFn
o/tKwu4P+LtV3kWwsUF1dRbwuNPTyqHHQvHJ+nA2MV+ctWsrYiGClrayHw+Zv5hc7RM133IVgxqz
9NyE0AOWE/a1Wkmnu43ddJj07MLXEru2xUm7rvn3QeQBoJ1yaQts61bxqvWfhPyM5JenLUVn8LmH
Tb3wdzFURDPTKCfoDyDWnAZ/HkAImQzSTLGwrh6YkzQ8RTB3+TOTg4i4iJr2Vw5ZX7jW0EjIXzWp
bUdGEeBjub4axXWYFlas9daRryd5SbJJv7eHoSRuZosCzVxUAk+wY6OdaweSztkFFZlaflU/Zsrs
oYEDifwZldHkU6VsyMODvJOGg0f6Y53P+yP86xtT80X4ri2MziTLIg53QRpNn5r8Mr8A/xy1LQQQ
JoUOIJK9jo9q6UcH/148e7XEx1O/uEGyNlh/3596MBr2SSju7DlSr7DMRYYFwpabiClmmnLfm/wj
KTengCnewLN9+zu79kzEjNDKTSJayFuRutvNywar9/f0ARDR/6UeG+2smFnApRs1V10kXRiqVtjr
eWPlCkZD1c/oqSL+hpYw70rcOntcFe7pOmr2undvFLLl5UOhGSml1GxJnMHiY1eJeP9/9iYrmjSR
RRrg8thMiyqhi4CR77Bv2fyIwkiu9bVJV0E3bs+uJjY1xdnuJlAA++zDpyKMQm3AvqR34WqwaEtF
kdzJKUw/WXvPnOmKzVAgqclb7YQmURX9ulhwemil+4M0gnsbvRf5qQbShkXFWI/rg0G3mi6KQKpn
Z6qbMGoWGmg2h/ax+vv8wUxMuGWy4noRptrsfLX1v7SvoyJNqKVlkYlaKqhy7ssssTq4TSyZ3aaj
9l9wHjXZ4GA/c4VSeoWvZkCxw1/zQmpB7fE6VVa7JiZNWlAx3ZbRfHeMh6c3XN+S2wwnjFrpovz0
OL4kz4RSxQQMVRT4S44hCy/1jlYrkURs1UKC11g4GyHoWcf+kILiuJKMwITUN/p8WPkZwin+olvr
lyrexXaDj3yZnnBAsNZjEfp4AYv3KmIYc/gn8VOVG8JSxLb33uu4sEtmbx0Y+g/u6/ODskOzkGPE
pnrx7bcqRvYR1PxbgOfy1EMaoeqjMrWbhAWE35ylgIyPu0PAWCzt4qn2naSGF8fw2hHtV39zl7r4
nwc/7qXby/KS6FyfaXyLR6NbuxdkP19zF1s6OR7og+cggQMYcih7dnt4xuDXi2FrJTBlZ4Ml5sUA
7Ayym0DrhyLu+yYVA0N9xUY+jaFp7mfoIB+M/6nIfcr4oCHiziGSHxFEfuDo9fPEcKbngn1MYRm0
4A9gNvW+5zMS5rTYxe8iKC7cv3iSo/v2r7515r+6oXra7dhcWY8hwbC3JWhU7nUgSpwkFcoI76xY
Yy/r4hz/sb/RwkdMVtMySyDjsmpEpUx1FcYqweuuNiCDxUb2ZnIV4EqMn4AIF0VE7rOkTt5Qv0pb
EPoJQuIPFj/d0T6AvmoTyLPG/CJRPYNCpsDpMBFJh6oMAv3OkZ4Lpe3mnuYLYqooq5rEh7oTeklw
Zmgnaifn/2eJP5PL4caIspbC/JvUUe+CZRPmYhpuGlXeifGdCOOt7NoZN3MIZfxAQPX2kcvHM52H
34CUd1EGfyE1MaACnkOhBhQrdaLvScDW/5086ZCRq4vN5j9Mr8bI1ypwWo5HTIlb1IXf60hUIQn0
LMKZubQhdxPJXKSfbdRYY96/ggl+r8e/bVAIWtJeOPqKNweQhE9KzNqcJaDaG5zqLqfHJ9O4wfHO
25Ykq/f5J186PWbOpoV2VTXT8uHJC1V8uKDrFBtJsb/m91OVM1n8MkjrkHh6QxXfmKftr0GTGiXi
ONkASK8Px2QlzJP4HdUssL+rwOR4oLnED5gcQNFe0+eYCPdlpk0Mni8969vf/E4pp7y6tpP8IeNq
xvcwUl6qCi0SxMCDJcJ3bNbjWfFPt1AjwdNm8HcZcsHU0OVwipw5qvAHUiw5GWI1GXiGeb755O7V
Jmbxf5/SrIr/vbgRngzBFuR0+ty85Ia9Stfxo5FSBvxCI27dEaDiK9KaKq825DznhyzybCmjQMTi
68QkKw24rwXNmbf6jHcHMUjpbdmdlZtusHWy3wb7ynrOgsTbdbv3jDWYJzt8rL9wu0S7cYrMHMKB
ZcIFRi28p3Y6L5QoVah97G+e6keh3y53VSWwvHz714tSbYEK8RGAYbNqN+g/hcXwHh/WJuvCBMZj
ytD9yeGLV1HG+nEAkWjC8i318LWin1AqAiWYWaeXVX6xKKZifyifkZrUjTcRifuDRjPFbtnQGqhJ
yscF0+TwDka3fiY7apIUQufzhBAl96fokVZZZ1y8w99ptFZeYNxScZjR3GT1B6R3juuaz6ZxOHKT
mCZ1zeQ2Yn7TLTp3tXab0MhOMxSBgJUUFCDD/Hlq2vtvukZ01/UwPuNt1MN1tE4kjDkuG6juzQrj
Pq2qCLAAMG9kYbC5FP+rA1dygNNZzW6l+fUkMecDFMrP1+BVobsszXfNzt2t6m19LxwtIkH9jyCA
zRkqjd38Zd2NqmCPfmanmzZpLZ2YTRjcpCa1hBm8QP/KV96XnNQLR9EAqA9FYObbBtHKlEQaBFfR
KJJsuNUt067Kj0G2MylPH5kja+uo4LxqfJWjyFmo1sGC1ohQMaxsWF27yLQA9zNQpNIChER2Nxsz
XctlngLHvSJJyY7dK+TPfGVQtjSiv1tsVvF//+SMKiik7cTAfH9rbExZsKZ4ReE1jaTPPBwjcCbf
E/jg5LwVm92WbLzLZZlbIAmWiX+XThSbAis2MaptdettfYukuIkrC2Xi+jwxtFNDai9agAgtns5T
qDItxZ2PfZfUvsCYzQ7CLUqS0kgESvGVziHvAMlEFRUklK+BkcLJhQpU6t2ppCWLGLvDFQXNVYfw
Y2SGEaPZP32gFHXM97XX9Z6ciBalkCBV7oEWHi3qRbkNkjgiNxMQwq9Tyq08bPpy2KZQCkiKE29u
AFRD5tFx452cyPm1Kf6ktVi/PIlKwwacKO4gPdRpdqpAX/8qEMYqYdSd5NlWZvvp05uirji4lHdf
SlmUubkkJPe8AgGtDwVNgZ7hXY/uxm+gUBR/mAE3qToP7b80gRmiw5ZphUYbjv2DkLfo1CPAAVVs
Zi/9wmGN1RYlTjM0mWCieId9ZLrF/0evUZpqVct2lmmnasoTnJqM+nQkmLk6kU9lGVYSI8nNvnC2
FSv2V/fFL5w7vrSzoATN6ZjZX4aG/PnlRkB1Ls/qZzZ3gUMMbaFn2gGfgH1QdRe9xzjDpXdhR8J/
hrpcbwi/FQlG81g6pT3onXdzsiBjYXP1l6KoWZtRg+iLrYE3SwJLDprTbAk0xrXzEtF7JPut1Xy/
WNghvEbLkBdUeXowx+UCrBqtj9N1LkQp7XGMwqYfKHL820YvAScMT3hXu7Rz1swST3wxG/vqeY7O
SRlbI97vZUOm89kJdqbNbiyLZDUTE5jz2+5ZP4HYCqIGEiKPAW7OtTvwos161ItK4glrQeBwlfvr
ny3YLXns2vuxAxxCcHfKFaBuWUoRUowzt4covg2IswFzgucWaHjNOMDJmMkmnKviYzgU7awfsVDT
azawSViIlsUsZJy2P5ZF6Jiv39wDWxD7Q6nmmuFkg/GNv3adf0T38X4LsnYCGNBP4RQpziABVvRg
s9hG4mtmU+5l9bSgvj4caISg31IE7YSrMD6l1w9JDD7f7Hk3X/1K2UR74mdanin1aAojXh7XDgZs
breEwVEAH43UEwlJ/B4lOqYlsQI5JI+SjyP45IXQzY063TDbLE2OW/eELlG4a1jo+Cbe0MbndOVk
SjRpW6/ThITU0ZgW0BWKtjasIRRNhjfuX8Uev/YWN4slclI+7hJ47f1plsnYQFGR3h0aXolPxs7I
xArK77CtLAQUGJRQp3+be7kmCw8UkzGf6W1bUFL1LsLmT4Qmc2hx6qVviXnHa+kJr2yDrLqBkPOt
39FJq3v9EyUS+q5Xahjsd33wFNK54grmNUiV6x63ROUMcauz7W/1kkZdqnBfowAQI+AcOmnYanS1
mjhf4l+ejreCbZ6WVx9sPiYz7QWIS9t1i1WbsWbffQn1sB/24oYEJLy2scQX4Y3Jq/rQHWtm6EbK
lq6ygyQAtVfiKYP7UbO5d91rDxYZFqnLIGbtuTcaRvXZiJ88sC/ZDR6sg46k+TC4KT0EcZ8pUTgr
ZqYxvcvIIwQDgv/CF93RUvGkJmpD0CG2OkSpPIC8O8cNBW3gXFow08hAx8XGUt4iLTVFI0m40iJv
leMRFG+gcLqfP1R1dcNi2OhhM7e8gR6Dx3Uyay4/V4bz36DQzZyTmPwsHocD1KXXiNdlsJlq+1bv
jIgtOhktCuZMfQLyYUZ0H/G6YvI1cqLPnWTH87ukkYZ2yacfZAelmQBT2VhC5S2P3CEg0jRGyfyz
dFEDAKrbrV04PIJU6DoXoaQr5RzEzu71WS9ONmh42ouGAMUOUCU0xBpu4khdQKBPzrRCtJja+3Ic
21SYa0zMWKdmstw3cpCyEvcX8RtSeZjPVxPdqHji9cHGMP7VGkiMmvxIk6AoFpNPYs40UFPgR0zW
9Cl+R3sGPPWsHjWyLqVMa4EwAfp456n+HfotgW23vWpSmfVlxGz8HTADyz6qhsxQcofxbd103Ch1
J/hoRLIEfGl8bh4037yCYD7uMNtmfj6HAZRlHioXl4K7Fc58KBNebcK7c5Govhp7yzQokcZAo0so
1fLJIlFF9OGies9zCNsQ6pVyHrxtSYYGEj8Y48eHtOVXucbhn/0nrj4pgKck0QIKeB83RXJV5HJS
qLbgqpLwIYCxFbsWiJtai1a8BMIw8IYuUUO5MCBXc5hb1gMMNfSnaEIBEDf00iNu7A+aRGPYIdEE
Ui7sXHB8T/3PyRFkWrAbeTB7NyNBdHyWUCQOQ0XiNJxbiPvUkbbTFN37VNg7YRITGKqOvyfBEMA8
wiFArNT9bq8sO138tLw2mnae2HFMOfwbGm0qvJMxWD47YWcewfQW//+ONhctyQqUWiy3w2zsoo9b
iea7kjKs4dnQip1Ay6paia7RvEhLjKdJTN7iX2F/uNh3v/ApQUgLe/zaCPEPchZaZys2YZvTrS4z
sYkpv4Y3yvniqyeF58vQwd9kyo2QBbd8S8u9kE1RWpvlK2XVjLK4ZNZ2nQjs7eyXFP/vcfiY3vUK
mC6OxTl+hjmifXBK6B/jjR2x69rb/WvJCC85syRORriuU7IQ8nuyADBssnyu2LQDkIlYb0gPk7yI
ikhImE9W8eJ1RbmFWgKm2JnkMS1KBJD06IWV78FmsMcOd6zwkwdhguaesQADvpWKKpaLPSKM5cxj
UYurmhGY1HHkuiKR3bl/vYMLVYGgnA6S/VRJxGHm9gHSdLs5RB3K5luRTURY8MbvmkVXvTrkmjGO
J+dFmox2n/m//ng2JNkbBkkSacew0RMIiV6rEwu0HhDcQ3u9OJRbaSuG9H6UXim0Ix+GLR83GV+p
6yf+1iiXNURXr/Xz6q9yQv9qy2dtuSze0xyGZ1rTY43bdobdCJTMPtW57o9s1yBt2lKmOWNZDlOH
rPfskeQCijn/8wg49osmxg+npC5MhEaAGbuTThbEm+yBQsQ+uoN+wlTahPxFZhPVAGyzDlmsSlo3
C9gGDdtKVeMjFmJiM8LSPdMeKCs7XV8mFSL1tfFQRDz6uJYCbb7JvFIkaKytOZ76wkkiEkFCqYll
8BsAf22fFsqD4zJMQz2Q1PbOJLvgI4/rSoJCogyINz9odrTL2r38BOy1WjIi9u+G/OLLB3T0YXyI
bgUFqy54Qv/2GDHbsh7C6nmCM6P8+hNadivFn7ZXJRuhze/MVWxI42pI8RwlJ8vmJZTJuDAy8BR7
/YS947nR01f4woD+rFweZ5RDI+d0hFscCpFoxMev7STolfvWxgaqad/uq7tIcHEBks538AAYPy/A
7zt+hrC/r8V9qijMZ5L/JeWWnTlsmXZFdVfFnQIFhd65iVirLw7L+pnENSMu3bAmk6wre8Y9Cyns
tqmqmRjX2smxvlYUgGEGvM7dExT61we3L4m9lQjSDiCVprJd3viZtLYgyb5i93D1YRiKx8e4zmYt
UPVch6CF35Jwefw9pimYV27+8vkVHdz9yEUcb2VLfV78qkUIil/ZhRmSjQ+Ql2RzaoxNPYAuR5gO
OIyQ0Cez2rIpVAKZH6O8zZsEHkK6MPST0uEcR9melsL1doJe152vTPmxii3JGFd5kxLUyEqaGqU+
wDp1dt934SLdKX10L1X9fDH1HclqZ3GIP5KOBxFa6op6fmMSBr5RpzUuzA/wHjpEa7oaRKY5efDP
CpYtltSUtyPWL5diQ9/TsFgCpHGFK06rlPjaNiqja3G4Exzrg7BEfyCWrYONq7dF7s4cXi4QFTSA
5n/Q029iY8OO5XHTdkEPE+baUSebpvpz3GkpADqy5rv2J+BluuRkYz4PF4fw7eJyuI3DlxViaig2
+e+eFET9p6tj9j/lbuEO2QjtbVbecAQ7lwW5o60DxRaFAGrABdC/U0kSwwIHlJ8sjRQmw9ux8ieF
zRczA5mMnkNy45qbpiDPAxBqACXTymr8om+LhGkwkK5Eq/gOK11iE6XiPBkxvqk22OPi53yi7TE0
+CkOoATeDW9mlBtfGbajht8XYKM5Vj3nJhhxPtt32oRMWFoPQckj1NnNovhChCBCE1IU0+MoYd0v
kEJPi28+xvdZOYotYfH3cWe4TPiiu3XV5QA5QPkNq2kal2a0P3v4idZqQp5ALMgUnixlwL4wmeHX
GydVzIllN9tMSTvGQDacJ90UspIFEuL1/oBjNmuZs4G8Dx3rAGmZz08UAtLhG2LgDP+5ZPwNAk6U
mxEEKBk+i41JOLAP3CdRr4Wg6FktI6QIlJ+g7FAIVl4SiCSlDKbydaFgaRxBb9cxY1lyP8wX+wWn
Dzv56lU5bvPoSy8SDR8FZXeYNWOORkrwZ+cQ6+MLTufLBnatsL9dycyH0etipJDHIHXQONB8BP4h
hazlm4gGvw8sWKWbnyGUMgFXwecw0er4zXB0y8WVOSB/ZRdiWRu1odWskijbvVID5D/swe+NnJ4L
zy+EsPsiiSIsyTZ4uYSx3OYyVnAqusc3wX2KEo4o1wfCsDjJPLanvxbNxCYG6qYB7IHNG2OBgel/
mKpWMQUlVzS3inGVzP9K+g4tfMRWsyk8A01IX30dNjJx2ESG00jh76VPT6yK6cdZs89vGGa/D6ed
0qdeRhhq983qWRbIlq5K7853gfiGtCX4hLo9qVIgWFUComIbalSJCxNusSmO2PcCkAm9cfMGOWTa
cpVaNFOSsyLUSr8FstOd/JnjF4Z6y/pcjdoQW33F8E7zA8kw7nsbkQT3nA4Op/I0JWpISEoO4k2Z
yDlvPoIt2jNiJ8ZWaaBFLRksCsbSPJ4P9K69c/WKAZuKhB4ZMjMBA3zMyyqVh3gTo12ZBS9awbmt
sngOHe6o+Kmoul7r2thi03nNEl0QoWKV7iwGUHE2/1CshqD5BrbaJxHXTEZGH5oNafh1cAixKu2/
kDbvPnVPJ3NkhFmsWcwUOLSJias4nfsw71NJuceP7c91DXfTbrsieUzAj4LR4S39dqUg43DQEka6
vqvbDkA0HH4AFO8LpwDTRebugEHTpLdLNeL7k6YhUmLErV3IFMK74gKKDwabOxsI/2wPZuB9cVo4
sxCb/qGlyaN4/kQdFVoRPO15GskZ2wdo2iDgHczXfWQH7BqDEROvXItSYMdPFPIME1vpO9PwJWzU
2+reDBCNobWhrZx2YqDm1n5uPiUmAyxfsFYSo+OsY32yvV5aweJ1AmG+Nq/MDgm99vBVBm+VVjId
5GHdszaIDBvQjHiUSeLBMPH05tLivc+91JTYxunFdS7g4AmEuJaFnEg2yPfWstiPU04vukBatWxY
gBteiLZy/jqaWmE18os9FKmyIXHHpM+SJVH63/kGaS5EfGnOx9iCqeIPJAw5FpZv7hDRM1CHISI+
uvcDbQtxL8s7or8+ufBb/qftk1OY05hG7PmeSDQXVq7/oIOgcYNwdRbnhP6olfJvCqw46FbkkFgV
nOVTmZ/K4fQdZjrh+b7TabTW6VfFMxe1Hk4xb/9XBNMshPD8irMeMOi74rx94Lu9WmxIOD3Q/mHi
pi+g6jAzEW6jft2fWcYqtlccN4kIvLfL827AF18V3e/RIsKYxuJJNHrQFLo9ulqn03aMPaorSiUs
VAxjR24k4j2sdwTc1UkOAJbeC748dKdI/38zqEKf5wFKTGP6WQOWBRYGt0VqEZcKs3ZLhjyaG+8N
owOr5NcL9O1dRLXSmfFMReX4J1ZFHIu4rckWOpqE06eZvOohK73AEuNV7QAelg/8CJkys7cQxfvT
OoYN4CRGDbsajLHus7bsQ49+CVzOj7Tp5BhVUc98pvTQDscUijiddrohwl7KyelTKWePQo9Eqt4K
zplNeWPaG+hLYQdA/rTnYih2ODcNd0bKOSEBGhXyFHb1byv75H3yXz5toJAfvxEaxvYG8FPnsVX2
ljMCjrlFmsnBc/kgTGeXB/oTkRoceQpL7G90h9A6QomN+fiT5frjPjpW5KVUydFs5UGl1nR2PI3x
Ff6CuFiXj1WjpzbL09ndkLF20OLEqDY9gfQqb/7lO2y07wbX3TiW/aPPzM0TiQmtA9ktILP7W+u1
Bjvkwbf9SKEisWPD8tDvrqcGcCicwfJOEcf/yLymuGpX+3ErO1rJNjjg9WP+UmxB0VyvOmRX5cxd
HGQoZImLUXfw7FSqkAy1RWmbs3j3kP60Wm8AP09gUvQSJOo/rVii00xUeBpAviuLffczSpMHRcY+
yCWrQyCjr8BiQYmrBbN028kONJPhu7GMTPOhStrRNUrFcsCw8dWS2wMjyeeVFrbmM/VZjlgdkeri
GRZw2FIPZmTjOU+8w1XFeC1/nXzhhUZp5dBTSZoYtA6JVx8NQ6mi5A46/lyVCNgw98zK0hrCGPKb
crohQ/hTxxSgzKU1Mlnb23PpFWwDm5uvKdIGM+969NcnBLPLS+i/6QpTRXvskc7mlBBbTxx2id2K
ka/lXkCMsQPa6XQ0uM/gBNKwRVpBayoFFIL58FBrC5lAqgdsfNzXvEFAwWxpiCBE6uB2PXd1QcFm
AylCMMpEl4NK/96siUu2lCFXUGdrXMPD2QWa4M9iBVzIMNdnoUCKRjky0qO1pBSC/KkJGnGbZoXe
sbz150Hj4u63mZ764RYPf3Klo8NL8GmlJ3pf+5SJ1G50Qp0pR2+AWquUfRyDlNtjtNoqKU4riWjM
9isVM0M1iYhSidkL2Cx+5qzcxLFOhk8jtk5I5POS9/sI/70Joi+W3iPGH9o/HOINCm6OxyiuiouE
VVMd3dzOz7tf1tW9UxLa3zp8qLh3hRAIlhqFydbceWUJZDpRPwbvBHwDH1401/y7btcH/K/1c85Z
jLn8tfgbkjCzYdQi80YbN+drXRJlo167D5Tf3JxfkHHMy/hclke6yP9BRk6n7944ISo35SJfDySk
OZZYn7/hV51ZqVfGX6/+lU3KFE5Qrx8ZSgB6pzNJAoG9s0SBvknMtM9FX7R8OZEZHc1dpEOHfQa1
MRtu1EKsEpap+aYwK6PCOoA6Yy3JVNAnBeqSOgFacgGo/HufxTBG0hS6r+G6jy6kHUTWl/3voz2U
+f3cOjuXRniYz8kM+LQKp4+LE6ML8DH6mBxKh6TOVwQS3dFgcO8JkwlEHw+G+TGq19yHL0fS0kOB
oitq1bUoIGxl1cY9IV66ZWlPqOL393DozLH5q49Xo+yNFxydUZALbrDSbc6xGAjgQRND/OeOpJzb
ExcIrzbVk1Fh64gJHFV1DEZCBOwKfmkMU/IbE3Fs4hmaQ4C5a8psLs7/uE3rv53LQEG7NhILp3ko
G49uQooPRcpxOLZxW5KUGn0LEZNfgy+xvaeLM+mPJcp4CwUaZuBtbsWPKaKNGPKO5pEhlv6SO3TK
COqwseKRm6k364w4zRns2R1o0abz0JvY5QxgbzBmdoiVyDEPSmzwf6dhrO+Qf62IlwWFn4LNX7JZ
B3spKAKmkzxVnpVQmlmNIpmcb/gtNqJcHrwsOD15dtZxiyFiuT3H70rigzzygKFyQ5vkdDndp7nj
EcdZPZBlnUhEEiZKPfILIrgaK5Pti/5bQ9JilJsmv0+Z1P61m5V93H5/n/MWRYrV1QN+PLSMcEfo
9mGCnzrUGfxofP3kpCffu4/St3bEfeykLz9c7Xd0Fl5RmYwReEs7gGgNrwxNrP3o4+zlWAn5KhDJ
OLlBGa4ESqseaQ6clnAwFI6uudONoi3ODQ9gYABUAcZegRzihbcf8VTkOowIoO46y9BJlX0L+W8O
ovEb98YiW/Bf2W4gP/oPcClBslyAb5Y6BCrTu4OJorg6xNIdEm1YbG1GLG8tzJ2RoePVOnWBoZ0P
neYGH3sf0Rfjt34XUvWYevRv7JEGFdRparstWd1r/b7ac4IW3olvsNETzZHExeTLQKqToSMVNXYS
Ixvy4hUfy+pjOOMdA9tJmALB4HEDuIKP+UB32hXenXZfDusrdoOGaq9D0K8Qwzkft76zuK4dmdqg
PXeNej3br87KSvHRvq9ZeMymTsVHO0AOo+TSZK364gbs6oml4r7FoHhtLjZgyKqoHrlC3cgLpFfb
SbjLty7Hg3BetnQUbj7ubxuRky/PxSD1hkCf5XPPpYk0BysBNChOuOciYiedSdYJDTTaG+BSD/e3
0n+CLdDOQRXcvWRlV105FrwxxmJgqj8HkCyvJiE4cJbBXcI40ZZh5s6SVmgeVisql2CIrNV4LEx3
qZu90Knh8zRjbyW7DiOmdql5YeWGs8RVmrVoP6wdisJAjAtTXzNkXwxuF4NYGzagnnVTdvEUGQMp
MziESvCB5NRdC+CgVtpYAz1J3bx3/tv3pFygjEKYSnncPgmXgXwW4kBj51vuv7CkNMcoZ14FXdmd
Pisj43L8nXQCZ8O9LAH9iXrVz7+7OaFwIxwECRuJCap+fdz9adyuOWxeBb34gzuXBEnhqAeL65tu
jCfvCoDwkhk9E7GJyjVE9GDHZIMOty3GfPOXhr94j1JS9sXLwBaGN27SDwCqyBJCzVV3Ddr6yXWd
EVijfRzzSuL488dmPMCe1jnGofJBwCP/21xxrT8xcb1k04apTx/Ks4xeHlUQXtUo4BDYmpR5v1hX
sLHtApRyNtaw/6H1H8MjgWbM5G4gFwQ9Podrl0K8JF/wEnP4DMSF5QIk0h470XWmcFo3JIqXfKIa
6qUmp+JHLujaW4+HAFuvajVh+ArA0wgtDD6L9TO/9pXVLvvLxFug9zFEBboUvaq0ANvA/9GAeybw
th1+pp1VVYYL+WHKvNX7sp6x/pTG0yxjVJV8dux7+6FH37AKdw/kRP6c9gH1PIH7DWnRR18ID4Y5
vXIBCfJHCpPc6qcR7GRnKlBFghqX4q3At2DLmvlbNFQDD28EUqL3QJPrgiwj2HP5gq0GT3zxySwE
oZLte78Z0mNVFSscg3cVQtooeiEdyXEb5pbsoJUmxv29oZlM22fyYt4isEmfdBPzoE3sL/YfM6PQ
fekuB/9XPeNGQkBbk9UIWMD4B35mnTqCD5rUhPYSnRcHi6dl+NHy0iEVswGtwHRDCPGXIOMtFmRe
tfRZMsaPZqzGYxyVEXoJ6Mm0quB3ZaxtnU7hjYUlY7SiD7vXHYTUkRc0CcPVU3THPsjn9ov03oF1
1OT1fOqrT+GDdugS6pZpkeHrN70svBODKhWYuv37N//0ih4sG3JTRmRIuT+RxJmqJPAFnRx59sXy
qAwIjHDKDAtXF01Q2iCj3sSjyr77CuGcKhkMkwvSXhJeMkGM8vL5cLPygNSnEsvwCWRtWCwo4bnE
gx6k5JmbZvo52TzEqnP/C9qzTJLCxsHwah/i1FEICyqDLJ0L+LBNu4KyELuZwUkCeuPrw/4+uqdy
1mLaoTLkdWTmAUme+52aFbgaf2zjVufhQp4ajrfg2qlkLcqicXYanhem8kRyoY0OcXCLwJnkRnTO
3STw7CUyxRnQXoyzqaSylFy8w429gAVGF71pRmrtm02a5XJnOBWbTol9fvxASsJtXN6aHf8laH46
e50Lsa3Ifk/Ej692EVL74KMTzdNKtvOUcqeFM25INkMFqHpVLOqzJUkarCk7kBfApQoS65u0NkQ3
QJcRU12Qurq5+S0ZuMyQxBPWm4VWLiX49wO0baSHSStNX8B4NEKpUB5J2NnG+uZJapEvy31Mq4YW
85gJYSFGkOQXsXco1NtMgcsoJ+HxpfvD/Ly0t3H0xVhgaObxQ8N/SEWRqkVCapMpvhOCXZB3z+0n
6ouFr8th0mxEBF3BtMoJ2oaagYrNDyZAGXx1sk15vsqURu6ifL8G9ZZoUgUcNn/U+GRTsLkyug+j
cbFrEwWRYvMtAz77nS9iYb835/fngOxeYajdhVguvKCR5+fIEp+MIcxwH2xapC5+Wkm053Q28MEr
y1D9Nyc6GdmfE4F5Ell9a9Uln9hw/aeidvhT1KpqlnJWYiJzqNOEUFUxnl9U5jLB6lILTsjZdZ6/
tLed5H8wqS3e9IdbZbUCAIbFlN3CSRKLm7cC9+Nu5CTZZ2lio8p9Dd6uWf0xXnWSParoIqNxTwPh
qYch6qD206kAaQz4n/BhQFCpwZSfZWd0EboVr8degGteAfMY1Ah81votVINWurdczY6UHQe9antx
ziQjtsVyEUh7lw9CotmGP8nOqydmHzztIhBBQPh1eS5RbRVvN9yZqFZU0AsO4ATEnh4ZgYsWQjZk
aQhu9IyzZu3GoxP2jBR6b0Pe7G4sW9/KmBqvG23m8nSyCXtzz1s4GG0UYDAU5E17r79FY5oZVEMM
vK5Cg5KMykvrThXnHdcO7EUCdfH0EBSRM1WvTSjcvHE3nHV68HTqFqUCNy/DQW78ViQwwWbbBi6I
aRlQH8Fo4tw2jStmkmRlst9D5QtwND0+GMWAG0T5T93ktQaom8aTlvz91qH9wYrXyHz1XK3k9Hwu
AFjEfqIvCqwzr8NKJpKY5lZiOno9zcXWB2TdLrGkp/gvO5TgIX9lhx86759IeTEu8X+Y5vqpYjU+
c/LRXHt3ePK9cCQahSQ7SlOyddTsdEMfmV3IlFExfa+9VIFI4JITrEGABPpTSzg95pfJ0QsbXQFv
cin/DF25+9iGaa0rD95hnzNAotMZMrUw24XeMup1NtBPJ1nSt/V/711X61s5CRtR0S36ZapCshZq
GOpKEJPUqE38s+HPb1ckPL8Z8t9tay9e/WbnIj4HxaE9x3vtxEMXdFMUTOcqqDr4Ah4oH/Z4LLwW
Y4xqZQnspYaUgliA/vbOn7oAPot+ZpKNmCCPTwi5uJBtpfSv7GWD8GHczvOVPJW4vXruwULneFq0
R8DchKHrW7x3lDal3QQBayNS40AyfpgHYezWYLS5gkusPoRJw5yKgeP+Str2s4FeYmURPEH6YVS+
L+Vv0mjZe3/NrqF6bT4vqKfk/2MiOajkZHnk8ywkBe9gur6miQBOXeI78UwIXVq6AyyhioAurXlW
dtoYFNx9GGUiJIxsJYCX9NEXihHKmq/G6z9pc8YWcyyXXnRKmOqPi7/vlnLmDMnBLnF6X7FTzApp
APRsa0xdzsnF0Yiq26u4iJXQw3lrJ0qIK1LcWSh0XM0lcFN0UWiFhTtaeReGWSWoW6umr2Ptk6f3
KVz002OKtNq7gghwRnESz3xd2omzWU78SQAANcVAZGyooUzeoV16RkrnhNq76OIlgMWvNHGofcdr
Ns+KQddrFysCGij5xoFMCCNj9MeFR1ytU3OmlmyJBHcp38jGP3ZycJqPnzfaa07Qxdj8qxiWTceD
5QDXdW0OXfBwQq5l4qv1jzZ9ERcHCCIHBo8oQ0BfdZIhYsh0aCO0aoPSh13Ar5PZFlwXQMUQR2XE
eYfBeTPEbgUGVfocvHf+BxSkEcB1kLITf3zQ0nx55APdZ6La7fDZPHqj3+/wHvKUJOYKD8Ha3fiW
/ip8c+9uEr7veM7rOKFtOUAT3l1Jjh+68WFe+QEnq7/NGAuQgtBrCEyWTNZT2BIs2mPHf3smarjO
fslHCIPqOu8Cgril13nEkvwtZcr5z8ps89njZnkwDP62pdwTdHlRPH0OW0xwomnaUqiCx7nxPNnF
WG+i+ryr28Oj11Y4HrayJwQQqrUEbIQvB+jJpc0+tPJi2QBCEZCTrWh9mr03pvK/xzw5Jp9Q3XTJ
RMXKEuG7haaLn8nNL/vHxzK2iYerV7r0jnZw2eAguXnYL0KC7f2S/eXI855eApkz/yS0Foq8xS2Z
ZSiMVF37MXroqrQ0eMvkpoTwAGlE4pD0mWk0SvBS/lpW+GYKVGe0DFTXMn6GRpdN1tc8RRLiEi5q
sUsZM1CPCRy8AVGIJ+PXSQKbBnUiTyIrhNfoqA03i6JzFTzlbzexHmhcqBXLLhK8ijnlX8b8B2DH
Vzkz6n441NbdQ6z20ReajvysUwfBH4+uiWHgRqVutvHMAbRtIBXhIPdP8zzhUAVTUoVT0fHqobbF
yTaC4pxn1U6lJjzpXdgoN6CFxpFOVi3D2+aRxt+q6whIQ1FRS43Z2E6HfU1GEutOsYU/spXA/yHI
rxQ3H64y1/Gy37wHa0muUcB2FtxmwBxat+qz+v1WdvApXYQ6i0c/GQKXgVITmNA1LBonWl1kIH3n
3fJZfgwAsgfdYXJXKhbxi7L5rUD+O52IW5uAsU7g5abHheruYBlCQe6CkuAPal5kLnzXSYz0dLOH
pBxdTu5gam39awiRSMlvr0P/RWbNEy/HTkcvXeBdpQRWlWjs+7IkX3NOlv+Z6co6MsWvmDrg/PV4
tCKhHJ+r1NNbE1X6HuW68eYTh8GOW+YNgazszGO/os5vvFXdKg/7UoBn+m+FZvn71uoKZUABDExz
3hNwlgR/pIfRB21QGWbuJFFpzmrv41Es+WV1gKlxm9SsnnVjE96EuToUy78NVpz6OMny3sQisIlH
edoXa+f/ICaOr1kGeu10hRcgk/gvT5ohGGBq4lzo9Ft2IwoJmIB32YdrjLxPX/md0jL9Iu76/FP7
uy+NK1QdAcroaC/d7qoOho7pD0QUeTyo/6EeJ1VqLn2oCdFWTet+SR9TWquQvTEBQiPaaz0ThJpl
Z8e8rhYhUq9COV436mEAyBpF0yNwb2W4gEawkyFuxiwjeOtp2dvqD2pmLtsPHymy2k2S/rLgvDyv
yPcWhUe1thIEArXrLZhEtMPJEwHIYSZWsfSxOTcZEv6jCMHUsjP8OstjXLNQ+uk0Ht2/542xglMf
fcCP+zNh1RsGWfHCdsHaACX0G93IMB4/hmwN8DvRK+VvjB9jlc7961jOAuOzhfiI7JEFJu3pxa00
zVO6FBKdsri+xPn6+fV2CKd48Q/W9m+5SIqPnRFTO+27vvoADSl8p1jxc0b+snIlVV12tEG1VrfL
ih+DYm4yRqTWaawHXPCcfGaVNb9PXSau833Lg43g09s6zlZP4fRiFPNtQ0FBiD1dLEw7VS1/sTYg
rVzuyQhubqjipl9kMw7eppw1ZlK2d0NmbZkd5zso4FigMuySgWPmxvLQdoxMedbDFjcdjyeN2cHC
SHZa4wOFwaFIpM6Vjf5sunOon5wvLT8Rbhlo7+ndg3st3IMilpVf+tX6uPVcqWtVenG4eoAyPnLq
lVNFzGFHHjsoZejmP9Z1BbEV9EqnDKyGldj9JtXh2BAcdfuhYQrh0AtfqqOQUgdrxALj/zQF81wo
kGE9NGkif0holiESDT6UHN095/be6KKH+BG7lPT1yhzmkaLUyWBIB2lLr7tC9MjrHAwtDNUEBFYX
rg10T1+27+HjUbKZ7v9+PP76UNGCQiV8fHfddBRmsaI7vyKDzVDZaV9CfT195DEFNdT0INCqg4L9
V0vdcbI8kbWUzgiK9qUKFYXT/5u1GGdF6J1DYlFsu+su870XE1pJfF9+S2FuBTX1cUjEwm2cWzXI
ozjZBDwqby16W/KzDIavqYuqNbNllzL2cACIAqZLnnX590U0N7YGQdxqUrok3Qrz3Usl9vOHKye9
hPVI6phWhULjoYspKJyQy/4E+kyM6K1v1+/Fw50D4FOboY0CZINQW+JUXa/jUaHoDb6fbn4UyyU3
uCILawGSafxu+DpdNW91/Za+WXwh8Kj1R634kBxK31CKsdayZepg9jZsg4mUza3adedOJvC5uOl4
ekfTlrHzRFHxlvgHuds9jvZC9t7SL6Kpg/R+4c385JPW4btgcZrB1/m6DriegyRb9Z0IdNbXpw0h
B8Sk/5hqiBr+oNZoZhX5iuy009bSjJnrSNtofEY/FU6pcN5oXHPhX4tn0jaH2QO5usV5q7BBEw71
Fs83syCK52bvc5u6HPYzDKU5pPb+KGOO4CXNQvsKGQhLIb3olDsXUxxPiJzN1lvONJKkmYHN2rQ1
aHRHhXUHgEW4ZPFKj0w73T5F1H9wcAcu+9nVTUc1Hh09vKADfk2oyA8m2W6AvZxSuDiSztXz3klS
i91KuYNiSie6AtMGQhcyI9HsQDL6J7aqeHJcgq2BzBah3pXltK7FyMsj6hHJy+PyvdqF1iBBDXge
xsngleh7Ekb8faAFqr7BNKscNY+uc4dk7ZW1mjoGkbSFP9rZX/1o9NFZ8RswWIpr7JN4LOFcks5j
OZECxrr/N775o9B0mLuy7WnwSlJBDkIqHz9C26XzF//3PMcR+NfL5JoJaQku3nOHe0Llt/Pv/CSr
PtOct6QCaUoFPpX1iW9NY99k+hsz202GcQF8+gjVHjUIUp+m333ruPMxohZf8XG4YTjC6xQ0Y9gr
AVFv6nQW3VZoCiZZYN6yKlu+xV2KzmKenT81Ed7l0ufvD+iXJnSeH3Cf1Elb38vnpH01Nr7aokSw
jelb7b7KDbzXV+DMXks0jRxpTugvJlJukn8BKfCgqufIMkkVAggITWUwEb+dZhGugkt1+SKLxIlp
S4cl+LQw5qPSaTmndpU+wT7LXsoySai288BDuSkybumOmpbkhnis5kVKRR1FDJnZwpD7eirbJSDZ
GAaXw1n5V6Fpyn+wP34an87BXg14npc11yDGojtiitswyDJMFKhfj/LkCHbtMZh/KlCLjHyn2irO
b/tS/yNcFSXIAN8viCc2X711IR5rQd4ZjxShD6fXL1G2QePXqIICNiGS+nXtmvy7qy5XBzcz59lY
FoHldC8XmdVRr+/6D35f9V7wx8njeJ2HTYrZxJmK4bF9MilkyQW4WY5tFpH9dsd7s2vaM5UdKL+b
EKtwATWvlTvnNvBFPrI36FV8AZVaDSF1vC+gmFis3Zb/H3x2UtgyK2cYk5cH+08q8wrStoMAUESc
jYOc8qFcgF09rGCsFCK1D1PejQG4NPNZwWSMA3QRv4/WLjHMuWOOPeespOZLguj8jTwjxP454/V9
19iY/TOzEei/KtwgAj/Yv4Me2nNnFqRpW2Z2U/8cfdyQqHMm5Vh7+wUdE0LoFz6cnqQQfeLLcbdf
UWcI3MISLHbeDsH1lGvHLw75CzzY6nm6qqViJ8wmDX58fGnGwjDPJDNj0z9BHuWWES+rQ80lYWUn
wo8bwwY4V6Mh9vsibfwfH/SmbfSW6qKgaLBOIvXsS4KdC2lNhN6Uy6QiQJn8LMSHz5SP0mRGp8zz
oBcFJAEvttzjQPR1XSsZ8YVWBxpRMIBfn6Taotdcl98Hiub9Wm6wSn8LVneXQYqqDO6c22/FEl5k
RaOTXrwDeNB1G9EBepPsGQmdArbEtyLGoxxIKcjb5akhYbHSEsI22B2nDTWGjXs1UXuBjo0K83BS
unuRKlQksR34Qasm3QbRrjPeYVmRHdxZGTwGTik6FFS4aGSk49YAl1vC9XeJy8gWS5ilEbRSNbmn
xQsng3M62xtMe3BR2h0kHkNhNVqF5Ui0go1tIyCLl4Xsne5n2uopUPYwDMXsr/pfr1sspCQkZF4r
NgShEVG3wKFij0sJelSiNqv1mDhduoPD2feG7CiFJXObW58IWWsuVKgB93QXilMlyHFZXaAlILo8
2NQnOPaE7MU3LNYzo7u8TG60OO7vq9lRwvIVOb+O+erIrPHR5yCI2yLermzos7kba94S+hijzUNX
Q/FRYNuYRrTHRBF3b1z7s/cYlZ+KZZCdLWz6lKrLt69XSLBU0/ADXv5yB1I8zNQBngE6zMP5kpdH
z6eWWdvYwE5Vv2JDMHD1z4A3MPvOPXazJDTwI6F59j1VJCISoNBkDBaXEghOkBfDmSA7KSfu6ieS
UpXVs73NaUavHZ0CF0/kaqoC+FqsCZDAq2QQqn2IdA1KtmhhKPqelUTO8i/bf4GBBEXx+OIe3ymQ
ZpcyOaeQYMx3Rj7c6KVB+RdohKi0Njg8TcMPd9v8mxKd3jbH8f4hYyS20gyP7pDbMNhRzqhc+LfO
PTvZf2XZTxXLps9MmFpJMJ+j+GH3z4zyezOkjzulFo1/9vvPtEA+e9bM8vfc8UrJzJWCumxypHNJ
YHxEjIWjxst/+B+6I5sLb/fGxSYH6KiVyYg336TDbKaoRHVYLXOTrJgaCuWXhOdOykVddhb3Hwfz
74i86slxSwVSsSKWia+kVwklharm+xY2m28LWHtjwn/b7bEUu8qLHlyMSpvkNdYWZwSsAekb5lBB
mpSOV3LjXvXFwIIpY5WEivBy8c5BrwhPfuEcXN2jr9OCtRO13zeGbRSVZjzAQUBAnlVVCmuC6HT9
STjQAj7qPjzwkkeUzdtaPD0wadoqUvD8cHGCmz1f7rKQe1+1u+3S9N1BlwPJKVerYuE33QpYkltb
V4+aQrh9FS0Va3IyJB9ZvLch8EQRWIbZJ+d1XPmFL5wJiMIeXMPjwQNH7NdxNlZHwsYk1s6q6SoU
f1yPr5dv/GIeUYalto90ECO/YXU8oFmxe/w+g7MEeUs1GsP+3i8HVCjWCsplCuuPLOL4Fpdh6nGC
2rJGN/rE9vi27MAwTSTMOAwpVfSW5CZ4XByzbMOCBR60vdJoJzv6kkr0rkiJjWuB0Z2+mzwSOnG0
NLq1VetpRrzTmpI/ZzbNA+5N36g94qve8Uk417kuXUaktyEcfAqyf5a6GwcWRnoXPslGAOvS678W
WNA1uXd5erPmb6QiiaLI9xXzRwwjhOO1DG2kEZa92ngQY+jxrvKqklrb85IOXnWjQYnsHqh2v7qz
3QbvG4qoVmj8zh77qSg7x4RYump24ZuwgeFo+5NVwdBsRbfRBdR5StH+eGizhhp2MkL4dtSjF0RX
f+YkUMaUXLAYllL63R+t3m1PJTc6sNbobBAuvHSsnmkd9S2ITuP6TUIKpUo3K3085JPE2hNQcVnU
aPnI+a1u0igLCf4iN4funQN2168s80jiAIvUDxGQpoPeYsNaXqBlN+2e3DxtBMInNfZ+Ooh4IBjn
DmN8b5jCMmqfE52MByVZKNARrsF4Smutl88u/lswetcpSKfZMXyUXoBwpHGseK3/mnDX5GnvSii9
a/vAya9z6zfx2hWVfXPlsKev7yTsBa1cyrmwrah6tMnFbd+Sq3eb0rF/ROfaHVk+aEV82N+KVfui
mKmZJGXUbTS8JnRvsgVcBhIhlSAswNxQqKazjLEGgK8DIKUQMssoh6rCwZBHFwFbrSAskycVAGw8
1WQmYZFQysmAOvAVV2cNy4Sbqxz/UfGxex/0foB+YpPADNnPyJZET6wI9kmL5kqZxdtcQTswtggM
Ywcisk+F6E7PSRnmTF5qqsyL4C5TvCNz4QdvILxvl6u5W6A0McoAOI0HcmAync/eYmZaSEPaJr0t
FA6N9zEDwh2n/KBt4wLrzzCcpoJowCe59c3+ATChTcZpWkwJEnMxJUiuYfGsZvvHJ2OOrDz78EVP
hZwf5ZRDY7tKMlOMrU95mtgoAnoUcn2+AC53xkm6sCK5ZBk+KvUfdsmGJG6DfLV2GL0/p2QS4tCB
BO2v0KDnpYrfbc+YYkfwXdVaf0YoUsTaOzWI+M+dEceI9e9r75k7dqDxVpkI2GTdT1CrePSV6uzU
Xp/j/wnSi/4cIkOUfyAcdIZSkhF3pHsRarafsbpuDV78Wxss4fwFt4TBscGEQC1tWhPtMqNAfMB9
3XYXPgBHSNUHngsrPJ87HoPyP/WLuYDdoGOEzqc3DQA6cviZ6xROsw+CWj2vieLGCkL1icPephyS
vI5K5/u9aKOz3ut6OlIdlhoERTwlKI70iKalVYbdyv1eHHt61VS1GIRektGQOZdCyldHht6Oqo7h
mXgEhB2jnJdjtVTqdfb56AqeGtzVzF9QzjvEJL3118Ug/bmthLmGvCCYgGU+FHCSMTUwMkI+H1aT
T8J+jgdOBBRhFQK8p1Xw47g7VF9qd3PlfMjwgwTk2d8PHnXOOOtyIJd3A3jU3t4//XD/gTQAZ8bq
R0AQR+1638/yTyVEEjRdtLhIC4bOCs6TGOZUAM4VmDuu4Gd3vi+DE3dWJkSfeD4+v4D3o9xEGA9j
gQDn7JqDN8r4T1Iq0urCHA0za18gF0F7WnDHIepkQhkxNllwD+wjdPFTQK+CEXTWEUArxOOag8Bn
en/3bVFYiyUTXPivSatCzZkkNrhMf5B1WhfBACoYCpcqWHLXmK8H1dv/3tpFSYpI+LbVmqDj8b4b
HQC7MvOV1jYoqmQNpXSAG3vpYVD2qIA5PAhUHJZN1VEf0ty68vXgQrtM+VlFXtvniCfYY/XQkBmm
47QfmLxAdMITRbFpiSmLYAhrlfWB7//5IEiF69dmKoOH1xD3tSv7CAfduHo4tbm4Z7UmqJkBVqKF
mRfh7Ciz53opWOdpStlQtLD1oL3HMitKgBfmUEMX3fcOJvfceMEHENM+P11fjz5TeU4fcHAKqqp4
i2/sdAqWbyyXeLyCyFtnA9dizF+2RtxGERpXKB7kgIljng3XDt3Eg3SKPGQR7er4L96vw9suTq9b
2ijDo4QT+U/0p8jp5OPDg2ahb0axfhyHSQzftfh1hPIegIKKqJL+TijNcEkGBLKqjcOq8J8BnFN4
KgnfNhxyq/YGeTNKQHnPgqHWj4X21FBCqkdvzZX1gUMAPhXuYLqdI4wL91QojDs3pQHXSDsV4b/1
qhs56Pif7Ko6DKiF2tr2hRwzlhGKojrdUv0t5aKhhr2SunlQdahT2uNYOvTGyICfnq8LCqCkOYb1
G2xihdVPCk+DMS3TyBiyWthTYssa1f26bGS/aNTSDmFCvAxTAATRkW7fvkLN1reWX3b+Gw02E+f1
89Jk392IN/4KKYlsLAC+a1E7VV6pnrLsJyd+YPsp4Ph0e198r6TwF3oSAjb7OX5VKtKrDEhXScGl
OxrbaCb1vZa4UwCSy5miuFDUEzpDEBIYbtV4zHONccZjqVCyuPvaeoFkX3Bv/rbc2USfKEWBNy9/
+xWwSPkmxIM4kIog5KyYboSqhr1J920CfUvAGbNjmp5mmZwyC96AYLdEcJodwTAqfMA3aKNTIvKj
LwY93Weh3twozH0jlx3m2WQNs7zCp8uS0KJ04ZB2xVX2VK6ZNaD6c8Md9a6oKY49IS45cIhKEvNU
jUjjI/mB0pRgKZnXm132R1Jk/0hJfnAp3GqFQYEH0Njf7AUHqtIaV6XmB61ggjaxe43beNd0gp7e
Iv3Xi+xK3ANOrigHimdWFqaoXFkBnEIIg1siTCjpf5ueWmuWHZlbwDS2o4/zyhsekhutr1hOwvep
6Si1hys7+6bZawbeUO/CEMq3xFTBcO06EHcHCw4Y3JrX61jJyo9l0sVPWalnpgx3sI0M9P9G7Eb7
XwhrZ+UGPnbwAxbnIXTRS7J3A8UekKCck5TaEVfupvajF4oEYMPl/CNeeMN7VNgO2P+BzdnfWbUc
fELTQX9JeK7ZFpISU8F91FIxX02Psl8O3PGbVfsHZueb9WBKuRhw5dzob/ILW/OYCAWAdg4gPU3h
xv6l79wNcEus4tBOOsF7reviDHS7BXzVat1XNagQwGib6I1Pce5wZ+s0Q0xzBy0HSwE5753CmgGA
aP2oaZ16dcg86Blj6W8neobRmpxwcdv1R5sbP6EccDIqpTfnf0Dk9yPwieuQX1X706UU5WeIde0e
0n82yzLoJ62CT780KY9cVCkAMmHyfQW54xUM9H9KRRvdOSn3LDH3zYjcu0gDIVLxOodPVaEpcxV3
oGt0NJJRpoHLloKs0iUNVXIbAb6IMiWOVXs56QskC4jZPSeTSPJEcNXiiuYcHfIF2kH7BIl+YV1x
6PrIYcObul/o8N2G/4DVxQc1p7QcyzZ9zxDnXB5ls9tTAjmC1L63gXV99yt6PHal3U7+0MOku67G
NjhD3/NDr+yXghx+PDea3ldezBWJuh5j0uOqDjAX+SqIX8hmhgXc4EVYXGtGRq6jdqE3wtjxmIX9
chyH34nKneBsjYqDYXvh9+xtpV3HInPMGnHdCMcvBwNTZCzPuR959bJdpXII0F0GnnLvsQtkyJgJ
wkozzq/JjCxzCLmKN4ou9iQvCn83hSOEWOwroxrl7pCFhGZsf/3GauW38KRcR+KROvZJYXWpBJW3
Kmg3JsnDYCd3hSy/jb8ktmqnsNRnPQOlAPr3kp3geW5lc2y2LzjJgAfM0uMelsmhrLO1w+FGd0cK
8SGDV3X/2tuIESeJKveidh6Io6svYt90Bgpo3j3i6zz64JHy4IwpetjPvuSbaRmqN7qyR/FgBZ5k
/zat8T9JQ72vx5MKN/en8jliNZ7tt30ohLxW8tcvNS6GhfN66z/yBctlhGIrmRJWEK11mHFWT67k
aOkVgw0hLUqa0GFBfq1+G/QbsygW3Cn3iGsL7c35zliexFbK8wkNBOzRFUmpN7GfkMe0s4gdXz4p
NbjT2SbDwW5tSNys5kbjegBK3x17OORKMlHr+KMEvBwRQ3C4WGxZTdh8xWRz4fJm6ogujYxPXj6+
fStnfvKOEZyC1xEZMKvo7uLcsZ/vCtpFjj8jGMJZ38SY9JSV1fkSla7BEl3wxHDp+c5K/6XR/jvJ
YV40/Fw/3nX/U7OQ+Wlwjawk5fDltEbC72t/dhFC9Xd9BW5hzBpeyRPlH9CXAemLd58oJVecVUNZ
QI6m2PAFsE2URPObk0wm+3TuDozKaDgbryDcCcf6r9NeMuXQQvm4qrWBTIW+ASUGKG7ph9JJb4/p
hJ11QaX6slfekq4kcbVS34ZGjkOw0Izn7vQwjpxBLSi73uWpiqutIwQ5F8LnEqFmKWxrf2iDbxxv
z3I+TmtCVuDutqBtqFDH1M3dLilZXFL9w47T0W3qQH9xsBxNCkCHxw2OZ6TlPNIh9kNJaxnbsazc
U10Gf1K/ibMNk8TWLaIMBg/zreytlOTf+KqZzcl2lH7skE1o9IHpgQO3ofrJ3I0d3X5SDFatsdWt
6HKgGdSv8IIwjlZaf073RH/BHt659EnKx+y5m/CJcYyWkUK3UN3VgAgmCfx4/nbcwQOglb9zB/Vv
wyWi2r+j4aP6dTtkZYZ2gJpJu3uF4i/HAiZ5AtPxbB5IUBpqpxjAIF9ovyl+lmQqXRSY143tyPzv
iHz5/RdtYywo5JtqB9ZU90pOPoHeU1i0XPqaxWfPXvRnm7kzyP3lng91AaPjMz6tL1JavzpnXj/s
WGD0wlLsFX+uR+sH8kaNLpCEgcVyf+BiCAKfL6lAnKQYTzv54kF5b6r7Z0182syYazAOHrYN3a50
QhTzEVUQGHkLKAFv/XjBpZqAq6fSqmr3dWvOe+KtHRWGRSPCqzLgwlYKWrFSKcF0+y+1m5kaSsnQ
yON+xTOKZ5EkTLo+ZEvmVR9SR223+yVwG+d3VocVp68inxrB3RxdgtD3tr75Ayl6T7ktVrUR/HkB
kCqRk7vBeiekG3ITgQVbmeIUdoO8d6tsDLfyiyRqULnsMwyxHD8qJcJAIduQastvtDRlaW5lThK5
QzvHiKulFjz2uX/nLVuy38z6kiZGcW9iI6NA9fqKsSxLTTkmvC8vyW5tlVwq5q5Cnyjg/MRqEdrf
kUH++HlI+xq2oXtSq1evzajfHj01Igdn/G0CUQlqChKTyEqq8Vp68tXoQf73kJa4TYCPzgFO/wfL
xwdvLQqIWuj2yr2ss6WSKRcx9VPi626manJKm864G4Do0yC4lPuXR3vMls8YVfjzg/s17r7IccWw
hen7GH0EU6FFsEhUzD7By9wqnoXX3wg00mJ1ihwzR4IH03eJ4u1oHd1tOUSQjfRbJUmn6tMs1C5f
MUKVNpgOTadunV9tiSK5HCVI32WgYIqsHAUKh9xE3MxxZANPjDwZqfY4hyAPJCzJqKgSMdkNntYz
A6m2nULThRaPG+7eNQUYbeTY/zoFScysi2DF6nV5cPXwwBPxrNFZR2f66WJhg9PFvbRl4Km2FuGD
rL1V+QupfVaFDN6FjfSj1uKG7qpZp0PBPVC14NMaKY84F4ffeMn1AOA9ZYK9NVOUDekRIE/tohyE
QzoPC5Cf3Ec1nIlOJzJbFf3S8qQr6lPz00GvUUmMldIfBC/ZRBSJDaSK+GXmwH2ZZna83qIqgxrt
hUegpqwDb+pyIvFxa7+scHGnnmXtUWJ7l0dHRdSYwYrKM+clowAwhnnohHNuoZEeXYmhzqcxZGQ1
Np6I8yZeehrUTlrY8QU9azTgePT+z2Vu5JEd5Wf/OYbKxIkV1w0wef8CjA65PW+/o3NKv7ymvX/7
WnNMwe2rsJFrTnohz//m4hgk/lEoqP9N2pqFzRX9GEPx7kFRXZEYVtP2koy+MARMRsJjc+4EHUYe
9wHGBQNe3P2vnN8sgOCnV+r1qtBAwlE90pSusXgSf2AE9nzehWYIcMWYpoK6fY6Cg9ixFDpw1LSz
3LV4vkzwFZ/MhaD1kZ0cvAf7kfifzVKwtHR6m1EPU1CUEMsAQh+Oz7wkusJwjWZr87xRisS9updV
Mu/OgdqXqFM+p3FGqoIXxkoGTaaHAtE4fNWSDEGYO5LjS0dSyRtUNyOcGNDcRC1CdnGmTW4z7TZ/
Bld4JX9ZDs3d5t/iYgSvN9JzpqSz8aqiUZ5KiBh1wcIo62tVm6gDG4Oc++2E12yoBmWzw8lWZMFU
bMANcpmgTN1NXRHe492oQWcxLDyEbl+JtjJ+AuLZ2UeiLKco4HTCaCzN9XiHUnrXgH92wG4cxb9X
0tbma8bITAg4VlU2dpnYwRuWepExN21I5JQ2W49kNNRcOlKap1DFiSo1MZb0P4fhbanm1SYiulQ+
gcSyMWZnXGsrIQIj2gT+4pAl8mMtFAjXOkco1STnLzkFf8+YQUY1U1PyzyntDifxO58404Jsa2gi
8N3pCg7QC6IOWZID71QzHluIpU7eMMRmYQ2Ya1sV++dqe2AycN1aOPCOOJr4CDwdIUZswdaMhQ55
rFXo5u2W0QZteQPHuUW2jIfSR4SVJOFtQnF1BLTyjpiwnH5n+9+gwgfke+xn2BIMdr99+ahnmbvw
AGqzegkvVL1cgFFSIPqtFMj2Lscchvsqg5HauIsKwZ9cA2CBuwWLn4BebGk/6QNK8W0EzSLteWjf
RjT5IH4a35iBfd8b7eIBAL4pKs4A1pTlmaIhWwOVYWCgacECBfaVxRGI4i56OTlt1TR56xcneXKX
4hPB3gBEyeY8EAy5dYha2Gruq/jlk0bNTzpf3FJg8hf834FLtsvOChBCHSRiZ4Jcj64J8IW/6+iA
Fv6WuGlIj2FC9QkLDbMxgp+3ETUCeTBSCwF0m0rvM7kB2NK3TwH9m5huWlMYBsGmR6xbMu7XzDeo
mFGc/4i1yrq5OQh2pqVB22Lh764+z3QNIdG/DczKRhDcPZHmFRDnE8NqWQswp7QEFFPrSCx9BYZZ
kYsWDFWw+Qsn8HuVm/9UK+PCprCcM6v4h3uc4aSbCycShM3h8UjteeErpbTsdXBo4r5DycJdR+Ky
tw2QoJVzeqO7SxpMERI7qmRX0evTrya9dIz0FHSFia+cCOWlxHq+84B+DzOauELVr7vufYmjzDSn
kJRrVyn/ncFliGInLWuFlH/lkNi9ms3fRayws7WUa3l0EHiNztrBbd/+HCBujhGBy5EgYwmaG9x1
WOWq+BrpnH2/QieBIXs8UlAXiPz2sznxPU5clZ6FPCYlSP8kEkHgHeHX2pllJoN57z/JQMdUa7gD
D+tErfLsIjpsdfDSIhLfizPqlIPCesyKgv59IyJ0tSYH4NPgnze30cfZ6OKREp4QpZlWA3NDddAr
mCk66FRZ6hQUkHNzv0aHviiLlUddgfSkpANw0xJc6ImO7owY+YMUe1/S6cWHCj+VLkPu4qo6zeqn
yVLz44EW8HjZpDfJscluakgrya1SSqU0SUxkabuCvutIV6sAjYeXSnyFJivG0/4+WlPjWIAHPVsJ
tPA0+oSMkgYYqb4CYT2vC02zoBvD1pQKG6MoDd/BVLGCYP+LIM7QTmo4CKdyN/A+ITuZZYwIetRA
s+OAjObJK8IqFb1YGFto1JwgDJV2gMbSwC8Z6nkrrKK5Dn+qDxJFCwuLt3FgjD1hpMpQZK7AxZxu
lnBWEorbyZfACiW4tnSrB4GvBRTDLDXkWZjW769T3TUkjagLtR4ZFtxpAC0rfu3s4gmq+i4o7vSL
ooTS0VKBK7aj9SxOefyjniCPYBdQGZoBH37VL31jZox68g9Hqabv7RE/Kskz0lbeP0/G3h+UcSvq
DboAd7Sw9a6ex/PUopmGqVrQw5FM1y3nO1bKXkzSHr3NiXjMJCn46x7VXeDJarht8Vv/x5GD2Xb9
LUxeHOwKrw5z0Xphz3CJ2IroQKJCkQc/wH/DidktADpY4v1Cj59pvxyInZlgED5jbqH3YopZkBVi
aA5iPgBPn1id1oJTIvDmWnCuxJ19YFwas31BVN1elVldErFN1DiM2370p1IRQmY4Ix/VYiVjjhOo
ys+RoinIpQ2se4AHzIKJkv5L6JklTUMWfStpOqX+HlyRx+3E6fQIYtzHu2IW8DA/EWCXL6+C505t
Zfg3TK+Y7UYGzz3Z0nWV3GZy9bRWT0Jns6Y4JGCqj8CGx5bXtDJw7heVNxZdNZ+Df5feUduPCTWa
fFHWBTl3IdGQbIjDrX9edTwJdm4sIdZkf5dJSKpEAMfam31yhl1uqXkyfthI79rzWH9OYUszSDzB
GVr36y5oZQI0dn3y4xFY7B+g/LlSG90ZwlPM7MduYyC9J6EbAlpfAfGGdhD+D97fgSw0RlUP0Nwj
DoWF6MAqNS5zYYPN4UZ6AGglEaLL8KqUh38LDvxliMunEvCixjFezmLz5vThzePknwjELOQxO6dt
bEyIBB7uy3ochw47y/5Y4r5EMgg78tXSfYYsIA1tCvfaK1O1/5u76fHzcWOSjBfIQeQU8IzoV02R
YNvi34qbkVvIRWcdrdWA//GEwJTY20kYq/IqSsdYPxylQZ4mZ9iyq62eRsIBKiNjll/PF8pXmELO
WgbbfTNUb/fekka5wwVYAmfZxLkL0c+do4S6TJczFwcvJhl1y5C3dHUH5+cb1TAYWn3wR40vphOm
uBBcRD4P3TXvRbEL2ML3NXsitV/LS2GyAx7GyWHuqiS+F19Hj0BY2/8dVm76hY/Ks85A4jRJIo3M
heGdnajDli+mCirnLpxYicnuGU5UryT7zLbuAHV7LUbMfGvSdR/+91D5lS3ZM0Nm4P3IsMF3KYrh
VFZ4XmMZk++SoAf26SvfSiOeexg8MCkHYfZgKGMtPvjHypLF6Hh9Mevx7oC+GZzmPVRqzpc9el/p
bnNaxl2u5K1QPcp0qVtnugpjAtf+8I+yFboaUDipAa6nvxLuNmLlyWIoonmqz/QLwf7X6NS66Qdl
kXLHtFqDz6iDTfeJgf2JoCFdDtYBW4RvX0T+9o6FcNqCFtXDd4dw68NxFshhTP0KI0ias1kVjAEu
+Lhzn1A79qjGV8gElQwAVdh5dJz95KcSwl3cwA/Mop+/F6Gm9nOIXfldcl9JJnXvBBdRrHy2CWkV
rXI6t+Q7G7ryW9DW6X0rsDhVoexSQ70kXhh6CVPfZn3oJqtbwx1hCk8G4SiHdeWJciPVIEhrjf2R
wqhLe+7ISrmtoWSOltaLmLBDkEgBdVsLsQ7j6LwHdOiielaTbKltqhKPPgVvxpXHvnlwEeBD3WDJ
OdxTNAljD5qaFkkM6sH8LMq6ffVYCjg2+BtQesemM8c47jdm3e8C9U/bwlS9c0ek6gSUEz9RVgzu
kq+xEfBvt5Fe0Fav1S+bCHEU+GTKisv/62v/R00MjccCzDc39mdpWmN2o2dfyscZJ8KoOJ3nYgIv
70/gInQxcgpm8OQ8FbV/TtQDdWN0LbaeyhdemiISkkzlAj6DaK/nPBKYKzyCIupKVEOLfvSMONZe
vMTzt4fHTcX8ojgfngAsJ5YFoi9Ssrxwns/qSG4nEJm+6EtwGl5ehCA8nrNYSqo6LZgjUPwCwZGu
oOzbS7e+VVS5D3J5vZbxkpvMcXhAZMzuFpYqwovNEqyjY27LOdjccBfjqkHEbH9G/9YIjDGShNKY
+ZbnUwua2cJBQkO0CmYxiJaP+dqmXxVYDqq+XRaTLgv5VPglv1PQgZK7i3czVyeh7/1V6SuS/Vlw
x70lfARzK8MGERPimQpA9u/IzTEMtauyI0EgpRDoLRPJWHtx1V9spxqiY/kLr0C/vyCwFObbW5HZ
OPQaYWiyJmoHT1ztPnSF4+mrBNbyOy1t7Y8s8XgmVK85es7DZPNOx13nURQu+SepyeI/qTKFBvIs
LqvAWNXNME/ZROUM5rrp/1JnKne1BUa0lERiMXgDyeAdbGh+6GmwOWkAg8gRr2BNTihDsZR6y3Yr
QRJSmHrl//1x6OU7EUw5f434KaPdOMaA87OE7ESbo4x1HVNMhUDnLC2+RGLsytIc7NZHpuFLz9dN
C+AriR02n04Hl3yqod0yAsuKgh1/OdUglJiJwSxollesk/HfpinqX6P/5fHxW/wXiSBNCHXrJobH
4DflTc6qQReR1Jl63370WhoEJx8U696JRrk7YScf8ViIssz/cv4Tpw6yxG1DvE7hEtQ1w3ZudnHb
djrzThQzC/yFVR0DnU4RGSqR0reYWeG6RFXFhoS5CcFMZ6enoOcYjmve1qqtE+hWyaWktvT8gdLM
pC8i6bqorPYKUmLgsWMMwS0yk9KIa/zxe+k6kfer/fIEHfXsXA7ls5v+OkUkQRYTLYgsoyZG/dEj
2MX96r+cDwrJAzxIpI14nRWvrgVsFoQlPrLZHLvrqr4JWMKslKzsXOthFof2YNlnrR0QOUBcLBSe
JGu3TqkHCctOlexhRSFMNG/Cf0yZ8EdW3eCR8qQH8BldGRkcNdNraTLfABhh2k2vWAOgy5eQQ8fd
FyT2WGfr/bZ5OdEvGQahatEV60v++8D6mcNEfbXONJw4N/5lm7yh8YsUphZKJ+wgsWDKkSQLsjGV
KjXM+gljfgqtCbLpWKWbOQDJ0I8IRfNydmoC7HBM5yXdivSvp68xszlt7EPJ6NcvrE/5Lrg9GMQt
Tgoqefci49th7Tb3CDCiQGJdLABZQjQkSbe0YHi5PRWVWNBzz5v9UHzG5+njayZ9ayMB8mWpf/fY
imPCkkd3Y6wq8IUcFzaZzDaR+pWqsM5WVRYQVIICHXc7ArKxde5CX1AS9Lpa8kA6mJNXUQGl4rb5
QxBM0sTTpvRNfz1H8XKS5mpZgdvqAppIk2sHRpkc65Ng0IGgR2ro5J/sKuhiLUCnGg52oaS91WCi
Sr7vFvYELt3Yd8y5Hdx7YAanVg+v3dreX2+/xAvX3gR9L6B2DiBSKxQtxO0On6iTtKxajXbHYQkt
wdzYq3c+hTqxW8D4J3hTX4IckB27ImXnrbiEEmxrdPSsHpNt4qoicRSW/aRA1GCKx/GyQyIyUTS/
FLr+nOEROf/UdDJVIsojtG9ZJB+2sEln8LOqKGa96sMDdvUS+MJdj+sxgWmvj2W4N7Lu47p/6p6S
qsTf5v80a/3EDJIqBoXZdhdEMOxjoB6gs8d2+rJUnnMchSKxwhB50ih4OcCTjRWd51fmu0W+UeY1
2FbVxT0YPCzCqDVgURHu8/pJ7QjvXwZgWrBGrKTaCKm1RUyBh5judOOhIOhEOIpvGMkjR0UTJuGG
Q7xG573bEHExjNKRfCk0dUEV8zkp87UsUtrGTqVJnwATT0FwlviYggYyH6lrswZhQWp6zN3SouBZ
NuZEaDOXThAPPhj8vsXq2BS6cyH1utgQ62IsJV5mjP8mqQ9zWoIxx0ROr8K6oNXMnjEL8fLz74Po
DpWkBHKLmnTR1Tr0Vg22pV6ZJNV+Gvf6gjtmgMRHV/E12FBZ4i2cuotTYbsxlZql4D6Mho+dFjGR
+DeE78iG9V2bVjktHfYO/35bVUPlkMfahFDHL9zfN9EhsjnJh01u0oAZRLgvYOniUqsyywdx2MjT
igq1SdFpzmhWqqpeLa5oQHijMg5p80nzO6KzZtzjMgFu89+vIUhPJtu/l4nN076ji/RYbKp+nXsJ
SAIZOVE0Msq4gmMUacJs/qbMoutvticwBdjPEOLGaCRa5lN5Ftk0BvdpNec7LzisN/MLrk0vJ+hV
BHoOV6c2IZ5dPmMMjWz+UX/eXp8EtyHQbPRV5k7cXVBvy8LATsdaw68Ws8WyX+IaiZRij0wIBv0Z
6XjB6sOxUUgEZSK1wQ235Ybq7XFnDMzd74dZ+ibACc2RWs4LReFo5S1LmdDGg3i2RDMHxklpGOhS
iQqpzY5OjguXQMlXFQA44AWMGq0G93uZrzDH6zz5tbS1cF7gaDXy38JJRkNrMHQuZHR+bM1c442x
MmAlowJyB7Xg52dwf3aaYvGzDMjHY33cAi1fSS9P9XOkBQ3r8FI58fr9UizMqhVVm70KRgMqMlI8
l0fKb9pYBIy5jhGBlca7R/gxw/rTg5JAbAa9M63pViJThIwSML8Ou/gyeQXOQgIa6w/IGfBIwsyP
aJp351Z0ju7m8Yi+t4Rt/FcpdJcNs+4PV8sLj32oUxbPXKjMbwj2sXZQUzpgGohOYYvwZBzUabtL
0QaWJk0nGXhGXDDfhPii1mH+elX43Ssc6GfQj8Ugtq/Obw45EsvWiSgtr7wVIL8SlwhP1aMD+upu
VuOWpEQ5tA4tqTrLf2VErqriIdqMjvgsclinnpBtxPgbsPEEK7CEbPfBznpn8qbmCWql94nRmX7F
8ZmsAE0TqJXRTpyTWMCohs//9Rob2oM8YHf8Jy/osXIq3mmF8IEQcvIZr+dyIFXQDU2MxY77VPWW
cERjytRxx9c0ozMApHiuI7IFCxUKd/oRfdRLK2rZ3Ob6W8gOMb/psnpp0jHu+HhaOy7iTTxGgI/y
S8/+L7IO//P7SnWNazjIcFR7aCwh0YDISoWkTCSweHIO21QYjaLYNT8zSTW4ylTeHKUVm5OMqg0i
zmxMjixwn4USAw+SvAs2kY1YKd0YeRsndlbuAAS36gaAcbAA1YpAOzq5vPslj18p75LsqgyAOAQC
igpELHXDYKOV8xWrZqa1jHCrWeN7y6+09b/Z+/oPjJ4BQadtY+NBlDZ4PlxkvcqdWxhOgH8dumo1
rpFQXmqSU1CBexO3oI1lTzT+eajdwY5IEN3A7pN0m0wgNOsuw5QDq7F+nDNhgOEldJam4N0jTPMZ
G7/I9M6HqdxoiOUYOtChkfvo3NkFJn/bpe56i79OVR7PsxEM97f4s/k/FO1DDwiQfUhO4mGXk4eA
1BLJdAkkC3pvtREmXUN1kujcXPSvOSRpsfqnETfWgZaqOSNZxakTlUbCCvQ2HP8KyMxG4KPEJWjI
X63mX2lJ2BvHiPazkMiZTNwGgpAEM+OTB9fIeprczRmhPt3Gyt4DJB8pwB82CthNhuClqcdaJknT
uGHhKpeDl7ZGK8Y6CbZYUyvYkkefPEpaWLGZKarUrBU3NkcbpRC56CFxtoQ2sOFvdB966aUflXYN
x3FmaZT6uZe2ZnxJMzNZ8bbPZHbxE15fj5tBVvVrWeppNcJNKyP4HaWGa6mvnaZZljhneW7IL7Ir
5U9M4SxA33Px+HxFJGC6nM+CRmt4wpmh4npZsOC7mAtlIgPgQW8dmRsj9Mzro5sRMBnH2JaJop4u
7PWEFLW3g/vnFQFv4kDes9QQqAS0oON1uVVZcO8EuEws3wzVq6OGkITgttrBZIuJ+DaNqDNqqMB2
BGNkac27TA7xJM2y0+ZipU8KLN9SPpnNIhpVjR5H7rgBoUjCeL6BW5BIu3xw2aPGGhBJBBvK/aFN
QFRMr3uP6/fLwP4gyhFDpweAhg/FuNVFmkFSUdbfEK0NEOGrqgw6e/fLQ1RmptngD23tNsa/XTNX
9X06Mn4mD2qLZQuDXGPuZfjVKIi+XAYNRhu/EnApyom3RMXoW0gm0UD6ts71Lp0JYpwtvkS+GHMo
1xIVn5YLLpBeSoIXfYC+1G34Sx0wocl2bmWUKWOYgEfUMVb1eO1B832QEblMGkyQ3+EV1IXoUMIX
CS5rStnvpk4cEYUQimyi2ii0zruglihRsnXlmKIZ5i8Y9dld5yWG4ExGQ2Hlv/lIfwTMhhuD3sA4
gxOsxQb/DDC4CkOK+8aDU9koLj+Bkhu+NbOb/RdNAkAwN3CNct7RDX1FFdgvNl6A6lkeqQ3qvx6J
b4zocfU+/PCxjsM1hcvMsTDbUUd5xA1hUiYHgp/AbohyfWvNdb/vjfBG40fxU4xdnZSNcLaEgWAQ
rBkd5VNNJuHGD3ERvfie3zCrVZ7DzD01E1SVs/qMEvg5b/OL8jv+T7gwaZ9E0T+4rEbbeIekufCX
o7ovs28uqVUXejC8ZMy+tolAm2pj9fnj4Q+GkynWqi1HK83eFrHyINPRipwFRXRA38KUOgLmLnDd
THkouhDCjv6CjRL4YvwF8u5NnxIoTBPTG0AUXsxDKJ+ipIiVNqPWLC74+UEevlX5OnMBf/LBaGvt
lbaGioC0fYKFZ0kTDGQ+jTcIkAzh6QXF0x0vkmhJvpe40Ek74FFLiV4wX2tn6PPNYvapLUNNWC3a
rPWs0NyA4L801V/KVrnsjmaijRV4YAigPDAXa8LAAs9JAo/VXwVWbaRsAJGLrXdzUWHY0Wk20n+Q
SeZs3429CVp3mbrfsyFbwX8TBmM5uerWQbtco76A1AWVmK08U9EZNHRn6KzUvHf/Viq+KfEFullB
sVNCD7EiApXu2dxxXAPltpF9/RBSvnr7ke1frrcdmH84qp74Nt+RvwBgTwKhPwR5yGy1hoDHDXX9
Un+o+GELkmYTU/0A/6CvH6zXGpQdTCBe7gW11hcN6ehmB++aOsoTMS2dNYp5l2npBfl7WQ12oYLy
vgZRYzSdCKaj2tOwbStHMvf6SIraRvL+F3bS2BPBDno+M4mNf8SjFbMRPtlxStUKyMcZTJKCZAnO
ifK7GQCpfNGR8WPDgzeC0O2jx9TOMd/Dt65TNxiigEPm4zX3adU9dw/7+HpOmPZkX8cGTlOjblng
s0SGdciy+1GpZO756CqCY+3nMiRPKTnIABlFFIrarngEpTAX57MG/C+zsL6bjlsA1SkbftIMHZTY
rFGU3h+4VuHCmgnYkaDctmR89k4yj2cSqm2uLx/VH8DtsuxQE+uz4WMNDLmHrvL606SscothM6Qf
CGPNcWPNA/bPEhM+o94RSMRC28MsPc6P66+pWnGh3d6coF2McLUjycxNn2F1AtxGyjcU3xJ43LBS
L+4W/tkfkCSBzc+IDHSy01XdMBPi9UWwwKFTReB1MbPPhtAtW54UqiAjQXABUh5VUsv8mzmrAla9
vdUDKBbcxEAQ+SvhpUL/mHqNLH7L3doS16FnZ6h6IjejjV8FOaQSC6yO8V+fVHPJe1ybhSBALQjb
9AJs2yo+k4s5VTMwZM4L+L1lGCtmf418vO1OuOidZxmN7SVC5J7tFubsncfh+2iuDX/4/mD0kcKa
guZjxM6DV+dN8Liazyhs08nmA5yoaxPobcBH+Hq6KdxoiB1UhZAOhDStEbTRG3HH1Y7D1JY/6VU6
1WAsgk7HxTTX2iom+3+ml+YklHeVuq/mSFW0V9axhOlq8pgDrvFWJ/7dACGe1rjJ6zLhEgktrGKC
XBegr5pjxqFMTYoHMWUATTzxnJ6puBNi2M00MoHdSlxfnYMFpZD6+K25CAzZrsBFB98fUyA060AX
GgE9ASUa9Sj1AqdfD90hCy4Egqb763zPru8kYcAwIS+FTfhbpt0NSGpeYo+6TlALEmrisfezUkpQ
Uphvg7/pCKBs5hL0Bx60wBPdqaFafZeKMVXF9NLr/xrFJfJb+IMbvOvgV1LTLgm3cdfByxo4ZUzJ
CHq31QJyIJLvyanFDLBP866v/SM/aqchamThrAirWP+lGaVXFhNborotq4xzLXZIH6PadUY5pQ59
NQpUiAzkBGLHQIaR6wRcrMIg2378Au1MH7k7RU89kJS+JwuAKYqSnmpJRatymUrMGDfx4HkkmSB+
1bYUYbUqKry08h5QMKNt/Qr08qlDjmjOzoEIXBhQlqVN7PD4Daie1ysIjN+xaSGFw1Uwl5xkdSPG
qcdQo8k5VVtWjXmgqm2IzcuD3E/LBM/qvgh6qpykumIRn/atmqD54KToKv0prJC+zzrgzRAaipI/
TJ7DJfipZpy8P+ACiMjFa8W3RfACchxcG2pby6nBS8rJ7ZBUN8tgAHGQ2BVo/jbJzVcRHwF6qG2n
q1Qz9ro17CEPFsTbBA6iEfE5aTplrMQJjRcj7N88iDWr3aqxwi3QbpxPHV8JnEfkHM1b5qpsn9gN
h5MPSUl5g+qkt41759jYMANDsugZ2vjWIqKvjnZjviotwjCus1j9Dmf9+kh6OVGWaztyDclISiFJ
mCCScSL2qmVt3bQ+PEPWLEpjFE4tPc/k9BMpK6I//YvHJ6Xa0IZqCnCKbfRE3suhoKkM7HlVp4OM
bgqlouqb456a09nrLgRbpfX6aiqt23ln9rzTanecYmV2EIsZ+VtRlJvCPTV3+ZmDNzNnh/joBvFZ
UmqS+R96LMo7XXP609bJiFRJ0eff9oeaT+oYfRCvkr+Dg3wRv39i+UdNjKZhWW18wdtlsLfLJWYp
bNwHWlAFldEH6AGEXH0UAodn11E67PJzfb6wBz7Dl+fzfgKIhDnzVZLblv2YzZoiHMIM1QYtjxEC
vJ+eORZ3rdF8NGjk/VH9CWJxtLrZX1sXvm3OW4Ep6fmI2IrDJzfGTMFKHXU/cIhfOOidDKb60wqM
y6apsjtNBb+54JElO8umRa0lvrGWE38SBH1OtQUHxW60TNuC7fv0AJCpjt6MioCXE3W6xkAfwbxe
Xv7BUSU42xpN0MAyAPN6/K5G//1S3IPuln6rhEx/AuBbbeuytb8wRNqMEVo/Fmx2KlxfXjL5Gh/H
hyqJ5F6I713MBHuTKT5LfeOBOUah9UXRwAcOImPEiV1SA1ZFE2mXtzyq8fjBF95E9pPlXVTpthif
46yRvdxlyilAV/9gCJK6IVc0RrS+eYthfQWxyFk7ig+Ux4dzxMVG/OdKlunelArK4oodiEWk+n7b
3r57B2B/bixPxTunOFcppXfzTjEss5UBe5HO3dmTIFpf9U4Ny7qxJ+3Wg6DL7JtBd8OKMGpCzESl
YVzfXIrqbRJuVQK2KdqP/J5xOvt6Q8cRGrWAzErDxJlgztWlZaEo5F//unHDlZgsY+4PeDsO/ISF
MASMKv+gXErIUQKE99TMe9ER+8DkUVO2ZqGhd1ZX+94bPOuha8TdGraaBrHEqD4cxwk6HXeEKSeN
Z2sYlP32nQtyBjKFab45yc9vnrY8uoYPe6CwcxKy021HyCKfuf0hNxfd9tOFL6aARZOM8VW7D4ar
QOhw9mvX52K5OosihlsRPXruw8gGFTJCZsQbD1f+iDPTR1AVPbXV64hFE0fq8kGc6621sR8PTlIF
FVD/oIgotmn7yYjPKg27JcMARLyIt8mZg7zWi1D16uEEX9CVUhq01/PWTU+HaYyb14G39uJOm9AJ
wn1n+GFQVfFg4SFCN0eV3w63xHTiJAqlI0viYb3Ye47keUy1qg4Q1H6RDETMreJL4yep5TBIhonn
+ugpuRHoFFkoyCz+M3lI2GyCpVxPLKM5vbAfSjTEvrbRIKLqG9dKTTXwordtDdXTb6EcYnzSIlFu
6RrLRVWzsuKAtTvlYyZGbQZVGnBScvGWfVDgV74Kx4tlDCwHvHfZuLit1Gi/Yi3NYNeeeEJpUpAX
xfDJ8/AtCV7rcfaaBLqGwslovWYryWRbkh2zuazk4byJXgdtpR+gQj7LkoDIhFzEHcmeTZV7M4q+
tDJxp1xWTAbmjb/zWEuPebGUcljpOhoaeJ88/uB+VXddX+DHXdcdhXwXFBJXcWoSmg/yBNMyP1NA
9anlmlalbG8q3q2IrwsZ/0bfQJbAuWdM/RrdESBUzZn94OyJi7qyqTVIp/NC6py6Zky3CoukwesR
aZA0vEZows5VXXvg6/LaaFPVFMvll+cL5CEcIM430y1CsvhCWrEGxy7J6JcwWNHI8ZpclXijpWd+
CpCAB4XY0UFAO2qXKCwNOlysbksG2jmLywVQd1Ng5iIJhVECBRnaN1dFrr7Or49EFcQUMXaikiCY
ZYTUp9NrKDXh3xwsNUJNRWem/ZxCAnSahMvXtASd6Ww6Os9C+WUFwwsJDa8bKt6j9yfkNeIhWumf
GM8Zofu4PTwP/m70rdTdVCP29jITolnSyEzQPkuXmWL359QeShqHpMFiPhaHvteYHupr/YBNtFy1
eBTVPpIhMedo9Vdoz7hutwGl0I2p9Rw7E0ObJuorQ42uuj1nUYvVLCmltc1CVivUZqw4O6pbKfP0
/dqsxtCud7c7RyaXXrUK2VsOkZ7ByKlHh9evusbt8Ju+FMyA0zYfYlFfaojVJoqHH+QvQZHc6KIe
4JuXMfvWIcfFUgJ4RdrDMtqxsOKn3PvObPN4O6xP0nElu9ZEiADdH/S+lPyBfZSDX06FAfaG4ecY
ZXfOYmH9scYS+cjaYYU0Y6FZj9sx32+YkQyQ+VCIHDrOEB87J0UHmdiopkve7kT92p0FQt+guKIO
5Gqth1Eo9LjPwvX3BXGqJ+Og67qYQAVvDlkYkCJhDbJyh7ip4rAaTQVlv4asIWEVQT4YHrecAp8A
vjscBOSKkeXB88O0tKq6Nm848CAXva8brdTB7eVErvXi1FbNJiDMgVE0kN5+q/ybAQEVxHzQjzcg
fkWhqHLWmwhjfOHNjbjKGXoFLiIWl0n4NyfxZLKyvl5hkUvxHfnPds+Qm+JjAiGKjeG2XG3DTUxp
vaDiXBpZfpIHaluGbCYttphE5rrfolWwP/Y6BoAbHxmzmcqxv5PYYtr1+POH1YaM/JHZ2q/3BLdB
6sKtDf1w9sjwwqXvbl+RzSPcy/vOf1Drfed/gTyn6CCLYNgLfDPLiNJOodN1rojpEn89zQWgLWB4
stfzpld6V8txrnsR+JFVh87QT8GYHeOjlpvBTorsX830jS9J9lTZPFqd9FFOMxtkg4EfN1P9d5mR
bkJDZ6vHRs3QtEUZsAQu5peOMlV2UkOyCl7OI4hRKSXGKq0K16ETtjswRIX0YXZNr/wFVDWNXWbA
NaKNNaM8OulXpFtVDyrngIa8m3g1faKBBY5k2XMRpN0f+1SznahXC4Xpprifu2BCWeBzPuaAPi3n
Heu9MEMi7+FYTUpHpGPorKaAPUect75AYyz2fL+fcG030vYwNcH9fKMTrHsc1tEUjez8A09xZD+P
FgX0pRtV1xRNk/Udxt2Ez/RfpcnkF4VzCMSsu5pKsc5QfUGaeJnpthuK+pMQZkqBw+PkWzyKK+xW
2jSW91jQGFC3usB9WKqgVaAqbQO8CkZoa6OCE22zG0vQA0qzrb4B5/nSQgpTvydC5cTKcMImS1WM
PxC2DaUKTRgDai3zWZvLxnmmUygvQFaMxjfCoZjmHZSILlgOZLviXYJX0Gke/wgwjbkBhzxZWusx
oJyy8HuL3GQnzJENedXCtFNLpniO4eb7nFr5OivSdUJVTnQXH7fLmyitPuCJHVLUYjVmX/uEwulU
T2iBxTBOOisM6lAJCaih1RmMM5nXQaWzkzi8UcnESNhGTvSpwsvvae1M5QjBdC6dAU+do/4Q2bjj
UJ520oAx+MTBcdXd6ahNWrxVGBXtszmbP2oDdkkxhy+slB3thvVN27vaDdzTE0nxUf8ZEWr3/AQ9
aZZ8m8eAL+zAbbbzOosok5SGtHHgJVVAUiMESVpD9y1/EM/X02HtO7i7WdtI3xcq6jphk1GulhSO
AUW0hi7JINMgS/3aHE5hHonjkEjRCz1uQ0LH3FHGAdp+sSTMSzYznRBL97iMlE76cq4OkT/CDM6L
Qc5AWbEBDg7HF5sUHOaFgFghBF6Uf8g6jrXQitHZtySZ0ski/H0BK6ndUjSuCpmPR9b4WanFzfT3
Aru75T7l+mH1heD0dD4mZVwHExM9Q2dIrogzd1UN5/52cS6MrPMh4CxwIr9KxvqvudQ69THnD466
qUoLgVfL27fgyHY92e2nILCuECdnZfjCagMIS4ADJFLmvBfOnj65p5fytBadTWu+VGGtH0+84Ci/
yQP0fsSSlyQo0reZvZIAPqHBcmhaOivdHiz4QyIjQb5EH2P5ZFIbLTSxNAsdq2dA2SZRC8XMQYcc
jPE1IZEv9Mrqli2zXTtT+HbKOaGcBq7du3eXmmBPiBJMVFYbs+hYt1hnRqjc908VIMsXKM1Tsv9t
lrl0tLO20sxm/YWiKOH4H+eGwroOgp/V9kR87ZByY916YWoHqsY8nQwf0oUudbfulhbQMxZODgsZ
2lGB6TsVk06O4MF2NztAqRTWk/81KJd7mEn39xf5GsW5ML+jKjqewwfvvSz7Kgqw3YjGJKhPQt49
DthG21Gd7+v876DEQkXdHjsa4IXv6bG+g9HrcKGog+l4zLZV+MlssDyg92XPFh7g8qvqTfkfp+Fk
egbbRCDUYiS0KcsbufkBMWEbYOcr3GJQ//w5E7Tp7QqNG5henq0VfpkwcLgrlo5ieNLHfAC66BBV
WE/8a94n0i7hbswEeELUlbiu5nu6D72BXD+Jit+ecvVE87tPAV8eC4kaWiwOx9F2WIv86E3tzBHY
HssVk/A9u3eqlExlMksL0jYZKd4reWTGvrx9Yrudc1ysCEhQTRuvtZC9OolA69qCVJ1LdvRxU3Qs
VuuzKh+v3PFhOSGAohpVUg9BATFVDxys332mFHqCsB19tDvO5J4UmQQgMe5BY1TyTkd4YBwyUw4q
0LY4YL9zHd3dGw7OmkbtnraTwuVV/xK4hnkod/vCB40TwoZ+YK46bV5XYDe+r2pDZXY5SpS8Rjhg
DnX4D3j9m1dE13jVHO0KEfwmEOyE8sa+zZGx1DzV7rtOx0CCB17N7ErOjS+iiI2bandk7RAh/4qV
uj/0MlhmtADoz+4HgS4qrti+uteKOPg5AhFWqjBJnRofnYBWazOr58Bp5dm/8qisljOTxAeHBXoD
VAVA5nL++8VtHtoGK+dEe294Etxr0zs4SAEpuR2NNEkREpg5/2tzMKL6E/GfKwjlLIuhe9+BYWM5
LgCEiW85UqwQSX82BR+RZAZr9gGzzTwe+E+AS7wQ9QLUU4CZD/GMxva9+XNMeGkz9jwQyxsTVKJA
qlzjPT6I3W44iE0l+Y2A/NZclMK32H8SMXNr46wqOk9zTLCOA9oW2ggMhItNI89yFaFCEg8/TaUf
LrLGfNi+KnVAZGipz7GKVvdDv/XH1055JzAAasLWO6sHItk7td5zphURfb2veEXRnA3NYAZPbdwU
anV0UblUGIWVAy/tGQIrB9k2iC1yHJB7zGpz28Mkq8fn6RdH588CLg9kbkoL2ktFWV1rpnYcLS9H
DoE4iHZas5moR7kj0w3QmO7rilAhqMa3A+Jnu6tFu7ARHQhLYBclho2TXlPT/j+3oiFsRssmNSjU
XfCklLcjpqSSS1Cdt3WpmTha23Or9t+c5y5MJDdCYY6MZy2+1ZhDm6r3mj3L+bkVPzMMaH6TxOce
pEpAmsERk7geH2MRLoO5qv+Y4/QiB73rRONUoJNLtUKLfNYfEjtuY/rllyEkRpp8muaqtyfXTOs9
vvqMNmVJkJrNosA14NkAgrJVMaVY1wI1hdMmEAroZkQ3Rubt+QTC9OyxiR7O5UD6990U7q8ZqlAP
sLSQQr8cPdIewvjURpR7qrXR7ixgIjCKf2qX+HnBi90NUf7NQGxHVkXwhDAgzZq5Z5eBfhpkUJcc
j8xqfp50zQx1+Rb8W7vWQOngsyCFEElhUqLmjx3DIpLOx6PRU4wE/4kbXMngf9tdcZd+7yPNT/dQ
LMbPQLe0r+/V+usetkJ8trz047QjKst6vpQOMXcVHQXPRK7iSWLSQyyys8AD8b0dQGSww3KtJl/6
6S9PIc1IJvyOM7XFXUN7/o1Mv7K7ec7jF0XdFaniP3fDkW9NSEpdnfBHByXzk8QfJwFwtCdnoOzQ
2/fnm+XXJIRy1oarwgPeuemhgjRFR9DoBr5wwoaxvL4sC1GdCkD5RmP5tEVhF9uYuTWfXpQj2MjW
j8DsQsmNJsiKnlPBygi9c2y2O5D5FsJf9kj6q2yaC/pfsSt489vQjryUyhBAQ4xTDwG1cFyz1nA7
6+WiheAnOVyeu8gpL4voar4e7bPaSuHgcC43ynHD0SIfVfyrdq1HVylrsI850TKzjlzDmsv99gVP
PlPl5trz8ybphWnqc1DLufLfaOEg8nHV1SyD4l7V6Nj5QWoRGdJLwls2ep4QJTc22xaUJdwkAb2H
aRZEsoJ+Oqeyh3bwJ+zGU1lYF3tNoiXE7nNZGqj6U9b0xYIvNrESPNvP83UbslJO2iKOJ3XN56Hv
gMKkTTpjyCuUGtsJyxEbLWOoQNA30/RkTlUzYOO8bkjh5CSnrxC6tnSZtIq4rHvEsEI6Aso8zTMn
09N0oYQmjncRhxYk/TbUvqdPsOEoM5qrKV+DNlIMYKO5L3Cq00u50DGsEVSGU6FlyTLc67wuxDne
z6XUa3HBgs10TGaR1nHmkTtoC7RlWUcrNBnDUtX0p8f+nj3lDLA1Rh5pDQ0scX/WojcjvWUzRxVb
YxTgAcPtVvgfx5oWCozuIfj4T9+CWZUUgysaodlemKuIK0ljwzxVY1Y2h26IBshrpwnLZvYeZA1A
z0QcndMik6YrLLfIMs6La6ij8TYSca8GNDVPZt/suPuXFKctXMHV/lefE8xfHhVM9OSh9xOq+ImG
RswNbkIJbo3oSym/4PwA48eg/rJ8sX673dhCKVp5WjLcv8kbrrvloYkornfGen8Dnh5zU30u4I5f
2KqrtqBamUqBmfY1oo0Jqwf4uuOgNPei/5QMOeF5U9obSbQBX4NvODDwwtvz/r2C8w87niDFtpve
1ji1hGSH/E8uyt5iiJCogF14e8y8T/Pk9qFg1DI0fTvl/SwDRUPiGJOJv2dscuqAzymrIFSEf/8a
iMxWFwn9qv77uCWo5tcjRwaQI5ZlgcGbucrnrQkbdocBbGwmz5ujCwZZhiQRigrWbR38jvgGbwbf
mFDn0A/O6ikgVF4bp5IbnuyroeEfMcp+BEWaBpirdcqhAFgrxM4L1e+EIeN4g/q4y5+VZOgOKR21
4FbxD9aT1NVaqhzI6CBgp6qIOUIeIBieO1PDPNShH7WLyqBKBYNBkcESzX59WlCeqBobbLCmXC3v
AIKVW5K+ctilq/hEXEOjdVQr8sGnLF06LTywRWrpzHV+BAg5AOMqD0WWcKkUMfIMe2HRkzBhmHej
ACfCiRH49YkDsDTwysDLikq17BwxfwpdCB4KNx0iZkRr3+GIi7BiEdbLscQnTanIVuAX/sYr7CQz
X2x0NI8sakZDzvah+qjtywSyJG8lT8+lyL9TRjZFkgNuI5vHVKrNyCx6TuXHoPUpS44Wr5MRtR7V
fpXkxNtwhSe0uREDUei+kWQjMN/ikGySD8NV6fbNsxxLbbO2UNXgT3qQpVWsTdBOE2BVuU2dBpl3
ID1vlEHqKci772a547X9znyxPUhUDBHEqsO7CLO+s4JvyzPm0iJQCKav2vLpFeyDDhgDgIssklRC
Z6UbLRaCanZaDXa2jB13Hu8lI2izY5+lV9bdrs0Edp7w+2E+zHkvm5y4ErhCXPdddHX0lxaCDIhU
/jM2tvjoVUs9pmAbwX7TWhCvZ4FG/oJYGt52uZPKmFieQui4KLxhDTtC32MxTt1I7ttPWBO6rNWI
oDmQSKZbhStNBP6Vgq7xiUDm/2KBRx7+j1kRNT5M4MRaAKeG0s5+tAA53aRPaKJMApRyWYwAUkv2
MMiMv3TnuhOhNwpv55uzIYE0X/vvbDiPPdFXOgV+ikM3wFFX7Wbc0yNvSpsBSwlBY0cZSp4CDRvt
7pOAbFsOgOi5U2FKO3ZHmOsOf5eyQXQzlFroqsZWlAX5eoi2hVtDNqOzYsPjom9YTD2q5vsSbSg2
7lo8BvwpwrceSR1qoBmFLS+TP+0tGk3EXJiVS1/kUWLW+D83mc7r5A7yOQm5WpZ5RnbHR1mH2hCh
Q/zMLkCRlFxIyUSbOQ8MVx7QSf9yyNJvrh568K2++xcwrEUm2OFVwSk1jeVOTWTVs2XJRF52PYu3
/Yk9LvOh+XPmllRUKKQCdjdBsMx8j/Q1te0RVhYBLm1llvutie+ghXco+JES6QaaY8zN5ZCYOCMc
UZVHW7XzBVbSaNKlQqJvJ1cyFFTYDhoN6I8UdSJ4NCLJ7xhKMBBF/aJP4wXtOWitqnC9moAShM0B
MpSnRLht/qwiYcv6SNHknu55OZuliCqdUEdBawODaTMNlenZgNdpuS13raHIZukZZq8PZAsi7J+i
7rrosf9HT8U7S2MgIP+u8WAqMbxkRqHGihJaoIzy4oQIdjsKxPZ34uCNyhHVRYE3N7n+SZuA6+e8
t/oMkrergf+bQAMRIkMjGV+hZbCNSBNW3yzu3Ew56j0RMRFNjAo2s8+nD3t9CkQEYmDLFxQd7d6Y
QP30Lr46ww/aXNCU/FUE7ztlfTARJFCZ1rf3kYy+JJPl4aVPDDtud1BiToNEkZY5ZnjyTx3u+PGw
Ef+cim3GD4E0xihrfcCgZ0R1bcAINE5ONXA+GkqNwtnU8qDJR92xFPqhYrxx4BQBgc74IMUmeFu0
YF9O3HFsUx2womEb11Z7CPVFhWX3wRpUI83oeeG8BuKKw3DRMCIRq1WwQFjprTgRkaQep1V5l1gf
87EYpaDBdkqQq8zVqO7+uXAE8QLlVzAwuxhc4OPf036UUigV7bPW46cWY3vtttG5QqNYpYTVJa5v
npyJYG8Mj81GdTGGpN8xJN76avovQMRaOVHpW2PREov+qKgvrooPzEUUwg2g45/TItjDhwTPV2v/
HUgDtbtne9Z5esf68agMs63USTSinMHhPEEtDt+YKIagEbVSOar5n18DHDrSUkfspXKRZPPrDtPN
nNyzuSrMkPC5LWc0h9pSqyIGwqXf+WlKuGren2rKO49E2aiwx6LPREAvT0XFJiIP/CWYt0T9d2KR
jLncD84EFrr6q24j7illObOeoIF9+zfudwYfN75SAsJrfAzt+ldVkKzScqYdpdDZga+ETpTGzSiG
GAfCdzSWykilMJyeGn6k9ynohMjBuUTiNytdETp23g5kQvzsmH7X4HGCDrnZx93YPhnn1jBj2cya
peW3cvDZMfRMCPZNddZoNXBFDSt/cTZ0+q+1OiKsKz+ZigXb8fxr92zxRXCm8iCIrluv9zkbFqef
UnHQU2+CUPg0YzWR13+spj+jgWqiCLJ42/cuQ6WHgcGP6SyPKHsPGyBPGy7I55O6O4Mf5BMYM+RL
eWgGOPKOGmClGlAkJ0uPFvo+HJsAOXABfXRVP5I+Xx8P0htBlgUI7cHXyh9pOx1HSc0t/yLzbzgM
pooy7PAqoGjl+qulPJopLpsBcWMg4u3RKVqe4KHegLZi1Meb3cXlizj6RQeSgruHVdNoPZnK81oG
jg5eUYeq05i4R9mUF03yVM85+jXjRmUVJBAFZzSoNh/xiOYGwV9ZaqDxDg6anp7JtMvB5KaLKGhw
SZTJ1tL71areiq5EQdcnfk11qzVZcajdNyuk3Xfn5N/T6EdyAvgkLmZE1A79cAImJda8luVs5qIm
NT7BIKXMXKEJCXYMoy7lpO0YWqgkW5G6FvOynt3lzWVBO9iLsXQZYyncUC0LSh3XG269jg8jqfha
vYJOBph2HTygQQ7N5Ra0u+aRuZcTgnplK0tDw2vQDuJ4ZTC+OJO8kue8FaowVnsM5ED4WYY6BUPe
BOHXfTzfR536dfVLESChK6T7m2k2QXTZ4K7Gsn06iXGCmOgpuCwAp50UZT21hGDQYa8ZxDG86YIE
M1HqVug5ZkdZnXlDNECYHFINxgGbG4b5QdnZpQj2SVZ2e26ce2Of3gUG734Nw5sokG2Mr+RDUIvb
bXeLanPDg014AHIxzV2aEd56RMl/pGoKhaTRaJgxmwN4WaxElcOySJun+5s1PHShJpnx1ap3Hoy3
4E6wlYs3/ezZWOWjdYmzS2PKq9qHt/ySmQ4/rCGZooot2Pans0x/dnUDCm+FkuLw2Gu7Ejz/qmGn
009hc2klWIYJvOULW8t7YYNghDKSRK/5Fk+7omy39yfv14BagdRW870g+G/vAix+MxVjXjVio5nI
AL6dbYS2yp3TNnu2xk9GDXygqDH7rXyMxhgESsk6ykxCmUJb9C1UopsV28sfncInAiTA+aZGVXfI
0HLYvEFURLA9mdWVZZdb+8CJaTZcheF1SC87qvuwEKUlE+vEMTutDAVv79cSG+iyRdZh+szR3Pny
Cg1vmRAdYNChjR3EtIjTPJyCPrDZUaYCdpB6XWiwKsi0RCmDfdNZw1+VpCwz45upJG6PL6Z0bWrm
9e+swRhCRjA2s+Zm6qvKnkwYfofoBrAncFA75kFPZhhgV82VIDgk4+4w2RlwXtGTl9Q4JdHCnzmf
JaBRZN1zMuNNwPqfVU6/ASEYEWk4As3m95b+txdWbhmlQCmYeNDpRvuU7kwKPWAU/wLqLigENfaO
3aWLOvupyy4wj1jYVvLOTlNB/tBrcC3IZFIAerFIrcyWzGYxeADYO6hcckh3IgZYyoMl+/bIhV+1
FLAbwbZEdoAHW72a8OxT8g2QCZpNAPPL9HNj4jWrokjTznYnK9RICtONBFTP1rNxAHGS2Uxm0mFb
8xHkwXbNkvSGg02o/KnvH8FfysHWuD7J3yJeBqJKmyFZhPuw9PEadg3at2hho70FhgXBOyOrISDi
FUfS/2bdoXR5bFIoNVJpWBArGwsAa4hlD4X0wJOwBZOX2YC0JMItGAeKbUwh0ujJM4Kj8kBvCksk
RAAMPuo+yURT8PgrRhu8YiZFu/CXfzZ8TgoO/+TYL7UPo+xWHl2/ePSNsAZXEaW88ZunqTbZwcI/
gvegLR419Us57J0LWp2ChprygU5yEC5i1munpQGI4nRmM0ZAE1eBishoFKZiC8dJHKBvlk2iGpx5
FEqzJT998vILqG7xoDwQWXeiv8xOicNwAxwzFnNx9qrFkOfDO4+BkjUcOlK+JbqOqqeGUfXKd8UK
TjCCkEphR1RDA5DXX0XWatSWammeF1cIkpYOTViMrj9rO0XanH6Is3rA/ZlFg7DGB10g+NBKsRjm
4dGb1WpuYnQ/Qb1ojGT5Zo6sCcqdG6tpSh0URuJ35y6clZWBhmfTYrSC+TziBjQgofF8Sm3z8Cqu
ADVWMI+PiBz1RuemFvDyFZfweJe8Ukrx04X+tFr/7IivuHLDfK0hBzXE1hsb68q2bKidXf9IOdZt
7PNZNHCrfBkPBZHXUNRxacYme54vtzoxR41KbG39spnISYEcdpSZX50mE11YZoFWJLOixcRVeOrU
UDfTEcqQNz+APCLFQezV58YEJl86A4WSjCBYF9kKeIc5IL8BrrhXbp8U8l4OR6lgyqv85BqJ/T/j
oN4zciIb79mg+4VF6WBWzdPrWDQ7hFMhEDxBb/AN7EztqASSyHXXtQkAXZeZDG2IbLbcPSnBCBe2
P1GF3iu+nuNnyxcTVSw2RVa7gKr2tE/LEmOnTEy6/wLLC8+7GKD6mk5BqhRamEtK+D49urbSrnSB
DSn3LEOYuzLUk6x+YbMqX7vG+2i5gasnSPdeSVOespQY+5+DUjlEBaYZaJ3uNF2M3mqvXwlloo0w
eFbjF3Q3In5SbtBN3f82nZMdt2todVVtuyL6PQIQzWsdd+42MsddKDhsJRqKlky0y4XhHrQx8Gvn
XsWMzlVw7o3vlpbbZyWMurt+pMmWPFjpQcKCajeAB9qVaQT1K+THUzHXIo5YqVpApdC/c6aGfg61
3h9NwS9Kcb6Z9fUdyo24Dw7hlvxLoObcmiK/hcZHQ0pYzj/3oSeFz++vYSeWHlQ6bKFha4DMLMb/
yNuhUIJGYD9Xo3u3enQtHeo8Pv1mP5bOs8vQq3aXoAEjgHP5/GMlQyOK9WjO8mY4JDjSYCGYd2u2
dxzgi3yLxOet/3GLqRVMXIdftdGIny9hCtGbNOADy1dI2V7Acp/pMp0sShpVEOurPG8MbBA28Il8
OVKRUddZOYfcrRnkCfvBPCr/SvduBjILcryl4B8wEOD/gVHey3MNb3Cyce2N1EQD1dVv9iJiNZxF
NnyJU9elZ7yAHiCsH1NHvc6Sb/GNcmJiA73f4mR9EKa9K50GZUjhZDCK4lhHLADevj7aKezAFmcd
HkdZGrOeJ1/XMKI6wOKBqNnPmidytDkY/ZLx4+3TVfz/dsu6xHWs7pkrnw3/tsaA3bCdWYNk0m8T
Mj9BRkDm5vcagF1cRtcsAYqwOX3sRkAo9zmjMzpw80ogCVTdig6jqXDqXg71KjoglrJgwd5x1qYS
zblOBEBPqPBUxjWKEzU/k8ivdeam/UKHxse0GSiXTG2LB6cfRp3neSbDUXnHfdiNA1zq0ONEgfKt
xNwODYD1Ha6DMsJAYuGnkHwEQ/vAtSKWzZCGswKizlzX869MUVCNUK4KbWSO5uDSBThfhLeo4NtT
a/zjS1mDXVZ3w5oma4A4wjbs0Z41fUtgyzvb34+k1X3y1xBJOtqtpibP1pZRvQfOanHgIhkvUgYC
Y6+Al8735W1fyBfNe4eJr3ZgUkKcsqDan36u3HffN3e2A+hnrQbT73xbtEEYjZJjGUdDYiASceJ5
eA9JLpADqdYBpQR+vEYWsY65HckXa9MptmhUEZ6S4+2iXiIpV2HJWkgzc3L+fDF/nQULBIkOOt9F
isvhYX2J0CX4n6kAtGQ2ypEf51QY8H66Dy7h/D3zGWNlyadwUOD8McFyE79kfbmuE3xy6+VaNNrA
AKQY1F/WeIrrLAUp4FIo2Vn8dqWuVMbpZYzJC0Hj86vmL7EwzNQ2njQCUIHh51tFieKzzRDvZ8j/
tQXFoC0J5MWDtQEokt6Ma/CPiIdA95+kGBzEPvu4PJx7ZA0WpIFy286SYmP/31vPcv9ASn7KDni2
xyYcPfaH/MYVrMWMhyE6TJ1Q3eYr5IsBHeK3lihojCljFpPcQsOcQhtgntgJ4bmkQHk/IAf+cwuX
jWSUabPiPSrW+XjYbgWzopDeVDjlgZaLzkBeihtWUhSox9Laz6w9HdCyoMFu73VqydiWT8kKcAkn
acBgaeYems6AV7e4TKaGCPbZsjhLnhbjnHjSkv3b5ugvz9mbAX4x3/xU4H8LKlba0HgoD5aMX7G9
4Dn7DBF1Hsg9XPAsvQODR30HHrvzOPythyyoPQg3M/HKcOkxPeCfD7IuNvCMjNTKYECGR1AqN7Xn
FyNTK5F4I0c7rRHSJaSWC3iKzSu+PGAbZfQUDRGFJVN5wHKjaJWF1BacTITc3d4HUQDgko38lVTw
w5q6ymcNVUN5ust3sQDSGeqTxsIUeJelm2V8ah3uodrFp+KC36G3VzuQJrVQnl0oBBeCcVHgkLtw
HA1fN9gPUUydbQMNy4NwJDWl1aKhrFKRuLoG0CvlYKTwGakwUalugqE2uQRlcIfyl7mfILIzOSt9
0yuTj+GCzk0SBlAOtOCSyBHuVC/3y8C8zW2UFMPC41tXtkqCx9a2GLYetB8TNNg07xMeW6whs8GJ
WXz9evIObPuxhxiKbLKo7GcHZoWReuJ8yH/67/F3p8oROZRdgvCXUA+MaaGEquNzQZc4Um1D4LSA
v6KxrhYQMZzk15UDSkfW1lBH5oN5eat5UaF9rmZljsfU3fQYopiAV6RxGivYXbPdNkbjAaXgX3O2
TY3TgrgUqsHwwkvZp3TG5Cfsil2nUzQC0yH57w+zA5nuv9+IFDOQmfzn7qoNDG0+FPnvSooiVs4L
GgpNzSxCazEA81FoYRqpLx53pzZEtKhGi0APkSKncVzfA/3jttbxU51k6naKPJkxjtBr61A9ZwwK
TwdI78qbTfARTZ/n0bIJdO7suLKYvTCf9g+IcNNHW5ulLaM9yFtjgXZNfbwWpQ4+HwC81zTEjgTW
i/eH6kUFuL6cpYDezovKfQyScLYHUaP3RDMHneO4faj9jDprWBGaWRpCUMwbpKkPYGROGuod5tHW
8hdcdUU1SwJ3IV6KH1u+fp5NmKr0b3YEDGl8a71sAfZZC+xa7K7NEDv/I1+CE5mzsdd664wj8/Pr
i7GBVN2HVENDaGWw0lXQRazCrHT45xQ/EN/dSzGs9FIsC6OJir8YzNdcfnyhG0bRs6rovi9E3Ald
v0FgGOvbfLaZzckIadpxJsgPT8BELrIsvGKKEc11YOOSc1wD3aReNs1Qr4iYZxKQptK4iZVqH8ym
uSVCOdmSlXcaYVTb0nOaCkcuTuDsMxe4DeuJy7vvH6GucVRupml0taL1DmdUWXyO58xehe+IEB1M
pV7y9kM5a6fKh11HoCP+HPlUHGBQRu4YEIq1TttEic4bnbNIcLLeBv154fEu7DGA5vSluAUJNCyB
YISWdmmUVYURahWw7/4OJKtNfJIKRGqziJ7RueSUBJ2Hp7P71HhEajXZ1EdyR3Y76ZRMFnvBzLx5
8YSgcNzWU+n9PN8akT4Js+iiUeJ6WtXVF8e/fk57CXGfYgwyp4gxtz6HF0NOGrInxUeEcgd0Ct3o
XfIrlkqek6WlhHMaqz8MX/5HZIa7ReIvwcbIZ0Go4Zw9MTTrDSEnD5Ds/Rc26lJvvK9Qis3RTOG+
FOKySIGWjCNRM8nyYirWMPiwtLrYzHpqiGyMwkrcnxTTRiGKZ/7i6ec+gPV63MkTbSqPO/sTtMRh
egjbl8OMIIrZYSFn9Pm1GYT4igC7kUf92AQjPS+bomA1e6RS1fONU7oZv4EtKGRYumdNoo0dlLSu
+vfbThbhj1OVynilMrguymXdIHL9L/+l/h/yyT8C3XtJKj+GXqOdTvWxuHZB0gZrvdgy23oPgrb2
x1JB25610IAbDdlMfoiFZz2I/qgHR+zTNqoffuTUNlRuUyI/Le+W/d68bHHosqRTRfiFiXRhCtUe
Zayz2atMMdDDhXpK/vPdpdcn4LEdOZnOm9i08kkz2+FSY8G/KRJuDfjKMFxI0sl98b6Y7YSfQtWr
sjUpCeG4A0qyI+17lk0kTPz8fh21ltJ+It8vEY85I4bRDAzLD+T5o60UAsMuJr6Vdp5Tk52yjqqA
w1+y40C2m31JWMu3fUz2Z/f/QSxrfxCCd9mDLCBKguFEBzcckCSE2YxE3zmNbsSVGbmOBAIkFAO/
ZJrJixo4hSeatCTQR+exX/CYqtnLKmlR433vwCjm9SwObqV8/HEIjzU7s6UBkXTFnS6yja8BHsk+
1DYkAEWU7c++59+yeMhFYguTdwC/vYwAZHzh8DWvXwntnNEr/RxaDAT8xRWhKOvLQSfRL2tEioTi
IpTR9GLvaP5urKPGgw/pRtye7paf7ZetkqVD40AHwNl9epBiz2rE/1hxMJtCRTsjD2en+XAVawv3
wOgzL3F045yUYGhOklXqY1iV4fHTT7Rhj1Sw2FNvFRxgDM2aSS57ZQ6W8hPL2OJroyEEIC0GA5of
SgYJQvAvSoi1Zq5Mz+GoNAx5v5IIAumcZiQGjPGfsZkOUnh8xHG0OjTkdoQj5WCxAYqxJmG0VNYY
h7togLQrOSfNPFkx5DwdH5dsf3BS9/uueVxJptaPzXkIyjmdIO+zcK6TC90ssO4yCGixUGIGGXei
8tqMR3WS5wqProXXLru93d8UWBxBtTGorqE9/EglDfq0Bv/0Ar34y/gGJWGpXpwStUnW+5t31l8x
Ugtd4TjVKPALd3PbHHiIzD5BjFwkBNdNzxocvTfhMAubrSV86Sd1ilNB9ZoW+t3zoAAYdnSol/M/
BZCVMW5IgBeDPscIOIDw4oUKxa+l0eqhEI8cY+SYwh6tep1p1GSltKtY9YfSKti9Gv4rrvYYeeOq
kcYEbRom1O3lVrHJ6tEm4vbHRjAII3DoyImfYuuhO0yBp4ESzcIcCHLi/j3ROmLPLlgPF6onFW5Y
mmlVJ8IKMsINyFvoDOX5jFPddS9dgejy4mw6vBo6FTPdWTK1OkjhCNfcXJPU8gYy6/fSh077vqCC
I7ewdA1CGS9YbKZNQcEKDFdnLz2g0+/wMQSkjcFVG/n9WPd5dwpDCOuAY7mV+HIaweeeThLAFp0S
r2Xuuf6DEN9bBZE1HAPz9pRwNvc1IiJy0tzoWRrRFRKDZnvPe8j5aix0KisqnoE9PuQvZeaVCcEP
tTUp/KePRXJln8RjrDuREtFp6kNo8QWFcnIekihj7yIHziaYyvMqNIr+VsCIfa8MuI2NUxVWy7Ad
ETuw0h0l4dDz7/EiAHA+YvocTKY2iX5gIlsqNnF9MA1SSI39NQT45EMcA/BGT8vFSaBU11DwtHTk
vjGzNQaUqmz6FJ8Zc2edgEH+mcS5MHtsxKo5w6OTkGk9oEyP7Yto4lh4advrI+4ZuilCk69WZYIT
MBffwUTzvtSR693ZZ/0Kosb8Hy5vKQxK2J8LKjRcCVrcKwo/8m8iHDuQUpDWqscDND0WEOf4SoxN
PNpcCAyMdDz+1NGy4kuXEQDil++09tuJo4JvkH569rBk2i/17+I9YULbGwcoWoz8GeaMQzMSb6Sn
j6t/7MbRcluN0vH4wuFrp7sPLP0SdNlypn+4O/gPxWyAQ2N31psjKW2ymCVa6dRCRA7v9DiRKZqD
2IIQCOWYcL31RuaBUdoTj38NmHRxTbjJSnlPVRwfSvZ8o2EygpcjM4GyBi/+CW2t2wKSqkzSg4AN
I4477XSPcbWAJgGfTqOTwHJE7K7X/FAMh5AGZACDkTMeULnvJ8ph5aU7+TFQjIO+x6/kSDF617Ku
EaeBxHwqFcqSWMirnl+G0vRCxFQaYcJjhlKYL7CczfMDPRmccRibKUx5MpoSrWolpdpepOTx64rY
w5xTOTNZMDpm3ZmnOijpBvd1wPwbPfKGyF/UdeBaiypJgjo89lMHK3EDAECEFn8gZi27dlhXEnQF
4x1CbTGee+/zYkMQBI0aaIRg7+uzEZbteXQ1Z3NSYznD9oBQCRnHXD2cMYnqaFr8YdgVbQ2GcKhX
mkPis3uhRvx/SQ4fcJUTIH6kahmo/z7F8ahUVN/Bng5llVJWbKGG/tkvuBksyrmtm8JmayBF2AgH
LN4CJVXfXHgeQsDS2nYnWYwaP6+vBijANPYP0R6YshWXJN+VI7YLGrNkAZBGYw2nG6Xj/fJJoi++
pCc7GUfWS6HtjcOltks7Wh7EZTX4eDHctxXDbrkM7KX2yVqT7tatsl1zM2Ii38U8a4vQK9Eb0HVb
gkP8usX6C6lhl/hE9jiVOYh6lEfGiPzo6JKNRnLkjR5OJs8sA5uwJg92dSUHaGKvWTQz96EDH8WO
FhPuWBJvwY44MoewAB5p4AYwP7JzmTtQ1sby7JAbDS0XJmspvEOuA3YOSlcpqrSxvo3GfcRsHvr4
CXVk88bBo/9llS4oXxacatHg9IEdjD1XNqs6Lq8bUNnuRAMWuSgMa+BhCtrZzdNzQlJTWZnrAM1f
MVasQqZGRKCqmteWLD+IktCgD8Vg7XFgBIv1nxPC4+UPt3RqJPil8sbnE5VMG0dEkf/0gx5qnV0B
aL7vtbg+qNz1tkweAjbUslVe5t4s8184oeuACOFyhUeCjSgxdt5wh7498GgQRiofkuAgxKq423QG
X7E/eSDbvpzgKuthSHzhf9lu5ZZQPfZHkGVjahBBJGXAwAh6Si+IaYDSCPGGzBtqs0hOI9tjhnga
3v3cSAApXcZ8oBfhToX6phQ0oLZ4i8Zpn9lfcdlQQMcgmNNWXA3joIaADWBJp2C0YxE4noMvnDJL
eLMCWlOOOAZqWZUuW2XGErtJ5lM9R+Q4rC+lRVwKocWaEyJeV4nwmGSliUCAR/e7Bqi8QCKB1nHv
Nj2A2jt/YqvnfEVvfzLp3JrmygdSeTHXNebD4OqQF/1eecuOWQTi9we2+aqFXTMmgUuhLq0iCKHh
WbBXwjTaXhIo9QU/dNdmVY7UwldYBpFHjUW4O9ZhJzzr/4Lop0DIHX7Nsf6KW8Bg1oQK1uDplwMe
7bPGkFQ+fOTHoJpVUN0YZITln1ekWsQsVZ2pPtMndd49Ky9UxqE0yKCBgKX8qypmXSLKx8BuLpk4
mZ8u5Du4Z3sThlTyFZimoOeegN9QP/MQdN1MjwgOswHXvmBZQi/sh1Fm3OAxjlm/CxXjdRJlKKkf
is5Jy8gUPfoaeALEUfmC39WyvUHDq1chEL9/hcu9nRRJd1ZsCMRIWSHURjpw/neFwtDmTOj9qr67
DUlr2Y8ElKIhua0M9l0OyHx+ORaCNtASXSwTVmlXPegDngXWKoIZ2goasKC7d7ihCLF7aTfIX8gR
KaC70maMtIdFqRuKNGwlXCGirSZjhuWeHmnfr67gffev+KZdWl9ubfFn+ZqdnqEC6VRpd/Jd1Ml+
LNvjzcf9hH9qkzjX4HHGIHYWUOXkC9odqhV2jNPnTfYe7vKw27UgcgBe/icBSg1K+4PRtBKLVD8A
Zhq9SUj5vf067ZZ5rlhTGpmk5VmUQBuZy4i8GF3bo0cfFjiNG3C73CvJK+sL+8arA7eX3nEBkFz5
hp4KvdG/0PZlih8Sx3okpNfrlW+Rsqa133OWsFjUbx/NTl+wBkG+PU9f3QntQMJfQjytLXuFb++R
XkIc+nkLQ/WSO/iQB4i7MH0AEhB0aWcDB+v+khMfvCwBiZcR+wrMkpM3Pc0N3LnuZaTXbVBz4o4p
Ighpvkg1pNcuVpe2PlbiouQYTnqkJnzxh7bDQJnTbXSlqErgmCiurvG8Uln7ECvoUx2bqQ3HXqQ4
TElvkyV3+tPc35F2Q7fqUVtfSIbsPR9dwI8c8J4geaSh3hbqorzOK2ox+ri3VKAZKXJG9utwL16F
V9TLf6JaMXjWllKcKzfOpVs4PEIXwczFa2K9nXj+v10IK4ofCZy3b95JhTzcWqVURga4OHP6UkyD
ZMcNMtvYd6Hfj9XdbbXIHtLjTXcPox3hXwsZfSi44X2oJ93/jCZauUNsPLVWOyecqkFcF0oLB21O
o6JA6PvLR/PysfkjQ7ttkwBampL5QnCs8bD+mJ9lXsfISuPuMGkrnQvoN3gMpIrArnnWY4ClkvwX
Bf0ikt3UEIMJkTm6JV/+TsYyZJGvPhEA25zPimpimwpewCLFBFvrJ5cIz0bfuftttylL1Kkqh/4q
2yewb2nvGCvheC3zO7EUslskexFTbpVDRKTPsJIfHcbdyU/8FpCrxE87hoCh2e9GYJF+8X9NMeX0
II0jui258FKzO4uLDPbUJr8+cWOYf8fLc9Dw64VBzDANZIeaJC4pZP4agdQTrpdVizB8yzRNjYgs
lEV95q0EC+c4bTIMpxAMtD5XwXHpNtdGYAkMHZSlPNrZnv8UdY25XdMsfPlXuhmJERElfjrfESI1
SQVFI4QcLYGdxerN3ZE92kyMHE/L3Xedwzh7EX1DcXYMz39epjb1QhuIqzo2RFVMT3CuH28E8zJ+
h0xWvRRVpRF/bitw6Vi5eI6KWNJUx7qw4HDiEam9Sfc54IJyDw0e1w5GrEvH9+2kzR1gxWSHFgrC
GrSyzfrTHADNHHxCz8di7ejX5w54/Bc9/ZIAsWApG96RKwA4UoyB5+rBmhL9uXvC3mI02b1F33oI
8pKLizpmhtPaccPO05vtpdLzSxRxG/D4iJZc4LTRqE7xxovQ4mw2ldtVrsZCfqRMiPg0UrwagiTc
o7UBUNtg8GJxoK1T4Q30YNsbFTnW4Tz7FyFv7O+upG5LJ/5vyeeAFWXDYjaBWVRvjyESEgl/Kv+D
ChNUz0GzZ24Li87avCTzkq6ZojxlrM9tzlY78Zle3+CQp5qjMJMP/hm9xOIkW+t6pL4cjiNrwpuE
rHBszFCE7RmJDGzKNw5rVeisSvi884zKIT2kyPQ4Mztez0TA6vTmbW7DJqJ67n73uKKu/1XoOVsY
25ZlkpBpGrIk60lnCYowIRqQ9VnpigajvMVzAGFUEacqBDZ4+68i9LKBZk1UuSw9pwzIRuvdNYGJ
GGWL/qCNfC6+rRjWcfVfCEHxqZnDS4HPy5t1v7jZvahm8+/WhXbzbOKPn9n02+5OGh5FdFXjR3Sf
YttRN0N2oJ6sNJUG9E2ZNEK7AuC5x9hZnWVRGr1YAdz4J86Mz+aKHhrn80oTg2pMXvh3VUgC1nUx
LBcRmuty83ev/oCyovbce+iMKp+GjbXKXZTRJWk72KVm9HxxOlPBoP4H0fR13xENIns7FfSAoxIu
sruESl6u27U6UdXc2Vp6hsiP675S7Lkc4u8Bvej7bdKUTWBYb9GYybXVT1HPiXEDcmyedycXdT6a
yK/8H331Z9Lk6HVGHAdsYTxcReZrDGf949q7o1CrbJv75uSbijxk9F0N+/eLypp3tEyNPvdIJXN/
0Ly4p+DsjQhtRhylDg/v/QQb2xTa4NKR9HPItFrEGyfsD6bV6Sg+PyxmSYJMcq15bkpueYV+AC4A
qoP5F/xOWWqHFZwLz9NlVGYtIG2WrpgMxV3jT+++yNWjdNVYluQaqxNC1O8qyq0aeNxK7abE/E/z
bQX8G0kEKmGRkWTkuh47p5T2lLPCc3V5SBZktvQT7cvhh+hTH7QzidxkmjEoXvefGwE8nuh6jReI
uhbeKacIJHMMfZIDM3e2YLjS2BGeL0f33YAoZx4Zjgl7KP26VTC08FW9UeaGKCA10emulibCGiU8
vHPUNnbo5SF+BftlnCQWeah4adjqyyE2wCgJUvesFmNDkp++DKBF69P7M9AWvP63b8ec9zwtap2a
a/5xANxpPiTmgpfDYc9NSTqz9WkgvBF1YaYXssfb+SDVD7JeVBCuUujKt6G++0sUSLo2CoIB1M48
jVt0WeoL+US/pK0mHSajwbj5LQX3ZdsbKm0++wl7+9IyHD095k3J+edjHTejwPrCbEzA3QwG20jm
WpAOJTesnluV8FlU1dawGMDu5aPrq+8Qq7ETu6guhTlWU/vMCtvBnkKoXcUWreCbVrUU/PKlp6TY
XTRLA5QKbK0+nemHPxpD9IqOC7DX/dTVXYP5oHWFN91tRY92WECDmgWRY3yQu9jGM4+sStOmbx1n
mk1jJZASZolPxsCNlEM3EDovJb+/wriMSBaqnW3ufgZoO9xO9XKYJ7XhsXWC0Mz9sSQFn6WXamdT
UgEc34pDlkJVhD/r1nMZe05MqKT2+IYqQZzDtwCGunfmimgQWzdB18PFq3Rs9khVUsEdDSvd22T/
0/nLsIEiLEcPXc8Y/+2y10/IGXmspR5Bp1NHArHAD2n4K0TSxk9Ruo1vJLymu/mecDtwFjglIMY0
hzymovSlAI/ZiWaJLiZrczt2aY56BNzasSAtYBC6tK9b95dZrryUWvtMgtCGqYuf4CFWmzDEtq+C
HLMJqdoFF04hVA9RY3n3uddxbtTdvQbG8/dE5AG1zAeZn/JacwWpdgeF26JWHAuGKs+WQvM6ZuRx
j7JrdSftInNG9E7macO6SrMylw1YV99ZK8HLWZXLlR56iqxFzKteE18aRS4Q8cR3PCK0uQRMzRKr
FZcEtK8dztIuRCbYETRo96cDumVkossDFaP5C2Ua9mVnD2/xHUJuwbt7g5gHQTJQ2ozEbU0GsrTP
ftCSPKbKAasJ/0emopMFQ8vnCt++bG5ylzbRVfWjdWeqhEUmlFtQ39KjNU5xHu3A3fUrA00xCgGf
x+YOY36xAZ9EBNGFyutcJeQOKfsA9HoFi/mErr05bzWbyYoXKKzkUF97X3g3ODDhyWM/6Kg2phmL
cdKzEtBCYQPVhMf3jew1pQpd2+7P6e4RT4PlK53wWpR4Sp3jz/GKYnWgD4wZ9ofmuTlc15MMBwrN
0E9BZ2hMcMInFjYAbybMgrG4FCygvmEc6AbZu04iuvp9ZAJIdAphb6bEO26VnpJc6GDb7r+SE+Zf
m6D5svTzzVeumsOG5l7CJpHvAQ3ZlwRz7VBFgvjt4Z49+7qG0imOf6ujvsddF4TbQ/8tkzTylirS
6bFf52JQpwgjOqqUdkRzjy4lOOmktu1zMNBYSVCdRouROUrQzHwqmyBKkJ+XbrRNHsZA0RC8VgFM
SWfhoONgLPxlAYvtYV6fjByNdVIOGJiw0l+lYBc0yfwVSAygredXlSODgyceBIa6Ke6xfopsXoOx
sG1I8mn4HGZmOCLldI1js04Br9gKTaX5vGr0+dxQrMZhzPSdRKxQnDus4BYbp7dpDH16mcbJCvHY
PdflWfPpP0GtmrJUlNk/fRdbWxspsjKws4EJKGYZzqNgYcwt2efSlPVmNVrCw0rXXJwpTpo3bCNE
LN+0ab4Nvv904LVvywjiP32RbCJYvh1hp0uFP8QOosIwYOon2CNabLj3sE/VbpVHJZtfycyCQdQl
Va6RjJCRf8fSMvK7C2Ac3+HT70ubZHjM1ReuWyaK7On7b7XNzmYmGbUDUE+mVw8yqFeYwJXkkaus
urjS/MA+23l83NLIi5KmX/JQH1rZEr8Jr+iOxyzr4X4XvQJXiqFbngLAubtnkoaSNjJ8CQirmVyY
FlYPwAK1MX1qSbDueHOwUoO3iVAKoCcOGrSamT5WVgpAbwtOdq9HhzRGxB7yYM5vA4G8TaGiSoGl
c3PVbQyf9XIOhMEHjj3h4wORscLoaOtS53f/9NMrrd5SSVuo2lNgaw3gpJtUGPjc/14qTZQPYApg
KG/eQjfXJbLZboW8+l/HLXn8zxHCH9u0NYjP7+HRdh4lcm3jWw0WIyBp+Q+udsrV7kF3ybd1uSjZ
qTKC83x6M3p7gCySmR832fQ5LjV7Z5fMsB1mrkk2oCHu5HKSPK0Q5fVOtQ3/10ZN5G1oGovcAHYt
MNLfTUN3R5Y57KdpSr1u0Bs8BauiNNSE8QbefrfVnEbTtvtcxPBGosUflEW1pZnq4Ka4BQMzZn06
nfnK96/rAjSHKQvZo94+SLqYtaHcLs+S8kgxQMa2bkWUsBb/yED3A9qIZOPykVb0FvffhXu/BciU
gIHtQ03OMJNFNiu8+pgOHmmcXxqPIXDEu5RFd7TttyxfTf4tkXeviH2PZQVSugyP+gdvpe7Bk1mH
12MRUjIJgjHMsWvzrjEIZ+AV+92tpPS3/V4KM72i1JcRH7J+EY3vt8iqsnUZUamOiMQiyKPCXZJ3
LQXOE1DWusJAV+jhgO4PSIZe+oSpcqhxdcl8rU35TiZa93+bUDLabqyOmO7AEjJuu+gHehIbAzq5
ILPUlA7frJCuZehQ5YOWGrGCRm0BFJgB4r02GXEeCg7y/SP410+Q8HjIscm7Y8FzxELFIsZ+c+zH
j4WzTJajxoSeZs66oBQaZedwCDjvyxbluAFdkxdslDj6qpyCfjvujKHWAp+kb9xnyHQ56wUhzKcu
7e40Lr2tPmQTjp3BojqGlKPeuPqGhvEjabKdjvqI8mItAD3sjkPLvmgxuSzWt9/qZt3MCuoMq1Ni
Ahqz+nbxMkfuhXbgPA7NB2nxYUrtpHWU9b3KmR4R/9HvApHkDYSQKrSmhL3Sdz46/i/0mAhMBmnY
J6p6UNQYxQR6IBXdZG11o5qdT8QB2MppI/gfpTLuR9cU8PUl+HubfSXF4b1ZhuvNl8llkavXYIcz
eDODxJO90tnpJ+iPGls6Q3x+wKBoUUuSajTqxXa7614BRDR/0zSbM9mwhINXfvZpDw7IWdaadVkn
Hyanm6XX/CvUsGmYy0Exx5RMDu6Bf3siaThV87OgzyQa3zOcvbNqNYvqCoj/B/O5Wg7pzbjq1AQ1
OLSoTpFeJIKq2H2ggwPalzPfgeSugWFzdRobHSe8xeOqh8BF02MsjzkrAYkjmb4Til7MoMF2YR4K
7MPumS2D9JPlBOhdNlCLir3Q/64wg8FBjkp0ypbuQznCgfHOwkh439co1BjUSU+rWzxnYJBpcEBB
kEqeIuVLQz/QKpAkXxlsBgOdkGZWYe4euwRXGrC1STldj3SFg/1wu8bHX5G8if7QDC29AoZJ5JmS
foAY9/tvPpLoENA6uuxfDrqE2gi/yew+e/fH0WITMYucbObrV1HiNvg9+p2SOXC5fAt7hNXtP2dW
qAIrQKOUHMfK/LkEyXx+Fx4fP1f3SlgZcVRBPBWoiNNTenUl3RuBq/o4rW19V07WpK7YwB1SanEK
sNBv09JZz57FQf7ZTSTGEouis3jXzEZdbH80o0dy5iw5noWmPmTu556A3TERBPEuKyBj8FS/cs0S
06/mLiRNzVrcsAObTSOfxqaH2L6e+WGkj5MZ5zeO/jHn8iGb4wnEDXms5lTDkAtTJOWQq+pm/dE2
ZFEMao+I6GEmu6bxf2jU9Ulcx2ffHGicez5iQO6Jai3Bg/vhYdjnSgMtQ47SeWZQxI8x7fENkowe
cZXd1fymeoSXvAGTxp4KobHA54C5/mpwYu9LmBcG/tE7bmfZG0MGH6OUOTVw8KdLuKKAL7wpWHSz
uPU/jO/s1arnIPMj6V45yhrKm09b7EziMx4PuhL69ptSvupvCDHf6jRh2uHUBpDMbzbWyy5oRfFU
JL2RjfO+adlxSnqJBG7/B+zjlMXfZIdl27mDQqwK/YwtWKCk1I+c/HEiNopbI6AXvqHiaKtlwFR5
NL5nZDomQ/8ajDCAp0hKFnfU9beRaQr7oU3W8JqcXStmYqFbDEpvLYajizK/+OTY3nkX3SmrtnQg
YSbBlW2Oi3XH2guCSSe78xp0xsSCI1UxS/yDSGNRCQn5jQxsxLzwjoORcM+Bs7c7XuXO/gWghUpe
ymoQhv1svbuCwMzsdyz5MmmO/3y9Mt70kpm0Bwu95guHb0E/mg5i3RYrOc0E4oQpvvAeuEKVPKO2
M9Bdyloq+DQHqm9b6+dnrBz4+qAzzKeH+Lk412P7FSTNxqJAyM55BXznGC0OiJUyXZU8WDXVVlJI
xAwlNDTH0KFo0fgf/diKag5c+e9axXZHNOBu5IiTh4Sp+U+9hd9guRPhf0jYCJvB1FpYf7/GI+oM
+HEj2JFN+E6+9fG5C1nuVBKcltn0RcPfASIk86905qfvZtXQxslaKZzZY1iCC3+qgFTIdBD7LJMZ
TFci1lxqKIDJPCFpS1rzqS82rUqzrylrVhiGcg2/IO8pD7d6Z5UceVO9ISEUjR51QVmvrPTrkac1
xbUkrz2NTjuAO32L9M9Rr+b//x4pDeTUQa3zYcSQXd2tpx9qllZ/tJe2/BPSdZ6XamytLuIT0DYr
GPp0izmFh1palKtglFYyRghfG8nSwkczpcSJYVZCme2imV3YQksehqhIvZxBkk8qhqvbTaDXlNYk
bIiwObQuADfD151Ir4PRb35JuIAQ9oyORd4X4uDZzvnXWCp9PlQ1ORMNhboUilzmjQ/eZp5sL1Aa
yPrWsGvflQe9GQmOH5vY5R5W0jbjC+MAu4WMZbLPVjs3UssJzh2SZx++WFhABeSN2bxntW34jxfm
RuaZjnagjbNgK0CeuLcO7umQTuLsAja4aBxEacnaoVXH++Yh3WK8M6TQhwa8C/CZn+ts3nxHUmMu
MdH4fG2g7PDOayChzx7rgk86TRvxWC40q1F7ZFi9R3HxcZb9ntBwa2js97oDPAMx33MPYGpxCWts
jkPSdhoV9aRsZc+dwdNugBWiYMFBDU1VC0CyNIkdIUrRr38Q5XvrMHTnKh18TKDM2CesKe3ZYtIW
tRHRoZTPYkxeYInh8/RzAwLj6SoK2KBGno+9zwdSZwxnMdq9bVgy1Ucu+cT0MQ6tWibPFh0ugrix
GAGudsFAQIQ5ESySgq4JO+nkP0LYbv4HQGqeTv4zoFOLUixzbpXKFeBKYhAUAiwVqXsZMM8ddgis
/mxxSbu7HNVYfEidm0mWn02wHWYye8h+yRqmEnrTctHvjHHcFE6xTUPqX11K6S+Gc3HvetkvJO5t
MEz7GMpAicMafG+rr2CP0td57wi5C08a0ZvrZe5qjGd9dfHXbyIWnqFHaYkOQouv0deQ/aYh8Yv9
z5EXENLuZHU0X6GmIya6ln2eKUDN6hy/IIHOlxHn07apM1ePu/cYGvqIYlSAhsn50cwIx1/ePHAA
M3BtKdsSAbBsOlw5P/bH++B2vd8Cm5G/pCT5jsiI5rAZJ4RWtyTE2CHVDoiYRm0YJTVXzUAheU/R
dmZS7w4pG1nRWQHnuQnC0J1zHWC+k9WxN/nqfbDiTG1cvqcj69V6xa/Am3bVgC/ewquz1YV1a+Z3
Nnn3xYhHBzlZ4ag70of0Iq9dBdV7CZUpPyp/IY6WW/Q0CK010AqfIdh/e3RYdtN5/TvtiA3paPIG
l2QXbBtRa5SUN8PocqM5V95UZ2AHpd87lRxftjVGMNu0l+Q1ePLAUFGCFIshYNAOsAkXkAs8HkWa
7mRehVGsIfpQojrYGotpZqj4A6qCnpdXuujiX5SljUWb/QRNeEMy8loSdsok4fVFjR3pFcee05me
Fhw+E/deEcmo9f28bMmrUMq3zZghwvz+oIixRU2KgJ7C1d9r71X0SBCSDbZP7Ga2wYzYttP+UGZ4
NdQCLxxFPnLjmBfUklQ/eu9IVV5gYQte6QGuQyeK+QQQMMLk4cWRI9jT16XvXUZxisoJKTgXpAOr
QZgAfTj6W8/BEma5hlQ1XZEGh7YJJtp9nKdZtEAs7elM7uBSO0HuJH7gealvgmWvw8rHUmY2eEWs
y71DXkHHmatFNfRhHVvM6NH/AJrVxudkgUH4gMo6ZktrZCiEky0FULsxlttdGczcQgmtpDY9Oz4b
OyZZ+1Cx0KphT5QDrqxBve+xObDLAqMpeKzfQgBwxsrOmNia1VzaL1RsKVhg2XmwcmNsYQD7ItJb
4GukTJxfl0/vwLNgPP+s0B4DV6ArNI8b/B3p9Tpzgp17crIL9p319dr7CkP/JUxHBheGZIzFJ7da
xYRNt4o6eZXOsjR4c0lYbKAsKDD0YTdyD52Ysy3pwwPxtLIyg/KiZ8ebGOpJQOXuvP0ofAKp7wxJ
wtaXV7xAvunzlQ6f1K7gsqvQih7UwjsrtU7CnDyHaDmSHNtjW2V0IvrkuwstCDQo4QbfNVhTCBC4
ZdqR6FJGdj/KdKGHfmIBFxgHJqtvV2mhTY4CgdCt/fIEvdceuXr131CZfdUAi3WHxtYHxUPzygQK
R+rnIKkpvA3N0icOBX1osk6qRi5txpxfzoeQtmstbxpj8UhArzAFpomIcOPaf4gWdNvUc+tOSBxw
b4AgDdtgXYO2naQ8uL7aidJTJ30H34ItWXktTKOchjk7moFXDQCWKuoyI7IsnuMOmY4Gw6h7q62j
P3kRjXRMyf1pofFUIhh+1oGV2UWo2QlsI1dfadyIFxNhnhEO6161ZXz/mOucbC8BrSugggx++Etf
rxewGbbO03XenliA3zGi94mI6yFghPmjZvd0Ky+NXN7m4nvjlUfh1hwD/tskVcJpKD+H82qVxjfw
SKyS++3o42BbrpxnGC2nuSNCEcpuMOr8QAWnsmxRp0ss8zpiEW4tJ8b1/ip27OwWNPKs5t7kDP0P
KoeJSFKOc5L5MZ23PWpdZ7w3sbNZIOf0PnVqCDDgmC2+BZVfRKPemvqnqPtqh9F+o14cxUgMT9sv
8vRNVutDKZNpAI9Kyn7mXLkMt0GY3FQqYqB4/sfdzaByanVlB+lyjL51eOiPAXu3HiUJCmBzfXYT
iDU8BRbsnY2gfMOQ8csL2BKY1Nm+GQmr6BYH/yGAglSzuxmPaOypvaZF9xyhpI9fhiYawpBH72S3
Nu5RyCnW7mPS7VZtGozWHyb6rs4afvmzVUUPlWzh4PaQWG0tpkbD09HH+7fcszeXEjM4VwL13Gd8
e1cuEjfmHxTtHiWzQI1enY//2bwr4LxNg72NCNZQNlsQWLli9d6Bnl9wl+1J4yhvEx1MZGyDPAPh
49+QGA5lCtPnVhZ1EZYjppH8Il4tMZ1Q5+y23Weomx+OxN3dDXUqPjyW3NKWNztpUC3I5+afDnT1
sPZ7fFXZ5EKutgBWQJrj0jokIRY61DgOTSeMnkZvu8AiWx2HmPIE/K1xdheVi7t31sjLHJ/bV7PU
300JzdyjfpcVgMX6wjIckDZ2PbMgBq4chZrSmDkMvGxyemLLBlQdVrxblxqncfjytEkLWz4sDFWc
SfClc9pFXldy46M8ZpxS93QcsUSB+jl8YOS9a19d9EecVzkG+V01q0EVmH3dTI7YUr6VWa9TxGuk
5sxj74DZTDrWP3JWFStP2zJw4FseNhGcpOorrM5Ikk7gYRvBzaCobJqDZnW4USjO/fJhzmIshzI/
SCBTbtna/O+S9qsWw1WxnYv2uRlKoDKwLMXWW+WrPqRYmbye7/VyDQaQKiu4SIRHceQGkv2d/7Th
upb6kOjL4GYo5548TusV8Q0WFUvS9M5YQb09KTiStXwKU1KRxUuoTiEHwVxAj5jgypeLJl1rM5ke
SAj+CUDckI92IyUKukdrrnWXUDr+tWz2XJdPdJj2BgzPzGjyOJ3HlgeqRN76lKJIgpJOjGgmVXu/
3hXfG8MPBL+ecJvPVbj6bFW5Oo+d3d//mfhZqT3Bc68mswBvhCCaB0woqNaOLeOE1ohIA9crlqBY
VTgNETuBcmmgIxKfaVA8bW6pQnsnGaIpHD4nhq96vdSeg4Uda8ZRjOFRmGW6/4FH4klPwTw0v01N
AEitmrDgZ7IJiP4kCMFU2UQwApa/n3dIJoUIY98haIa3UWJbv8oLPlm+6Qeiq+9hpCnN9jdik0Pq
1uhb8bc9f2xagTY2CRhub2exfaog2NLbBV7MtOqQ7tImOfxQtQPlu2o97iqzR2RgS/rvBvYkMnW4
XnaHWghX0TchheePUYx4lIzL3xxFsITh/G0YnGT3xNSg2Vr+blsvS7Dt1fqe50W4x11JkCQBQynZ
sL+gLysQkJyNO9wTqarrUkjyJKDamLqrJN+0z79o6wD1FbuglyRZouZbDAw2y1810LGL04pK1esv
xnDbJqQBaN1jP6xjPMr1NYdcfKOnYf2gtjwsxWDjAP4krJNTkgPZVlG6wkcZp2XcHsvFYGaMlkU2
fTtvpbxXYYSeXR277CdiyuA7EiEzY9Fr8h+Ze/WUN9BG5hkLXNHjSR0e3XncD7PzCQr+Lz/+2idQ
vfYA7Qc+grY7vKvAMMuj1wdJtmpGq9NoVp4TE57VZG0IpA/T6FWw0bsC7eukh9JkjvFef4te81II
JtSA2g2tkiVJe5byf7bbVjBO5TS5PbqhOmRuY221ZBlLq6oGPqUGq7DWtp601y/pf6W+NUT8QP1i
EpMZZ81wPtgcE0pyrX1j2Gp+/eVSVKjxJj55wIxASUwE4aDXTj2HK8L1nonF1eIYvXzCQCmsMdkc
Is4V1yljseKnBqRUd7gDwp3jEAuZ/v17eVrNTjGbZs7HH+LDsuovSgzDN0LkzmLkXBWAEoc1IVKY
Z0PEoteqtEaTV4Q35i5w4KsgQI3yols3U5rsZAhx2oB2XW2vc1jtzPb9lo9os8SiSDPtp3wSaJfG
YwW/dOoSktWEK3ihVHPBdaMUltnjxH55TGRv/bcFllNuznUmWrYuYSeCo04nNcCoD/eHeiAn6voq
8bDkM4DrU0zMndR+G9fg9yy3EeQaGz/f395FNIZvvJtzsB5B8Q+gx3LvIynVEkf/2AfiC/ilz4em
IgpazOGNqwfj6cfO4L7jtcTLOJX8klnE2gj8MS1VG66hmDnbALEYv9DVuwDfBm/OqNubRI22QRvj
9dXWq6oB5M5t3sJvQOn5rqMNYEkKLKQmThy5zzzk+4iuWceXVzVTqEM+IzCMIkVyVGzNSI1t1oFO
Gau9wqIFrRXMyEAjzNHezwwqwL02LvnxXEK6VsPD5ptKW33KIOZl3UGqdGnzbRl4sejmZ6re9ljZ
x8tRw2bn4sHi7HE/P0iWk0fNBoySRIOttmaydPoIcde2TKiFfI+dRjp1FlLNTDjgM734iMcKFOmD
jxP8Qv5J5Uw1zDtkxwIRyXGpUN8dIVIRFYmwS29CxtzHMfFjvFrLOS9beriS3r/vjVD8dhqrvCMT
0APSvK17jmB8Z1sKvFmW56tCfa/g4KQwBLsO6xjzAstW4YTWlbpodkjTXu40u3RjfPoGfUsWOw03
QDoKxMB1GmvlNJZwiPfAvzf8Iyr8H7M+9voPbDRFJqcQVFB3DGGzVQCAgsYjPg3/IcIVVo0L2XT5
vOC+pkJ9AwXKThYA4Mcrz27l2QknfIqEFoaVBA2YqkjsrrIX+NEaItKRv51HlH51C5RDmcaWSgz7
hyZ+RqKs46nzcLiDS7VkPdzR90O8qYe87x5zuLTJWAG/EdUbknZUUFLFpNYyYA/2Y7X8FgRS9sIJ
ygxyrsKeMBVfaNsPy336jqcdYRa0vMTHzpk2l3GD4+VYFmuyAnEDiAosteivrBqZYiiUNPEqOHRV
ljThUZRcOQhRRyY5dA4DR/UhtvR1zPWBYSOzw9r9bh/OKdQjSHMouFPRghJaDAoFZZryk4N9qgfC
qh+nzFjVxFPp2Q1pA8t+hXKGqe6jcoZVba1JGh6R9qrXxp/JaOpXIsneuk6C7hu3KVxqjOu1fWKA
0d8jRwWVTdrhG3UyGGaD7qG6QniOr3luXGbpAlPhMElQfjdYZY5+1FZlbpDNZHKCvnE+zI2WvsTE
70TKKBytTpnJlZG57TK19Z42x8dMaL8g5yRayZL+rqxlpcP1Sqqq1pQ9B2YlrxgLpXV53eput0xz
XCyEy0zigLLGTFAfxE8Cz5olrSzw6UFz5LuLTo6PuM8sXFOWVoa+s5tgXPbt9mmiWmPgFcoM9TNF
pILoe0vz3Uww3Jg3WovAW03CzfCEsdgF8YXgWHWuN+kWTbRZMo74VygOylmBulwdqv2U1wzvY0a1
cbFTzLRkUYNg16wJ+tlP71GbEeqcYhLRF0sHdXe4zn5XAy/IOya5GUa6+0OU6rub6s76u9gxfDg/
Uk2mUWmHwfvJcoSpHdF3EHil3o97lpFByf6x2wcjhVVnEKTBnIK3OUSK8JLn1KKV+VFupMMyp05c
AMSuFsiT9k/SlykEk/N/V76WBGNaSLpBke+icoRU6VOOe2HESEuk2veEM5rkXi9zUSuYBJ6tcOo5
BPlb3xsaCQjBLqGP6RMWM6xey3sKSg70YQoTuKNnQMMfXe5y1/K2GgdQ4uAgUnpGof+rr2OvwpCA
Y/C+Zso0dNPE8XCYzBMp6uafOv2xIG1bTeI0g4QpYzpWnQunAxHb3Ns1zfAmskWUQvKWDPR5CmOb
sIa+DCEV+CHvLd88RlzKu2F7pG4t8xMzKkAJXOO3OLlv2ywdnMn7GMFGJxdhGgCNaJvcECq77ivP
3XkFLOQJPj0g/jX7ZQorQPpyiFmycRW7Wb1yg73/MZu7OXhDLdIFsoK1dDL6QGiUVJrl6G1CJT0o
JkqE4Zt63J9St7HjYPjTKoEd14xOW5bdbiWZd/yduaIs85nUAxMv5Utrmqckq1aafLJ+KkwZgeHK
KcG2K0MEsy5904ILhyX3WPHALh3WUUo2p+5A7oXbw9ZujX+4UTJSkwQN25zFR7uy4aPVZkClPEg5
UHED3Z9rbbtoAgLDcOljE1zFFFYzwWhue86zMQ1IW2LO9HPhvBK5P2ueMdSnxLh+qZbkleTAvhuC
pHFT9D2PdE+jFVJTEu+E+6VWfRUvKXbLQ+S/H5mNCd5t7IDh6eLr/wkxi/VYnFjvY61aPz9GC6DA
9fl/4Yz0quLrRofNDFYj1xDLtREtWK4vcg1tL9NYatyAV8Gi853Am/YrzbyrcQMzDckVG6fO9ukV
k+ue+8FGpGz0hpSkIGdPA6p6XF0N/QW8c2573MGeWKHjHxLoinq7G+XqLQlP9vjY0MldP1pZiI6D
HymBWovt4hlk1Gauo6IA1TAgi1YCL2Lo7zrLLMuY7eNm1J8HbkDu31zY+vlQPpvftNuIsrjBjbx/
5R1U2L6kbebhucopBF2YlVOHY8MnONPllJ1gG5qGVhp5lx2zj0sGA3u4wtytJw/7kjjyagqvKkkS
ZJ7KGK4UJPICQ2FzB3CqopBiILJi79ToAE2ybiPkSkHXUPOSEPucjYy8x10HuCrDJzWELBRqBu2o
v7m6Pw/Whwd6AvKzSntYK+qOD9IMwutvCAuwfiO4fnNX4r7Di6rx8PRfQOjzCWEsaaHweH3ZrU8b
SRmwTMSeVzOPl91cobSdoiMewoxdD6RLKqEy1ZVI7Xdx/toLL910KpnZHGh+G4/OThkH9Py4lk0j
leBflJhnIADIm3n3nFr9H/GqcwGj2C6HqwGpGmRfYa/GifZ1NuOrOYitWIFHiz6UeP/bTWU0GLpS
n7Dr3DP+1VjetdGThlwaC5Sr6w8ROuDk+eGRtYP7VsbCBMGUWRFkJ111sNsMaKm0EMKQf4E+IehW
OiKXkAysKBn1BLr0gYOt6heH91XMyqzyO8kyEKzXuy5JnMfcvIbJx5qSSODGFzwnJo3TnHCvjGnn
5o5rHJ+EninL8KjVRm/pjBLGLrquDxAa+Ng3OGMmN87T0WOVLODnKQIjfgKeF2cVO6QcKlKp9o9A
i1S+urL1Dspyj/FRvjuQim/FdsRlIGHnP8xb3Bv1XPwjeEIC2UA+M9HOhmuQz/VEzhSU2z9qlwRZ
zW7GfdX9uMVSGBsB+jLHBGTJVY8MoqJD+dlG5xnhlAFxza4oTqDvD4pguOXUABxFAz+zmWqzqnOs
scZKaq2aQ3De9Yioef5qX+qFvsVEk9O6coRjw4VIjVQlhL8klJJTiL4MyPTurmJSd6wcz71rw+ia
jtb0w/4xzllbvjKKu49yBlbj1pxKayt8fEQahx/VxKxfH3MELNxzcTidobrFMeur0UfseeKoVYd7
ClOsuqFFG5m7VZM3p+fMXQIiADIh9gd8ejgYdyzyEnvU3oCgKgwsh9lbE7oczAABI6ddomcf8D8V
hse9UVaZiB0C4XqWOzlTaXSTs8dCQonUfXw4FrvhBWjkXUi0TC9pnLVoPJ5u/meTxjuHuLYxWGT1
WM3uY+oDJpRd6zrywdm4J+wo2WxXyXYRjH4FjqHNEfRx59zs+HMNY5u1RChECRi9IiPq0Os5uDD8
CUBHDRflrufYr1rDGunORISnNslMJnqQs/jytkWqvQoiIR3IjfE16Ccta2TGbetxXEVx2OC6g+su
w2sH1l2+s/yUBc3nMMvCbcNpofnC9SSE92aqA6VCm1a/ZBEz95zGiD4FpcFuSZfSg9NyS4Xl0OLM
xlIOK1yZxflMucCWUbQDiGcAs+dc6nDLS6FdW+7Wc8v59Pn3SqHzclJAqd8X2MCBh8OEM3Jx+vFk
FIkXX6dGDz9bHI8o4AAKSY3PYqNVUlai93pg7q/pXZfalYh3pIY9bGvHrhhUYy/MrgnQXyV1kBEO
qzEB5CuXqmH65nlZHt0FfNf0tHn9Zqd4mOaX91Skd/Un44JPyJYR3JGMm/n9mgaT3DyjtAOBQzIp
kQza7J1UtQgtN1q32wlT3EeaecXTX/P6W16rLfrHZHh/oRQUVyq/viGGo/B8YEC/DiAHIE5n+KYa
43PjgYMhBhPdDrEmr5KnsQ1GURKQxpqzbsbnUC6M4684g45ituJCeb+zybyI0kzUpMCjeIofLdHY
Xs8kBkBRzmJ9tG8ZV6xcUu6mCCmGYbaYWOsJ9eTPc8y3uz1VurpKTE0olcocisVOFSdQpF5ym1nI
Un+8cNQH9Yofcf+Te1eMFthAVDcqXWQ7TijY8raPNp5WqFhfNq53pTBhVVcXW+oRFrXy/2mYjK2Y
y0nn+K/o4Tkd8kCJK84dP7JQv79sLJStZAi859+bnSHVNlJqlvGTNr0qMq2enR3SIi1Ned31P5pn
bHlEBJJ0h3qQRI20E+mbWIbjPG2IVBJcGLoA4utgIASNwrfuVAzeXWFJRuGfw1LyP/DkAvlDyBsI
Xvz8h9kJd5YpkZlnuFvqO0dXrpMhZlRlBI3O6EkyYhwLmXxBCFI50gz7J56QyGEM45+LvG+yz1Tg
HJl53VZwLhL0qidBaGuPe3U0fbbdDb5eF47Vvg24QPCKlrNjBF/2kNeIZ0ZPzQ6ymxWzfHmWMtw2
1p3SghAIqjobbUeD/GJosd70K9Df7HdhOwAFhrfQghI3gjI/a5SBva7qI6q9ffW7njiatXdL5pzi
5afm841knV4rsLcoCVRqN0v3FF1kk/mEzT3hp0KxZBEcYugADzedOgTXkf7wnL22smfHdOjE6qqN
7BM6Gcg7slIir7a4hJOiXLWA2PqYgBQ37493nWCZ8H7U2XPtIv7JTEWxXDhi+P5u7mKxQZQqrrLW
gbfAe5hU9k05VH26EfIBGZHCy2pOUtUAMuaNgjateQ2pY94y07j7lpTh2sg0Hq2mGSawUv8nc3Xn
w+e2JKG9MRkzkDqIXzuPcKA5xeg0KsQabYJMQ1J5z4MvVxzNI/cL4pGsZXNgJe24Pa5e3iULlAch
wAd7mxup3XbBoP1deUH310OombAqVK+pYmUPWf8JTaPmuvYn5PQjP1HVFgqBQs6zDwUoLigzt45M
uUxedymKlzHGsSyBUYgexcnq5ug/MrKN+QUllH+tLfWQWetxSE1GJDGgmxED85pHF/6xwOyNTO91
fuxDxF7XbDt7tD4Z9GoqxZvj6RalarxJs/5UqtwPLhEheKHk1zlTSK6Uewv684vhcda/j8GebGyt
1NCsZBvwA2TvNK8XMBnzJLcxyhpi8g+NtsnE9Jp1w2o7REg9KYGREi5LJT1FIeqvOQhwdyN4DsK5
OPguexFp1rwip6tV3GWPNUCvEp9E3WR8igfRBOAN2Z2j0VZaAg4MwryzRW48ykApKKNjU2wv7zOG
Nt8CmXegTEwFZgs6EGA8GIyqmPH2ACIM2cXsN0CTVjjElr80K6o8ucaNl89HgMMd/2E/tWUFjPx/
x8Q+25aPXclz9NwLtNuC7s9V4pxL0pd5Kl/lGnFyAMWVRXiKiiUBjbYfK1+N97sIy651fiNwEYs9
d472JF5nK3j5WngrWU/2Jsci6NDCBbsI4L48UH8CokbBcunm8z8agVSXLqyw/mYPg6I+WVWAA68A
ijgZhq2sfXlV1hWuUVYnFhX/TUSS03OAcaxT3H5merqyVAS9qikwK4C5u5XmxhxVZfg+5tCCiSE4
YaTSEgs4Cn4eIl1zCZvB2moA9ubWJ3/ovWmdax4wSAIcL92iM50dLneM6K8s70Qv+UJE5F45eqn8
8FJOvHzhJ3cGttN4Mj6lcoFKwm97CpmZvRfqQDbqz4EK3syHSneLHVD78o611cpYhJZHrAAMNE4T
OQR13DNZkCTs+rtlztGdY/nm+WJ26995b9AAFbVweM2gSfuYHJBIEIoKJ+PXWQSborK62Tpzpm/+
z/RAAvMSeNF1rZNW4GzG3tZpAWBbi/lUzEk8XNgfSjt6Z67+UBNkIefZQ+cvY8uCUgxjpTLGoOg2
b4SCcush5mXe2ORJ58L2I4hI21kRm+yAZMnZS+H2Rm9PB1MdFnCxqWzgeoeecGqvERPNnb+jUpEo
O9rJ3sDELBfElVoFTBB599Sug7w+IEZuiWi2It89FzjtDL2SCzrKV2UDW38739/AVF/h/rtYQwgN
HJnX6oc2QXiyMxlZdXXjoPTF37DK1bKP2eDN5EtdSmvjgSUZbMU3k+D6/9/jUZeRrN9si+bODZZa
7w+HE9u135N0pQGr1FU2qhoqleP25LUVMV6AA3dLN7V8bsjIpfB2Z+Rw66XVtufA20fjVLTd0gAI
Al9OZJJrS/wmv+qdScRezQ4wvD1M4xcgApW/bRwhkPZRrydTgzqqJpc/CTrVwQcGgVTyveTlYxOh
jnRQhTCC9NY8dKOS6jIKlUkNaGuSFlu7SU1LanHu0HIl3lvNpOoz7ou8sLzdtMWgRtQ7wUXDU7cc
sOeoF7MT+Bw44zgTF7zr5y+wb/3hVbNoW/vl5maMMtwUMbLaTZ0LvyO/z0J6I7N8S3FdYnXd76B5
bQjCOS7szNUWNj1/zXlfy2CqcGLz4H227+U3G78/59qQbeiPiMy/hd9jR2+aUtRyMathWVeS+0SQ
Qej5J46Zr8PGBij4k3icLViofUfQSTh5uCTn2+koelhuB+Zvr765Gj694xMb1XY1/r0T+oatvIUc
KngUiKcMyO6ovsupJwT5SbwFX5XVAI9VoA+sfZmgpvKPKrl2V9b8pR/Hdh9PFtJDMDFV7pvSbZan
Sn7kMxmP057sjHvnA0eSF87ITAoYVZ3RROyAsrk59+rsbjpSathl5H1yGu5AmtylS4sm5MXTLmzx
xjcyhhfXf8sclYIDYae6xQffkaW7v1EtGDDlVgDfQTtGgpYH7fNvoZp8M/OG8R4NdOUVifOdFBB8
0YZqzSL71WLR+xEZt19M3kpREVxffNXUiIydK6DRdTmYTo+DF0BcwZo132PPuHhAk+cr6dCpfIoJ
+GfZd1jjGmSH9IeALPwIYvAc3sHe1HOxpfuUaP7LyML4AOt+FlPit4PowPY04s3SkRtI2+fIF3CI
MGiDDGxqKR0HwgU4wQ0uY+cSn6chNtWrEkDcM5AOcb2dLHdbsgAaeJ6KeuJeHEwJl1xV3H2EvN6Y
Li9wJvMt+mVDGodhmBPqUTz8/ug1EYNB/DJOf5Jkwn0wFgxxd74LhoscpLjm8VxydlG8rsoTgHh4
qkzs58JazWRqNxyvDWp2zO6WBx8kzq+QCIoLayYnvSB9g34X5kYRoNfS6J6sjTWV+tSUXWrBUdMy
8BNVlx1hmrNDcAqWu/5YXFXgYORSVGs0LlFyjczhFDi5drRu7mCQpuXpE+gdu8ttNvJsMMr2eiRS
p5xnUIDgiI5Cjtf0akw6ZZ29Wp6SbO+fIFWJgNHvSQuYv1l2U74StDtADoTi5ebmIpYhdnGqXJlK
zLXE4iwkRZ0Uh12O4+SFQGFYRHQW77fbRyjaRKkuRkdT4uRMfG7J7F24ed2p5+fk7qembssYZVcP
63HbKDru7dAh78fAI/9Ljwcs2SSv2Dh498X3v92VOxKn/jiHFUcAPSGbGiUQz4UZ31Pf3gjprC3r
IqMuugL4I5iA8RJ4LE0C+ivMmAwsed+PtEmRA4ZTp2PHqMi38NA1L9TVDkpaWwht8R2xE7KHjYYK
QqtPLtx5GlDhu2QjhDT/ZgzW+rL6PHHO0Ex2OvvVsYTNEbzOXc8NreyOV/ts2QA5pbTQDPYUlEMA
e675QrDWlsMGKFgzYh/DSzFuz9GEB1BqrB+yAKUjXlU0SKZ8hZgcEvxtWljx0flEYaKfmd0D8A+C
IdcxhTUrkDPV1fa4TYptT33xDlNIlz7vX5gkA+mb3WSKS709D8QqRs7RgN1WOl441e/gryxVgbBA
ceCM3LuhrDuIp9dmXyZq2SBEQ/hBZTYSiK6NjH04AS8U2USdALoQ7109HtnvODiiLZwvu1j1WqD9
eSBD2fmJ1rYAQwwlGa3qqixbN++NxrKoAUsDuKB9yW03KI8Rt/c6nOiGOBU7yr3Xm4Q3wgIWm/4d
EcBIPJiP3lFf+nkJTLXzdFSpsZZ0kQQSxJ48A3PchP+kPtX5PjAfhsCNDZEy7EIFFfXGZkvx6tFe
H6TvIeiAFjoLwaffWTWCPh2rzXv/9gFlkbx5UMtUDrEb5wwbRjRh4ru5ScywwI0dBoVLGvGBa+Mc
/UbT0ciGkGCVn5+3PuoypSLra4IrmYwq8Der56T+3VWGbd5rC2uUFcV1Xe4ZeiSMmvPHYEfBGHnN
PHJ/fpyn2LSHJ1Zjdspe8XgmOfmG7Ap3odf9R9DpKOyCkK+lwDyT8+rMiRFI9YviQCPAEU+PY9Nc
mvhKVWxwyJlPXCExujqJrVHO8Xm/cLH+1tbe9TNonpru6AgB302WMbWtjQq4O5orhHlp4+6R4Y26
VOqwfBTWEGnXXH+PH4OlZgCo4u/2zZqHUas7TinsFg28Aqfoz7TdnsK+bfKcnQWodhL6lf/15fSN
rpdb4sX+4jgmhysYk8msUvoTD0+cPR1gEh5yvGfz0ZNuj5EkN/sZ6GxmTkNLfu3aiZoNk2lYci3h
DiDK3m1eAbktFfROoCT8bC2bvBIHPR4E7DyOOKovrmYcGcPIQ2zNUritVe2AzRfIR6q/7qfRkzY5
HTJW8bmH0nmKDr7c7F/BqyWTJY6ci4q1zDKhmhIop5IZgcomjJzqtmsm7rPU1bDxXqOKyo4RVu/Q
eNdXyrs6Y3vPUmp9uMMSG03C+4ketb7z6phsXA1OlJiB/i1hM9Dv4sVmIp6Hykr+5xH0nxhm55PI
DcnVKUiY9xwMWmw3JELAPXxrvgzXTtJDFFysFF4NTb/32FNFvuzSmhUWItGdD6lSkQ+wecJ/N7GX
ZICLCxpt9mOk5Yxpur74wDoS4fnzvTmnNe/on/+LFimtNBAU4WjMJyBhZXQn9GqXgsRr/v0l62Al
9cp20C3hBTOs+x78DtKMXxVStvMAk5Vdr5LOV5lzkHKpUehNrRQZ1UMFEWeSaZgLShMua7sSAbHS
ZrCl38NPYoEektCE4a6u1aZRz4HS6nUVpZmLKi1TYqh1+LZy1HDrVruUtXnMNFh3dt1Xkxo77cvo
gqiGtTW9KT4ej0J5t8ot9D3OkEbyP3MGC/L+7jEWJn+vEcOHJSoB7wsKHFxpvEEWkgUqbIzGAMQP
9U8+rBwKf4xSIq912Y95AFRjqqTM64L4Vm8WHluvyViT4qjdf8ZLA6zOBz4RyLZZR8GhN6EePXR+
oiBfvpqdyAatj0YZ8UabnL5R3OJSgxP635in5IHJF9+ycaKIo0NmJYOQZCEYtHcynR03YRySSs26
sE5lG1lzYCt2vqHmYl4E/0qCxdIV1Prp2AeQIkmuQ0gyvkZecn9gzvHNcNw2rMa2F86/vJYJbkWf
y+jMUka+3IObADKFUCupwmk9gKxRbDb2ommxv0WrcRj4DEqA8CIeAmaywdk9Fhu1s/pgEdxjOE44
K7HtiKDHMgPLNFpEP3iBj0dK8t2MT8qx+EDi4O5aQL0CgvxX1yNxobCpgZcM9KAeDPd4Np/PA4m4
+I5nWKRZGm5pbtKBbSpXVZuY/SibDwlFpAWSsTbEBCcNNendvFXbl0NjlExD08eJPMCWAo8EmLQq
jHW+SN/lt4KfX7q5P+PXzlIW5VvMl6MCTds97zQ9BzqYUrLeDlIRjQLZt2/B2canku38/15qeWH9
RFTo1lQz0KDGsQ27Wp2Jb8H7C68mKcWC7QkFtNdTjS5VVEwNNau1hXU3L/hwRhv35jwBdC7tluR4
F4Bf9w9Epqnqk+28UPBOq9VOLBp0yK5RQeFj8KfEPw0COfebCheqvAbYAt/h/0I3uADGsqzSvF63
jKxKRgz06B8fEwku7p8f7FLq6uTsiEX3MGCNNgBJlm/AA6ErvuAQaKCROutDEf8dqg3REurGjIuJ
ZiOP7HIfEM6PJ7tUEU6cKzE6usTqrfMiDUTRiRMTZbzVJYNnPmY0OCGBCzm7VS7b4Wo2+FYxjBq6
3BrwJTvD4+QXSM0wdLhvJf+G2OSpGuWAuowVZe+lvP5N6TaGBfJmXA//1XWrG8b8qhncpHlPaopF
coxuDeki/EoxzTRuZtpqDPClnqjVAWWb/NqVNVR5N0oG7ODTpyP/Mm+uvREl5C6usbdlSW+lz+ji
nibkHMEBJS8JuzwdePnLJsXLhl7+1kxUADi5UNA55cwTJUeRg2JSaI/W5Q6c2e60A58FMH8f0xQR
pNhomRPkFP6QGqceiQu/WOvkBz6e77fxvk5fu5Yy+PrLw5N51vwARNxJzqLcBC9LdncUDu4zlrgI
XOk6tFzKCKW2IbTxpxMdIvAyFEiJhWVIcPa+0ASdJip/RNS2ZrH2GICRzzsEh4fwQuyby7yHLImY
0DhBWW0B6aRR+Kk2UIR6ZQOjBQCSQDV1jNZKtaJ9jji7a9QHv+WhVxJ0t/UtZeZnXkF1M0HT9k18
6hENVzwqCRi7GumHHUqPOU0TY+Hsvx6200V70zw051fXoJqzljkQw51z4FTTYFJp00+JynRiRcMw
KyLY8cLTrSElPlRZ5bPUzOeyXgjBOURiTI9Hfsmld9kixLOwYb9Orw2yjGV8UykPPAQR4ChaXMVd
EhD92SDPNrcskxHd9L1RKPUZNCVaRHBjUYjsS7DV0GAWUOtx9t1OZNFySaDmPL4wTTnknL93q3EM
KNJUqCD7x8abj1aPTWCNVlMGoYtoUqP83gXOgalgtBz5EzM2yGRbK6kd8NSxqCF8h83yHScvVmL3
3weukUm5uueInPVQ5TTOW9W4SdJ4fPoewOOqZN8ynFlHVwoMC7/MIkU/rSwMAvNKTd/SV6X/6fcp
59IwoAw3XB7E0cPKetaq4jQvXrOhbuxo3O0SvuKDiML8w74lrGgUedyprA8gAOcWPMYE3DPxBdeJ
QrWvxEAWaBONmG3Hu1UDcuY0lY5uZC1X3M8g9QXme0MjrnQv6LW8rcmvdd2T72hI5Jx29f1oI3Y2
U2r/XKLOHbkccLWHE+tKBN55XbdgCKMqzUdR3b2sTY6+GjBVyTROi1D/1VvdAlr3LfGKnZdveOLJ
XTyaZsxxiydOA1uHg8uMo/yk3VZkTfMatpApdozWkhRcMMLUh3h06SRlZfoNsexlOXSqV57Mzzgk
UYXvLQIHn5zIEyU8hXqyANBqUS5qmBqlQRetP608Gc4jOwzyBtvUXU6flogW3ZjZXIFyPCLYBstA
aHK5F+2ktoQ9dRXMnLKFdaa1T04mKvh1nX3XWPOBgSFRDhWHhZDEsnDhqZ1Mm6bVJMzk8WQyYKVZ
rUgEyPC+AuAXfBxxmS189BEkYje0FRMjWcxHBTMxhFnABcovKRA1sj+uIkcSDEkU4lhWprdKgN4M
neS7ru7aWZbAi78+YYkP5WWf1H5Hk5a4VX4mY1H6CtUUu1nSl0LTk0UuSbwPwoZB41dm9XULmB8R
bdSiOnnAnwEFJE7Gvk2Ja5keZURkybuXq7aZwxAfO24BBFUzkQy5MP/X0WLwR/lsoS/KDBiY0EN7
9zQLaiBq1x+UWO1+kcI10dtkcM4OGkbLc0fKiMXjGKXF+eFnsqTbGkx5kENZtEr05e2dsjLPmedM
n+xJTeLGBnPE8hRBpK3fef2HYHa7iBuu/Ke2vdaq+UyNX6Am1/pDHzUj/q2HIiUmA99JRrfgnz4W
2J0VMcZ0NuNH4aCW5ARS/cBaJwviB0y1wwupnuhYtH6YCbz26PPBVPBmW6RLMQMTuu9AkK9x+0jw
T0Y91/or9/p0FF+yL2So3ufjQjNDMfHyXIBQB9Od1eH7h6Fb70qWx1VkTGzYcAYhY8+DNMGGyQmt
QHiZxjHQ2T6EKA3CIo5aeANL+SpyxaWIkElowEx1gZjbVMzM01uVTumdUF3Gfm+k+nBrYbeo37rU
sLNZl9W10N/cLo5T3aBxMbElT6mAMs1U6U1RmHYtrtQudsWCOtozG6J0hj+SvzJ2WNb6yJx+4MMV
UPzl9ffGVFRr14PWAM4sRF9EeujSGJdNbJuoN5cu53K3VYsZnrrc1dr8s0faHeftgR3wKVyGY1lx
FJZkRVpMZi61vjHlvhrjiJymnSIOebJINM0o0qHBi+JcQqrS/+dNSSBh/gXxcP9D3A+WV6VHvL/R
8InvDPRU5+hkJG2O4ttOILzBB53bcfUyKk7lcWPiMMPcZiqTaJmyugZ0NQDAqSNrZIfn+K6YZewI
HKFlVxweXGVi4OEiwWSu8GAmQ/QwIA/5+QqF95kbUv/tjhVDf5oWFQetXH2YoavdYEqlnFj6wpv6
TNJS0103DWPoRYWbDPuYtHg1fq6OvySWzlYpcrWCOQgf/t6XtjJ/d98HwfYfXHt7FMyeWe2ElPHl
S85LoYo0IcXB1tBBWLfm1MUNKfTDoxkF0D8qMbjJtdLz5qT9WL7P9Bt2CGKi4VkvfqRDqWBwPNYb
2j9GfBSzNCtBP8bA+FTvNQ0zoe6Vd4StAJGrmwyz1QpiOKQ+pPL6pa73fcLopBc0G7AS7cXMOkGH
aiY0UG4VClD4EdNHmTppI7bBDdb/t0poDGSkGNZ20VPaOZmpsqP5LayITuZX66bVhXUQh+UaagW1
IQ6DYW07zowqhA+cWh9vOj9KYYEFli58g28fWtV0AWYlOP+S1zzg+SM4rQQbx+rK4R81mrI8BPu+
t5hkizylrJ5kEjt/lI+CYGV7FRMT4Z/GWxFPGu+qkzDsN/KwxtGCJGX/pZsXjsVNghzM7IqhBk8k
/h42uFC9J6+iy+41ro28D+WAsal9EnhArUGrf4kvMJl2FRVPLqwSLqDlLm/3wtBQ5QgQVlGFoQae
qx3ZghrmA5McmZdJIxre0Q9pYxjn3yWHCl4NgDTAm5SqzOXAcj4bKbNdYybcAaT9u/bAgt9teduO
vl8otoJnQAkKHIcME/EnieANwsgxdBhjbkxJ3FOBDZ0xvPkcOsfZ4F3hhMlxzqgvhSp4V4909dJh
iZShi24dKVWCJ0fHKk/kYpuZVNwg3scHtTH6AvtFRzcfjX/mZFR9eZlh9fZIxxmLYHPOIOganRz6
t3m/fG1hg4Frq/HMFsFQ31fqCCqt4wn694b+qsFqr6QCi+JivOMGyT7de/JCsKmrP6h8By+CRpkP
gq06PpLNH5I1DBIAlUZjmP2ZLZxUCbxXXpO7zs7PklmCM3255O01M+L0fdpGP85lbk81Q5RmelVI
gzwBmPi1HumQISf5kX9sYT+UKigzq3aS2+wmLA1N9bCotaND4p4sdtQ5ulLafAjrLuxQ48fmUGfF
ljKaU24A5dg3jRMsDHUlffZA3ijjxM3ouSvlD8omCX+A1zDr1JaHtPH38MvBi6D9mdtfctiUwV45
eHG9H0FpVaVd0PWfba3qPXvzZN8YX2e59L8U0o9ym5zBbP7x8+7CwSZZ81KLpvxTufJjzgkznN4M
DHv7063v3sZiWrmrykucLuAmVGdoZpSSok69fygdR6gSAJ+totsh+pzv92MTBYR+M99aZz1FbNki
60bTPv+7lg0So+vKYqkTekulUh3TNfScG1w3W5RZF1APMhT0/6fyCQpFcbmMWzwyd+mcDji6lmGj
9CGzCHi3zZJcLBOxZTz/n3zD+rbmAD07PLyV16eotlrJ77S8TVyxpltkTHBlhq8xMeOt0+YAnXen
udVQkgtyMbRGSRggU0VjQSfAngbshN/xuWhFLyAEV2NGmvCbacyavR37br8vic343/urBgv4zP4x
R7XYkfa+i+J1cOzTxd44le2gAQyhKHBiIsAz1V4/iUSy8KSiSyVc0RlIHcLwXwy4N6m97iJeYwhU
6w3Lmn4160AT42GCW1H3EiAEB7U4XFS2a7HM0mDRTdw1iWGfKB9sz+kMnqyZW2ehqvG9E2CDChLW
gBjCiT8K0BD0T4Gw+4hBD2Z2MxwBWsh9kax0+hZSlXl3nFtQ0kkv6Vd1/6D9ZOxG9RwOg+OctyAu
ie9DEXcj5Vl6gyjaCFHL8PBodz4hvHdCWH5VmMZ7HPSPbbwZX1UMUUvr4YxMeuA6epVqaWZk5jMA
VDLHLmYNcqOzSpP73j74iQP0td7AJSygVMyQRjZAm1Dd5VhXE1rLWKlG6TDNqHBbvDtNf2KxUAxD
TFUfbaS0YYHPl/U4iGtISnOQsUUsWD364m7lf0MeJ19Dqffnf+O9m18xJc8PFXJiTwLaDulE5y2H
slGkoCrwHHSYqKEyQuYOm2LsZqfS+z6BDCH9AXWZLOae1drs4cRMVuRNtJWualtkCj7NmzVcNzY8
Aoak8b7WyDsv6ifRofonutonE1D+mUWFzLzBI/mUOJwS7pPztnZQ5sci5hY6yDhije5pD7ApMjIG
fUb+VXsaiXrZ6e3nF35Pq7GYgE8M4xoizHduGLP85QsHu2FAMb7ve1bR9ugTbQqMWmso50whIaHI
PALz7noDJ+FimKrlQJpcqx/djnUPrL4zWxKQzhd8jWekqz//U1KOSmibQYqx2dssY41GOq5pXuPq
Vf4zE4FMlceLpkmWzTnXfEjJHyNggupso3VIoOUGH3Tm+CyOR3ZokapLevQZ5PIqZ9EfgW70pq/x
O4J0j9rhAPiD+d8R1aqF5ag+Abt88JzIID//I1y0qiaZYrC82FiiDMrJUjSzJJdTaz0mCpAQyGfl
9bfjEGyodGhwzcFRMs+D7/bDq5Qra5RqtD2ZLUMsiQl/BrF0CzHUcCcHan+3e3z9LaQgUP7iIX9A
uysq4soQHvJtDxCgvXdv3jbjjVP8Br56hFbDFU4zVdKwXmXF2b6Aqxk1lznARMXXG+uZ5ByVf4I6
5BdVew5acPJ4LH/BHErnNN5Uh/xFqOYcdtuMQ2YIViJeRhetssvezSmCrVGCBDLeQQ3QnXkBLKPH
19wX3TyG4honNwLYebgsXSulkwfLZbt4Mb5HKdNXcsPaMeZTUe6DuygSHTo5SSnuoe2cVkIQ0aZ4
mmx7/D/ZHYl+VNQvi/q0qOQw1k5uPse6lE8Nx+qTuNVYMuUMUGuGYKuAyJ/zxhsrGCcaXkKbwGDZ
hLTmYwOZoEHAmmhXWyj1x8QpYZP3fkefRAcxAB1vwJM4/jxymiqzby191e4iwqmHMmtnbD3n/O0x
R4jmIQpSGj4/E2BEKAMQNqCvxSvHvo5TmvZ1MGUQVf3+Ei2vHsdCUNOreugPErYB6kGeRKZAj8lB
WVmLrGOqdxqhJx37BgOYPQogVrjL0Dt+W7oTPI/u/cMwqaAZbxQU4bn2rGVqFWt8aNvc786ewqJ7
3iNDKwo3PwmGjBSfsa2ewvNtl7FczX36WRhI+PBBZnUGGs+NfC5uZmLVL0Eqa3supBJLGkjQfrb3
zWx7IMDu2t9uO6BjbRkyUykjyOj8oj1fMkYgJFBurIwYJc4RC2iYOtRUfyqY0ugFhzQUoeNiH457
N92qI9p0r5nAwQ4qJG+C+2z1QnxZ02AgQVDpFKsv9h9bLuDxo4OBzGXmAIG7m7LuStD7pryNsHz9
0njr1zpmlrk661YGKmJJG9w4BmxyYCrNsxnaVikttUcYPG2UpaE54JBD9Vtfq1Im2Gw3NZmqkMVF
MswLR0sjbTWPth022qWNtlku96WpB7nnCM+dvbxl9IbSHGd0dmFwdTeQ3msX36Zswrw8Di9Z6sOU
4RrPLmfh0VLjXk9FLwrzuEc8BHoj+YDIZluj4seceJU6oy0VsKV39mR97WBbfKleEoqcQJjjgDsk
6JYBIth0ZAAoQAcZNqeLkgNnB7nwczAosUAYngwMwi0ehBZ3evMMqcKz5N6CC+jLFq4154YfIftS
chvK1rmzo6NvvLRaIIbIDTYdhADXIST3FykEnQlMKD/r6ymeY6clF1FZXaepICK6hblv3boKOZG9
tyiwU2d5clX7UgKh3d1ROfiXAiKulqN13OxbiRGYlb1tGFSJ0Cp2zv4TIx0AffsTBl7fBgVN0KlX
iT+73TFPMD02ZWFFQ+jZjfS6qkfIfwviVUy3DNCORPnRlLzbM0cJRfY5S6fTnlxP5tknmlWbcECf
Se/LK8ceBv/HkiaoqLM3bGNyfihY24A+I0oq72kMTplg6CD2PuiuWtgdCkEDnMzqkx4iWDuFGaC8
PxrECnqOU9DJNSaeowtFa2LBcgW+Ndfc+wT7nJGeQZorznqRBCjhhHrFE1V8fL/G9KOMIDs03eQH
HjsiU1DflChygOBjP85KCtZb+G14YZuSHUwoMC1tDUor6XcaI9feyTEc1S5/wPa9ZbgdUyw6IrW3
dsuf4OIehjMMPt6xzMI+gjZOUsXuyON6JQ+DsWHbPlO246KOZ0rc0Wzqw8+toUSMN5VM2Wcj98b5
V16GSYGZgMb/2qV4Pz80sGUxwT0pkCvKWFMrRLRqHzTVeGJMB2iHeQRSCH4RC/Vp1NXjBT2D1CFq
ZVFP37Bs1uSmvHzJJBGHlKoT3h7AEYqkZsw86MREQQmIdTG0XUf1G15jl+K6v1ULbb/gUzadm/Fy
HZ6npZashPAI94vyUOSLqmeiQg3CnsBFJRW7BC8tW7WyjC7bY3UGvbq9tLSGHEPMjnPadxYyE4fZ
l9W3tlX+h5lcc9UdP2TVniUk2DqWBtQR/vijNLVCHyndz67WuZvAqh/933YLQvP+NbhDeysX0U++
Uh+w66DT/SwZ4FZLBYy2cbLfoCcQI4LGGOOZnIuTD/hIXLpcoL3SLxjxZjZHYSWyuVuendiT2Pfa
CDw3rM8LuxYOfqqinNjqWQlhtaS0c0IXpuUoWP41iC0OykHY23qJ0O1KcjAQn6c7D1z2/8txa9jO
7yhj0e7D5VDzzFnb9XJivR2oVQ0NUokmx7hW5LYVs+w4XQTniLV6yQwMgRgnWo2HSUg3mX6WU8Zx
FIT2O22zi2HPcUvpUL0ijZ1dzrLAT5nBViqYSFcxCnFJ+1vLfsuddGyGyzxkVsaQ85tpmgstmNLs
kxZYZ2trc5gFmiXDnMiHEtF1Yk8yMjAC6HuFBkwTq0vEXDPecp8TA/lnsC8Yj9xUzul0p/t8Jm0U
+aEBaZTgMMqB6Q8NdzmlUPokRzrIvbE6VYRWSQ8MJTniwjPmmiPz3egM6Ff0EzcE5hZxONd7nVGD
LWG/riS33L3Vlq7hcj9/4Np9tqv8guz2e5/+fOnVuCJJZypB9dADNxsWSVT7CfRxKFR6mnUUlQ0s
+iC/aOOWG5HLzKoCOnd3fdlKbwguX4CYZXlOCkI4cDvelkjocOJwtRbcbsQfJP8JLOxg+T2mJZUQ
1VUW46i/fQoVYIB9fflx19blZx3K9vsZgg81cQsOieYDio17WuP55NtA1hATm1yMmHWq4i4X5xvm
jGuCHod4XDjSIUm4DaxBhxmflnpQEFl1XJ+DKxlCslLXZduyjBq9ZPXb/cS2SJFKmWci32puekx6
UHfj8Zx9vWtd8h1IGsVUIAMllMOzdh09Y/8PD46upvr3YI5hSW8G3XmOt1UIerNnZWkyoCxqd728
pjGTPZf8KCX87ZA8suNCoIGixK1cAuIsrlBgRZ3m6xc8tD8BAmXCZ3xfqRMO3/r+PMTBzoUyLHNz
Dx2qH74zrVDWBBxbbpZrWWmHbb32e+jYTfef2bLL4ppoz971jCj/XpK7PO8n7NXB18IJ+o6RdGfL
Ws3/vA2SMuK2qcb0xUaanBGyAoaI1G2d0KquTsMywVTop3r7K+4eQ4i13T9qTRuXv7pp1fC3roV4
GtkBZstLtHZIXutS6N/8EWd2BM9Lf5Z7FOHqQE3lNIxe7SMNLx5guTtaNfvk6DQ1F7rEtS2WioLl
hZhKZnrF2qqSkd0ZfCqRtmGwpkF5F6wyNt6HEcLm1AoZySMTPwkIy98gISaFPlxy1BtXv4xA6Wdv
i0TBQ8JCjU22viv4MO8IBNAaFnZP30NwgqH5Wkxo60S+UtkziQXcPLUQJNNjl3Ey3jZzZFsc+iWl
Z/tJ65aAX1Glc/xVvG7OEUovRNnG/AaH8hOrbAmO/81pduBj0jmiPcw4ULjfzNR0W8S9tmXouy6M
8U76fbnKYkA465WhWmz1VdQz4UFunSPTsB4l7wluNSX0LrQPWahAkRFfCow63oNZ6DDW6N/4j2xF
BW8zDyENQUJRWULCzg3qy5JCwtL02l6dmLVrbMvpprvQyDARjVR17SWMiEDa8Z7sBj3yKZ5Z0JCu
VdllEGxwBdwwI98SZyjcfuxWIF3Oz14MCZfkD+3f2CGAjMhEVFHB+Lm2f/Q3ATee6mo2yDf+FApV
JqpdrFsV8x85nvFATAAOWgKM0PfWNzd52a3HDw4foBVoGXXRRhOIx8y9QLLyA3jZcF/HWbbepwIk
gyc4QMYhDwlqQZQd29ScUzNrv4rWUtVqyKoJ+aPQrYPhGTYgX5TNRwiGf/kYNyn187sSZxH07iim
fKb3ip2MS2F2sgcVESeNKmnF053tel9rPVScIBdFbvDxEFl/5+g1kBRP1mCONR+GVZnwTTNToT/l
1dng/bZBVz0CgOY5FE4BAIl9zX8IvD6PqVC6dIi9S7lIksbZjeTInTuUhfLY+PS8zKdMdrhPnehB
zyyJ5C9JEGJRrx2het5M4lAUMVGMZByh+toH0WayInmSf3N7lTm36cX+/gfMccEYIuOuRskeYnPn
5zvmpTsijCrM1OtXxNW4gKWjLqhuQTPJH4KydJ58oKSKKm9xPGuTTYLmiYBCQYxrom/iehYQ0Sbp
miukaIs6S/7BJZlH1z0v2hIIN5qrjwaBL/ICQBwCWFSq/lSKBly05LcZbjl40K5Q1v90SYYKDgF/
qEqtDCru7SJ3IKCt0eqceDwH/HauWANgIt+dJTs5Im93UXzNw8QlDNEMPlptDPDNxpgau5BALSeD
OQExNPFUQJegx+PMf41S6p3OvjXjvCzDG/7meRmhAvONMho2rSMKJR7GfWuWlHRKbHJiczuspxnk
lHmqMaeoe1iqyzhrbAOVh5A7lLz8GmI1jxE6uHuF9pf+nV6Z0Lxv0ZBCViMl7HZce7XMIraowzf4
FqkAdEFO10MW3KGGNzZ1WMbJiLRNhfnEbOpESMkP6e8Izvp3gx0BvIeCHAQYVAaPv8ouPRkQSkXi
GK9esJmre+Y03U0XDkLSL6qh0is1/PloLc8Lc9wdLg3gW49/lzeDC9N+jSb6LtA1C4n3q1SvCHfi
HhXlLGiQOLjOxjTj7XFjW8Ogr4Z1aWCoQ0NASJ7xE9rIzf4sZ7VhvX28SxoUILxwFIC/B5XU4rsg
SZHrEVUCVGcDUOmTW8Sz//+nMEGU0oTD9joitpEWBxiPzq7BsalGXmj338ikrAvNaAhkZS/Iun4I
cX+Xmz2K3OS+iWN450M607SE58mI7ipvvp9bD++PJmcS6Sx/UU0Rxonu7/DTXgk/AdylqbjKHGeS
31u5V8/psZcwdTyMVwGgCgQntObPu6w3xctyn/KXL21TAkmpa1hWEVU9xQsTt3XN9X/Y6stDCfsv
zz1OFBAboR6J+kJ/tFsZOMh9we5ZhoZMAle6JM9+yV5eo9zbg5Ta/QIbiEh0e1lGxQ/rnXtxvIPN
4lwIYicuaggvgknlc4AtBjmxo/V9KwX0sjcbKoAJ/aH1oX0UE9saPQ/jkEeW7FTay5JazYEpgi1C
IUQGRRKob9ufOSMcl3m709aeaC7y4xylh3vZWjf4fcSwdWH037idLHWSIQSC6W/LhcwDa75N+QCp
94xM9kV0pRFj4iWrPrwYLex0YSlPiLdmumBYI4iKQ5i+qKIuQ3G4Ut/6+msKuuIsVkxKw+LOOHgy
0vhTNB5E3ygV5h7BXCVhdP4n8+7tQq08wuqsHhPf8JvZBV9TpYGKySHz39Vcfns/bsR+MAK2up8d
OncDHSWfMvlu+yzH7Oxvs4Ixv4EclJAF6SmIODzJZAV2fqCJz5+8czqmy9OLXGOPFZY0IG9JGJ9j
p/BIHrFrRlK9666sX3iFAQZ3eDHUbi3E3bWM9gbnE68G9m6hx1zYZ/ng9uRq/ej3isRIfKIPyvKD
WkXaxCRzcTZULis/EPSC7fQKSldnkTnTbpbkU8EPLQE5/2C11Ay1PjigQMLKiBJvlShYx1gxZvf7
QqU+2HteyTm6BezJYE47i+PgYqKF+0o5jfLgdH51hpTT54Cp6iRoAHGx0SlY7R9D+adIHivv41e7
GH569Hc5+DsM20KGz0CgECkuiRdb0Snn6SjRekdK1+rD7BuVYBcx8Qn1UOuqzZbysnpymli+gjme
G4kKi+lofjfQ0oKG6PWq+rJnSsNOkOw1oYwx2sNpIiYrqC/JWr5lhyCdQIxuYfwQIhtz3+Bucurj
zwHPi+6kZO+9Pip2gxq5TZuGLEr+xGI0cDENuU0tbwSEBqOBVhmKmolC13P4/SvkirF5cGnaDyyr
txuIyexgxaN+/oGxKFNFqH5EizdAbgkRuRxS+c/m1CBaeoPO7bD+lv1AC0rvBae4bikfM7CDt9qh
OrgDbWN4B2uxE2ozo03WfS/ZLQzij3kPWnu+i/KYCwq4KyWHukqF05u9013nBkGW3ReZY6TTRv++
OW9dD67FuVFz2vXJFSb/WQ4sLLqVwrnNgWoK4UFZ3bzPxqz4jCP5X9Sntaev7v+pT5DplGN++NpM
JHOi3gTpBDX1FEbqIhHR24nHIQ9uZrKSTfw/xoA3V1gFWsCBz5YHBfrsfhyA+MOYXfF067drC0Gg
BZZNArBGSh/pQH2u8yMOkr8V9sZs/EDmHByYtQPL9v5syfgcs26o8NptylcuyQoCELi//+XIJqAq
bS/ZDA81SPNllj6P4MWpMk4hEnTSLaWKoZceAHtnTQ7dw6BVFeejCCKdR8fz7BOUZB3vEuWNMVyl
+LPMeSxQ7dJonJob7y6L5dE5P+EzZoAG4zM/0fY0fVw3e+malquKg1Pot0MP7HHvdU5FTnVRWPyE
amzJn7GerVuKRrb2NSx+PG/ljyoYozphmUMGfYsmks/8pOTWsYhVPB9cNTuQcOFSAiOsfMnodqCu
BAdlsffBv9yjMfOwVbKGJs/Dmx0e4msrCmw7gYDd9+GNJnh5gE8fw5zw5oYVmyRgD0ZCZIdnPGNa
SjZvnUp3I81TStlSb0zPG1GcA5XeGQ0bp6VF4g3MpuMg5YR75hgp0DiBdoumA00FdhY1xJ2tQUeN
z4nnJZN7b94IfR5zFLI4ikikN97aUtvMIezPZxc4fVFRH2bETtG6U+I0/qhv+Trh19sZAvmnAcnh
NcXojwtcQTXld+DuD+UkIdVmHuPHDnoXbclITWr4tEA/apKR62W7FCPCGH8zMUqY+5YrL93FP3+F
1ysCrHbm92ZnXiUotflJ9a88p4Ib5IO0xG9MR5PHxyGl8RxO0xaiulyTF33xXzK5LKHYp9ZMNyfF
EJLaAQ7DM2o8hyDPvlz/W/MxCWrW5cEX32tIQ1LBat75faBAdj5RxWY71cOFuuvqkWuMhSLWo9z9
agdy/4f9JtRyMt0AaXSXxuwU+ln7/ZDC++xn8MU6hpfB6ytydqouQH9svxLvXZn5xlnEAmpjf578
f5vfYVgUDoJTjokmGAwtyS5ZrG72z8XP4HUGLwpRY07GdBWLKh7/yDeUvPLi6LhxHHEHkrx+t1TK
dpv+gRnXj8WyG/3NhjPGVFvATMiRKE2Sy2ERE8mMO/hBmwyYQkL1VWs7NKSdKFplWaKNeFwa5xcF
kdDlmvQvAqLOxNI8tVH3bxRCrQo8NOx1p0KZAHEGH0t8la1/tb+GcD/6ObjDA8kPQWHA7Ve5GpWN
JJDsLEcvJz2425HEbrv0nSgxe1A4jCXD1tmRbmBd/vJbqvaljzJbKiK8skZoayCjbT/MxVWC8f7E
mmHQZQdedsci+UhQP25sej227eD8XOI/gMNzlUk9DPoJfxSVvtP/DO8q4utvODFLfG+xlqsldVnU
ZoPyrh69aEQTJp0+T3ga1IEHXq/r7qm1HZ4J0yh3QuCC3N8eogzvYCJvMo5lHpOhTQ+HdqAkFX2K
hhScNmBNZTgtvPWU1bsa0aFQ6e0Iz8POfY6T4y/023V/t5Ni/J4t+hMKtKdZi1D5n4mSA60bZT2u
YCU4yZ6XDkgyMv3TiDEU1qmqqJX2VS7Iy8x3FtB8f90brFr8ws/ykF/zp0k2H148WYHsd2Qw5nLK
6/30T7xjz1ZjdcaeRn42rVmsWifPLv+Mc3RSg3BSCFkKJEQ1t2cgmpFCobDka/HWYC8ZCdDDDMmq
m2aLqxXnAyPV5zarsosqNpSCle/HltiobxdAZ34FBo3ncTzVFsQswzDEcCe2EDRwIFLDKRrxOzRb
OWzMABDphgkzDOvSs7PnePO5YTGnjfpLdIubyaZCZZG/8yXhi6Iy/P0BIyy6UPp6Kc/YO4zlsB+Y
3Be3RTl1cLEpG8/yM5mW27taFeZELjXnAmeHJprzm3ZhUHXQ4S+rzSS+CKmNDTKWAApTR9xB8HV+
6xWSHvbtc36FDWFQ0pgNLPMsFqrcfLB3yrwawF4vU35wvYL0nW57gSYhRLssMj2Mkf9bOEVhx36/
HNrPiSp+R4HrIdKrpNPEHEXrnsT1F5c+rTvBGy2hKjkbgmFyUfCRnJRNZokzk2Q/L3FcQsnL1lUp
GAH7mRyTlaM75IUXfGAcQ50DpPDrLHDJgBBfG1JECv1zj2pTPA/xF9dFbH7PwqyWPh0p/ncDYbjN
0logSVl68xcg9XHmvWzMGlLJvfNdZw85B9TFXuPnckgzXvywbFI04AACPB7dq7LPjzJas0c4zKXk
KR3ZgcqBOkjK1rl1YRycKiS1Lk8kzIbDE1sk5DcARTiBiIO14NW3xmIRJYNNbCQ2bm7mxkzDvUMY
YCtYGBqJ3Ap6+S65fWx2J/eGG+VpCoOaOSEVtd97o6sGfiKUwapn2q4WENnw9mAz5tv74Td+XLyu
cokx754F7jCwcIj4eyD0b266UO9t7/coCiHObtUulD/0f4jdbiRST+o8+vzRlqKdD1EXY3hDgNRz
3VE+tT9zFrDobL79AnDl3Jz3vmlJ/mOTDZXj7qnh8/K1xMcoiA1sf6sN5T82kvDOhluMKovp36Tf
CKt87xywgf+j6P0vhsM0WYJXb8qdD5VY7sPJmMfP0qSNijp55d6+QrQMANABh6a+vz/E+PNvBS8e
EeCEdn9gwCvAK8FtlUmIp5TYJtnE0/pBD3TcwgwCBwDYkShAM6uAsFEWd2/14JH3+iE6BEsZd9EY
Jsp6Cy10zld5I3RziElB21ar40Hkgc1U9HLAjj1XItwR0DJ50K17fyTjuVnkVRz5zGdpRN9wfoWX
i6M8M8/N4h0M4OMbnSl8EDKlyZx/Np4gia7pfFMfthXu0oFOfysVwWqcroygM9+abDqImdWDoyg2
HsIqyjCKKm+0nopFRk6gDWQDThg0BXL2ESH8bPoroKy/Ka5ZtK/7qbH52pVHbR/kPFnQZ0iTiLVT
W6+ZMpTzI4W+9aRdl6nXO+x9rBSxO8c+Pgm4Fa/DRxy5pQHxHP3G6pPiQ56BbyE4AgrdVmhRVAO4
dog0zWNbijYH2OqJt4SXzFxweChsnKobaZ4voO9FCMRMycATbdDjpi4cHn9hRhnzuAs4JrjZWuW1
n3N0R29bogsgIjotx03Oso0ZYEfKdoTiGN0nCISEJ/ygifB68dlHkObkmC6bpEf4evqlOaf74eb2
F3Z7gCMSVJpL+biogmuDMo8C8sOYQPMwmhPqVQhg4qGmeS8/86TdP5VyzFX+KT4E6v7foEf12cjY
T4vgi38dSJgKJG14cTt/bmu13hWhdoeQHaC8UQ0G6OPR/u5uunCkEcgZ/kAwU4GGmTPp+/Jojwu3
BAKNqAZHvWp5FL4N+DUmVJJTecnngEwIjhYjio1hRLwBj1W9Kdhz3CXaO0jepNou0VR5FptknXkm
6bISA7a+N2qZ9pa2fafVKnqLLoyt4S1wD7eRB2WcPUnVcF72iMU0C/a8sGD68khuvqoYEtHVxGaN
8uqxvd8uEkSSjjZ/QktHr0oEjdAInYqgBmWfNboSiB5KWQEyXqDEGZ5DNrQTcmGLZzkvsF94tmug
WOLJ9MZTb8S/sGGbuWKSO1Bl0JVjVclfvJxlgdzuXN0bnJxLUZGGZe7ddl1iSqVOr3VgUpmTSGB3
wgVclDdKMy7/ueNbeuOPWMcQWXMBjtyAJvaPjwIeXIcj6RA6EWwJuxyr+jWMmnPTywp6HF0R3Kao
QaErtYH8keI+nXpeKsjl8YklVTGOzpgF+N5uXR9jXab2XOFNXpmdfbxH2kMn13NfFfD7w75fjn8k
UOdW1RVv9J0hYEUdrtbTwH+GHyyo7j0rqyd4kR3XhX8kEhubbZGxRRX8Me+ataYAB06+q+VkyLLj
vwsMwznatM4R8chUczNCQc3xFA36CpmxYOhu/jyHJ+A9ObRH+UY9frghxaS/fBg+oHlh6SPk3R0p
V5ZBcujZlWxtHZ9C7uC/9SGIad3UeDUhfy54G7mnHl5+ZKha/iqwUZZoSNZc8KP03W5UXIXcykh5
2WOmZNYxVMhk75mLWH2wQYCofgrRi9UdfmqoZyLt+0nPgy2FxqUEmH9W/7Zgc4ifnVpZqumps4tB
J9B/PidEh8bz19K6Y+tR1Z564zGwGAEZbbSx8d7+VYBJifh7dhIwifaOQx57Ba/HeOIjBecT1Fod
l7j9qHTN9VlMoshwCFy2lcli4R4GCFSTt0txupv/xrWcb5mLPe27+fP5bYfgNJMegIMTbxel2RE1
IZxizJyFuaFVUETqzGY++cu4kJCwktLt8vk8sl/4eLonDbSmuGWKwQpYFJ0SYfVHEUMwhwxRWcfs
wOmgj2K/ORVpd5z3UVbNKPt+JwYWHVEdtF80KyPH/a4w8uIcrfC5BpcYLilnwNMduFvhKCdN99xr
9ktdSyG1KYrvKMyl6MDxze5B33wmygQD/LUa2TjM9mvEp03hBm8TtL+/lFhxnFL2LslbhPF6GOGL
v/uXSQ0rKqkae8TdHLi1qXkWrQNlG3paao2LAQOvVlJvnvtHzlLDusIH5mkaXnkKDLa4VhdNl164
6Uroq3Gj1UtCMiaeI+wkj3gUvubHBGSqvg0SuJPuzf7C8ArWTtFwhu6bVxe3RKrLX2dfvS/ctqM3
PZGxmJ30MHi/NNUzT8OWa/0AJfAyt/SLzdMrQ6PcuHUZJnZRmj84iAMRuL56NC0p0tzvoLgQtwG+
FIaU4fTzPpS0nihbjUMJ0zIosf+TP61YidC2pcknz0ME/eLnEZtejVzrxu1SFLi/PEZWooEAzNw4
XnOF0oZ4uCO0FSxB+z+jd3Zj+oJAxgLRXDwYlk2ut3pEMPTinWPEJ1IwE23ty4r6IOi8N8X/A25L
my2CP8WbQ0ywMmvz+cncbEkK165Kqm06c/qw3XpZtmbRF+3MPPEq46IpMZiuwbCJNyvDJKHj+imc
DdIJDIxzejPit1lPPSA9PRUvcI0y7MDco9uDu2nFJ1gxa/SfPUGi73EB2NFzS5AiqT3OXs8jVF6G
gRbHvOQLsRzRIFcHqchFKytv+ZxEBIZzc59BD07x1/2Ou5enlV5O/HkTiP47q1MJb6TEzqgsjWNL
g1bd9TI+oMzw9KEZbUcObxUc+ecqdHOgzZfOBuDBCx7cS/VEovZX+6d6csS2eJfjq1uY00OK9yZ5
Ri3Qxfc8lkk1Qot7N1+8vd7kVsF41pd2yq4LmwhqeL9DxV/KMU9xBzM7BUoL3t+h4iNcUPSuC539
GjqoCc309RobT+/2KyK+bGjeM+2N2I9AYn9WI8X7DGGQkhCdm4C0n7z4RsU1FqUpteL/rcCiRnHU
+t+ytcOTjPUOVktgGPJm0d3Idn9SlHYVptTAp1hnR/WJXDBLRAvbyvEzSUVvS4wTaoFLyAXwzHwq
EP/N16o/rCZQ3vF0TRR4sw/Gzw6hoTweCT+s+iyYvUXqXokRkK1cQVx1ErB2F5WZ1bY2gCp4VPdk
sKQFku62GtcAGqn8XGAkM/ndKKSp62TkM1P3tP3ISVDNsw650NyCcYilmQ72YRSlIM9+4QP7w1L2
uelDNcvEp9PQesrDeMe8QgQLRW/PwAf0wbNoRjJI2+o9/bB8aMmb4uffygno77P4GWeGtPm/K9iS
vRnzJzM5//ZO53AihPHToahnzUK381E4EagZsPFhNma+h14mFWjPM1FuVqDjy1UHuygqLLZYG/GO
K+brSwdsXUyHbVRQ/9Bgi9yd0a+FsvZUEYaYWKrIh/Ywhqat6f1nB+cBDY64EIr1ziEyB9oWzUwS
PL7fqLIlF1RDcu2M10DRTRGS5KV1loDyoSxgGyFdm4E+IbSybSQ3Ci7Rkf9FGvhLtbhYQDKOEPVn
WGErO6sLWED/zYStzQooMHDFomo1tZrBHTx+suUZF+TLSDDJng2/ii4pRLlSTqWMfXGov4hbyaRM
UJv/adLCs6aewTmAfe3AtpQqBNIO9sa6CujAafNTb+BNlzhxRba6gEOl3re1pwu12w5R1p2Dskta
irSjFRJJUdIUn+HIl79ZbMVRLbpNGAc9wq4Yx+Zbo5GTnBot5itWJD6IyNzgD2bzCg+EU9EoDMlr
z3ATBkB8GP2RwMdJx3gkB6+AU+78zkOxtYe76ePw6Ed6WWkjHceaaohAmzKVqnf9AvUNblIGgCzh
07Tkgo+e++reSWaP960myrMFqV3c7GKcT45AeDm1EEDvXtlP0eduHSMSQYRTKfJ2FANou78QJPv3
S27XgVlcVGoyi+7XgOGh8xYlAA4ZYMZWAm6Ta2ZUE7jsNP0UanJIOcMZtRghijBOYFHI3/0QehqB
gTQ7QG8/m+weMqZTfuC5OASOMmmTOZnUW1PIlJrXhAw7WBZXN8TviwtVlLSA7NxaD98S6fwTW0Ni
G9m+WkOljhYcleIvkz0WCAwO+A/EyK/8EdoW7Jvm+Bi3L/Bse4i7q/f/q9sRxwzBSUGdl8MPmHL7
LkjGnRK76pO1PWA4A5aIHOtvLo4L2aTvbLIpRsLhA0pRkTt9f8IXorqb6LyBoDe2DifDcxVSzlnm
tFt6DYQDz7fm1x/cAKnWdgN3NoiR29Q4QG2YNDZIiUkECG0N1BSLpK8M71fvKHhYNYNl3M7TC9DA
6bACdJWQdt7Yunr9ePOdJtuSTQ8reotOTjDcOXUJgLZMAK040J69wCz62z232X+lgFGvgLN3GZlK
22Ntl6zieCl/XX3AT4Tm7tpXBWCk82fG2cnzEFKIgV4A9Br/Cojddg6tEBK8PJzLuOa3rURnRFAz
4CQpT50UpA31BgEjConnEBaL0J8721ZkuZNJHpYDg7JyOls4Bqvw+Mfm6FSIZZYif0yvahKNHB7J
A3fnelFZvRCq76iMWDPeGHGAWLvJ2xpWZVxxHs0YAatY8y86ZPqFx2Au+YkhY2HIZDWs/i87zuSM
HIzYL286BJMq6RkbiSxKhU2J+TBJJjJrYdD/2T4hzKzva6G59qM/5XACgr5Kj8f5f7EG6qWu2uWm
hcwIfcGMDVQqKYWUVyQrGyAYTBSq0XSBTR5L/9BXiUSrshKV6azbHpgidyHkqwqwSeU63M6B3WT+
rsA6veXPWeROG1BqzUsdeI5peLLdrTf9xt9y+xut4FJjINgQ2PH0PiB0L1XZctYOnHfzhaBSs5n9
0tSp926UzvM89zb0r3Vo7Q/cvatvmEaiV0iqRKQFt3kyaOLJ4dvNCG7ykXI9TPoSZEjVXEvLa+hp
0tZF4t0g4VbFvNl2FxtpYLs9zq5q7MA8W1r7VmLPVTKk+VPjz/fhk40QTLPLmZYPJQ6vdGmOKT04
XQ0wkjrymQ7+cpGCFi6heGiny12g3cl66OTg2+k7pJ+OIv62mfrTb3Vz5avAT9lvczdcmzLyiIFK
GTXM/KLNzofl1n0H7RLEVXl06v1M6EKlAwk9R221MuuMfS0BuAWr7iPfxovJ6+hK3OKYMn3F1LnU
/8PMnX09jmu7/HagHpn3mtNE9gJJ9lh4Gzar8mPaCkCSKgjgK/9O7HCazIImPd78HeBr5IA7jNBW
KjTsTrII/i6j/NbOogf6e8jnAKRMGK6Ji4qxDaaTHK+pGMMIAuoMaclFLIPXISy1dbRGU/CUSUkF
MXv2FJ3nEIv/6ZUqgfYWa00nxLq/bLKYTsL/cd9KZO/+BdxPfLuNpliHAYp5jmbTxaWHBu0tHokL
3mmloioEuENu42gx4jYRST8CjpmUjX/+ZpuhvfQpPI/K/UuNYTzsQOOlUFcfI5eQAlevvLLw1MnF
QRya+D+24IGq2pQGHnsnBI5zZVQA2ZIRkSV+YU7slWtyxtKzyKIEetmkKyXlqUXBVDZD7fV8hIb0
zlNo+PrO79HnTnm1sIqaE1G7yhUNIzxRfYKCikcSs3890Hxzrsm7BwXr/Kos3Se5OrnDTVa+EFJD
J4kzGfnL+ssA2ivjeOT3eQsNV3EiszSYhlzj7os6T9y2DtDQK8PyGaW8WbMLhAUTsLNp/elN9dkz
xq3AyJnPoMARTHoEENlm7x11GnYyvnVoqX0CmWBdy1vHf/iOgtM+HBXY4vptfv5BHvyKU1LPMyH5
MTzweBYuh61wrDnB4g/+tvjYfFi4s9pgoTOgVYih2QXYI8ogaxvs7Z4bEhu3x8L4JszX6RTnlDEs
36IfiMgL7KnmXwx8KfO44otwQmJWPgrvllT1IX+PDgKV9MGVJcsZQbeVZ7UxD0Qro98umFcoFa/Q
RsfhBXQCoCmTAVqdBGRrKFAOPoON7B5++SxhsigskxDbH/TbEgSAcEIp0GiU/pY367Y9YXCbmkPc
gmvIW9O2uMCraqzEQPQR9qN07EGcgGZ4nrMnwMoshTQk53qE2L1je4QPkRI452Z7PTZDSMCyoJVO
yJYz5vEZtRzgNiiuzmSfeizhTPO6bB5jspqpCvTGF7a0JTgBBftJx8DnVsqdEwEIn8SIWuZ5+b1R
+cm2WLQqnIPgRhaVWjwT6ZdKc5sGTmNM2R36AO+U1jYdLemH4uQEy8xsaDjks7M3/NFHZBJnvymr
CteyVlMjQsQOncyCmx1h8X3uxY6CifWo4Df0JyZj3pYhgm1BXibIEEO8dsFFrQeeJJC/19Pl2G4i
nptEJn1ywDxdfY9hmJtganqSWJWeA0Z+TGGGqvVQvgc7Yh0ZdllT6TvhoYRp09SKtrtSjPaHbY4+
nFqMU/D7emLA6RthLegmOmmjMkzcjwKrZD4XR2ElFYMx7KS1oyOZPtZPk7uMsn6SZfBP8Ga+sde1
J9uhYPanB0vl98EhBLArs8HVDJQnjNMIVkVsRyT7Dy6FMLYqO092LK18EKSlMgeDQ0qTlFF4tRSB
M1qRuRThIrP5afahrbK51uiGbwIsA6lw6s0vGUpyUOa/c06A3ZvAntQcbL86rQzSNxpS0mqRWOBR
TBq1EnhtxZ7y17W8iBy3olU2Sw3ryX6cuZ9BG8+HZbWGjc8GidmGccy6wIJL8Nb9T/Si/kp3sXXy
7Bh9ZCYLi/fiA/t9VQkHr27hI2zz+n298yZ0DluwPYA2F36FV46WG7CzYlK8LrTxirGph6S78zVn
KwJFxCG46Wla1R9xymNJ/DUz/AH/G7fr4EWb4MFSOAk++gf1i6IQB1hzJkE9lJ5HjgZLdeGLYvc5
NHvyc+c4Prl+5q843jcPKm4zORp1u4ilUyLd0UwoeZ3HD/fOwvQIYAyWleMkjRX1FGuISS9f7IlQ
qKhSW11JTfzhjK0nqcek2UjinfY5lRFJxiPdUVCAErqqr3N1yZEBc0YpG6q+vkho7ABnvyx4rogQ
rJK9+y6jCJ3PUSXXk25HRx7aQrALvj0jeTze6Pn0RmJfV939+ZdwPzLDl7NeVmY/fhr3d8rMUPuK
BZytNnrUTpeS9L+Oj95lhYuy2XcZZKh04Ad6Lq/ypCRmR8rkTqYve3nAHplYPRYTSxOOKYESOSTt
1RBpcALWex5VEEkcgakJovWuRDHG7kknaXx2PEsgxr6C28prHEmP51gFsHOBTdck+Eovsoxwx4la
ADCqqytn7WcvHregEuQmwLJr8odiex9iEu320SP5BcRBpmIvC/FhOLZnbaGhRSRJWErFc+K65ROh
VUgt66bY3GrlkPUZxL+0xsp6lXAWZM86VzX1NBTkKmpXT0a7AYk0/glEM2DdEjq228COoSUzqKLT
4DjqvLxiH+3XHYOARibkHVibaT2vF55fB3Ah9wmVYjH5PbERhadtUNZE729TVEwh31faj8KXBLYu
MH7aZPT/l3xAtChqNdRrHjFRadR4W1STynDXOKwKpxjkdGH1bhLPuiDMihPMPcYIeDpo4FXYfoDu
9Ja5E0zuYF1d/YrgtyYz+pD/gEkhnCRH/JDAfuTBCtOCvvCgqJ1BQpmPjaeR/W48mX/c9W6n19v4
W6Zar1J9qMEr9XNo3AuzFEXKIMNWxMhScLfo/uFmuUWN0VkCF+fYQUeEMrzZTdj4a65kPQ/ygmx9
ABTJhARcmIMItS15PQbEX2dJyowgnGunYszkwOacbglF8T6JYzpqldiZ7wRyoG2rXxB6SAog6yPe
8ufEFpNtCjJUoRSorX74qfcuy8i5fDo7+kPq9c6u4hArYEE3iu6zAnEk6btYUx2AtIAFN2N+J2hT
EfELtYUejIMrM8KClJ/RngH9OZor3L07G4AIHWd1+euBtDBeaczRF8D0KCSDcNm/RNrpPOxWQdl3
ZXgp48vDs+aevr3q2myNAaDK3tQXSc/9OO4/odasKTqXPLjIVNoJYaIsuCOH4+1KGzzRIqSIRz7E
SHLqFWBG3ZbzAih+z6tUMHD8LL1017DmvCYh7bYu/XAfhko0DguYyijIWh68kRlRnlAY6nJ9TF4x
MWYdXpTakBCoGBaKk28MZH6WrCBg5eaN+CmEWu/ouZ6gdH5aoqyux0dyEuz5oF2akGOSAkT8cXH3
yaPtb3r6b0rWfScdpiHQVzrExP8luhvCokTwJL9jUNawGWrqe3dqRXVLKO6s7VmZsPAFSAOVwByB
93XK9MGzdaNerqX7jLoKhZ1OBvTWaQ4a9nWxbc9gzlWg+d1+tjjMKG5rOku/EjEZ47sUoT1Li7Pr
sFFph+IBPtZqeovujul7atwbHNvRRckNXjTtoTyYVtOuCVr7d3id1YwsgUkc8seFrbZXTgBf7+q6
F7JvluMpUJKRGu4iKXJSdTkNcGmWH7jO5jaOHpchBlF0dfz0nF10pqKTw8pPJNY5+/dUSJomOq8K
2sHJc+BDBhCQxZt1rmSkedEBITvoEXI8F9CqHlzCmUHoZxG73j4tyUTUU/u02UZ/oPeR8Isetix5
usOgzYvY8JoG8nHdWLxqsv2YfZTJ+yFZT54lx8wxMvnxEvnYW15CH/i4PUbOTT9FjOPcO448SQks
B2ttfOJYqCgf7OzRfWh32y+zrNaxryPHqKsJVFcCF1T8T5YEDP1n8scw4E5EWax7hm9gS4jyaup3
B/RSx7BuH0Yrqr1HjxnIX8lidCa8VMffbgjDfXXYFFwoYSWVwtpawzN/7v4Q9iQJrOMVCC24sw2v
vgVUr1fa8Y3lgFba3YF0XSx1PfE20qh6dBat/j1C6HnZvWZuKwpdPjwM8zjzgQiNVc7FUENBQDl6
yB7s198oOgJKL8D0FFf/Q9Hakd17i7fT93xk4jC7MZLFXAhzAdEY4B9m4epoVOshYPBo0QBTbiZn
ZN9azZlyy2b4+9C8no/Rt5xtqfHhzcJ/54yOQLbjso7NBUwgyCv4JYmwsvq0+Rt3JP67qEiZFqwg
vSicj8fToPNjEW/3kw5mTqE35AP2wmy/rBk0LIr+hAP9mshrOHkGFcyTQm8nmJqsnlxCZq3vyfDf
8FOUDIBVi+McLjbjb6/XmGcG4OlBpN55ZWuFUS1Y97uqyg+onn2gr1l9myfHLLTcUWuf0x462CNw
oFITFzPnJqL6Nl87HK8vtyr4U+CFZOvQvoZqxc05ZsgAG55kBw3I33h/QCdn+KxbytxdECeTOy0z
eOPz5C/mmL3yJ32UZoYp8N9c5Msuati/jd38LBBYqqEtu023vXsEovg+hywuNaAOAtlBhUyH0F4a
qAYyIYwa7AkO5Uh+Q7qnDsw7EXAiqwD1lgaKoZZ3ekCYieJdXv+PyrZ/WotpvX3RGLX+ZZ6DW0QS
W6MI3l8nHpMi1y+IiLF+9TpeHd5qdDbCYtOo0hW6Xv69j8n5xIvnMA5YDmxd/XFle/juLC1+JRU9
btLd8YmF62r8/DfdkVjNrcmxojhDCeVgTBLuKog2wA2JYgEFRmugN6l97PjzogK4FW3OltBsro0j
2VpkT3TarqB3rb4IBjb5Q2K1jZbPmqHoaBaVKw6jsqt/5EfWgoOwiSrlncOMbNIRW8tf6iPWsVIW
4ELT17WUNf2CaBm/KS/35auSt+ylNVgeFBDv2K9LSyelD/pIRMgs/T9TxLTtP9Y/nj97oMt2aNhq
wLM60VDFV2kV5MmLeJXbSQwLvDCt4IR8qVEW0UFQxCpj0lt4tF0yQyPXX5+jbbRn5SsYClPV/q6S
i4kUYFnMLVOs2xt5oX1AXXSsy7wvgdmCDX2wVV0kynF8HpMbTrh+aDPIHBd3THYkrUXEsCysvX3V
V1CvJWEnRFQ9zdLURSOY1tVyDvmyOH33AhFKnKH98xOmLnIo9mUrZzuqqfnrUQyuIe7TvYjic7EG
5TTiKz6KgpBhEDJivS/CYEezw6s+CBp0N/WQIrHj6Y1PIZLfmVOzJaOWer8GGYgnxtlg6cOLG65e
H8QQDJ/gU0MBJmWwzV5pGbRxIyPiKkRCn9+DkD5MTUUiZjWs/cEvvUy+oEUTPE3DyzvWX6jJ/XOL
ZGaVeOZomozh5bqsgdkag914RSfef0eHPV/KuB/6Ur/EXZN54famCma3re4U1vsQknjYgU1RKgp4
YuOqu13XUfJyi4BM2Hn1PfuX+sCfD9s8agZNYGSyaOlijh7VXE+WPZIekNSHHPQha33LzYNMXHGR
3zoPdU0ChrXgdXPb6Fq5TP5Ftkc89uzBhcm0Vs0vChtrHnCZjO54em1ISfdSN20YCwJzFRoba4F7
F0cxGuPqmBt7Pgjq7ql4tODLxEGLb7LOyngMakcjsTZB6wBYRLWJtPoxdhCHyE97avwe30BT+LJi
wghO6WkQCw5Yyn1jMph0XcT4jbMhwAIZM5PhD6SxuPKvl+tcmbatKBYNdFr9JMP9pg3K6cH1pGlW
yJqPZTjAbLiVlIgDYW0pPQO+v0/m6NdAnDokkyS32KZxgi7wVZOi8QcsM/mDTpGEALhnY5qnunEM
ltq9Ua/4qljlnmtnIE0ZzCkE2uG1L062x9dfTF2eVE5mFRqT4VrKZXMGc+lTbXHGsQDTQqAD5UpH
8MEyA2mS+/zq6j4dBkMNSmnoQiulUrvwh6nwdLB8Fk248rj1KbYrVmmIc3GiecX2vwGvkj9ICOx5
DvCdZ8UN5781WiTAIySk+MHwnN3e4L43B+qr3tjpzK+gkPJ5FWPmgC35K3mdScUTDZTEOWqBn9vc
AF0eekjNGD01tM4X8DUCKney3rUGf5vEQ46dLPGATEvTml7IETWEYzDtvvO2RknPO+2BfsGaqjcP
kwRyrI1/1Uk9ISGR3grP54ay19sXCF73iMNIz0VXvyCe+dgJ3kZdOHjSed7VeicI9hsQ6PjxaIE6
7HlkAlgrBxt4uBAEDWdVyW3XKKqbN8EZAcadXTj9xxWuNzQ1QY9M2xB33lKIJG4bnY72F0XB7Viv
3GZbsQc4zPlAa3YCuv4EPs3NUQjId2R3GkHpBaIPAMQyMGUe4jGIJEm3epxjUD5nL6BGuCUH7DlR
bwwgLR6wsJzjgIZ2Pys1td9JXBB+5OFCniDNPPwZpwS7a1JWD7viX1qxsSMYtdYKbRu+QFGUspzK
XY8caRWCN4tFxRWkfHEXf/QvUYRvCOuFSGhfD/NewnOfUIoRbRzyR5tAt/JpMkEc2owtEdvngQcx
3chAPzdv/dJBsgQ62sHD78QpcAMvTiAibAAwv5fErXjbENSnSpYNBAio2Om85lErYkwsJjeVpBxc
8Y6CS3JS9R07yulxDP27m7d2Ujr5sgP378eTKqHhx5ijLameg9DsUOm6DvCzPB927+pjNJQfE5N5
Caf7NfsKaerEDZi+osyTMzhD+InGl03g+GMZQ0U4N1Y/iYMGH6VnC5MZmIMMEeO7JOZCWygLN20O
iXHuABSbtANDoe55qvFx62vzTWPpVoPJRjdis+d0hrSq3XhT/lRZbOZx/9SJaE06PNHkO92q/D2e
4xMNymWQk+5UuxuFZQ5lTAjnumE0/6oxIWC3h+pn3o3b2E7Bxe7ArrSVOuibHfAbdTfTHlwQA6z6
hPV2a9PYPH8cCZQnLM/BcqZpWaBIshhaTyOYG5zzXITDHnHMg2uIg2SFHfG8LTyn3m6F9kDr5rr+
zW30ZS+Nn+dIFZcYu2rXWoxyIUpMJBFy5i55fURhEwuSBN90YcW1G6iThcULuXjUD+UQNkMw0hEh
XFXILqsoM1M8n0+VSAYy//O4zbSj2FNieuegTA33kO9yL4wVFHbx/i7F9pZV7K64586LPYcxLpoq
yxupDQ2ng8fXyITV1fiaQY0K3ixnjyGcvhIn9dqxiRdHEMBBHEUesV4DoUZkW2HwjiHeejITpBJf
kae+xUZgnsA0LFnv4aU45/CnZD2YhpO/s+SAL448V2vyLAt3a9dysfsixJWMjf3+Csz4YpYI5Pr1
WfGGGIuUn0NQL15QzElmP0my4L9JVzKv7fuip+U3va6RJpLzA+mhspwch8OOKypR+KAWtMgRRjx/
O/tOazGv1c8v+emDsB+xL7RFKd2yDTY9rZyZ1hQ9hGwaD9JaG+ru9jJCZPF1HrI28FpyLsiVz71I
rb764PQ8v7LjT0IQ3Xbvu3O0Q3gD5BuGm0wL4hnYVpvhij6HFyUhY0R3NfyuqjuVQ1E9Fg1CIzcG
jrzie5NAz6dLlYD3AjeBzo3nIbeLUEwVYCBQ6B5TBHNGL3hapGu+YaaL03BWmgZ9nVCjT3J7Ey50
d46GjkGII0dVWPLeR5NPu1mj8clS5LSYkMgHEOE2ekx9jFnJgMIom12b0Je1WdmBochi2dHvKLBb
lKMqLGHgCi6Enx0RrhoyfpoffBW8sWv34HyIi9TQXQXhplfuBoCnA4W8MtTiYgnyOdxjjUIMq4Ps
kbkNeI+X8ee/gk5m7+azQNZ6S6EetFdXde0kycH1BMAtc4ATNPtUYJ6HiztHTvxzjtXMdmaikP3L
iq54CFik3jx9OlDdQGjKK2g/93CqywQuo0cQdprDN1Do4m/pkonPryjaTeCvMPi56/vhjw9JagzQ
MX+y6pqvc1eC255UIGzOBtKUk15Dss1iuxi2jB9HzEll46HAittwjrPB9QBk8jaA6i60+WKpfI3C
2bVJZmi6UqZvktqN17XXPvX+EwOloJliObj5m3QCjQbc741xEwlPasGW1mPRnmAca7msJSWTdk4Y
6VE2DfDQBbT65frwrUI+Mzv9ToE+SNO7GaRvp1pjo/wNlKTPMxzGEEhK04IfcCv5QjiOAQccLf/f
cAnOJYAP9sN3AIvJpvRyJfpWs2hL0z7MqMicqMQAvqZgY4KzTpeW1/nBQNHI3SSaj7rVGSRUL1kG
KXyzymaoMU0ScmDKgAOzN7Y7PtqQIcdnS+VJHvx+oHj3iQMjtoY8FmtpF6w614cTZmPAGgDhNtrM
IU3EQL9qQ9WG6whohelPlsZgvnXdILiu9EcSwGrlp8Nn/EGM4gJLpQPlvnMfZzZdj1GpgvoI/C1t
2/29T95mZvUhDTzsZUqrrJ28TKvIKFOjaNF4RodpzrYM6ghHoatxeLRCu/sLQNts7LT9SuETQ4Zs
x2LyaFkFGIRuKDPeXoHx6dS3KacsjG6XZsZ6dgCp9AsWUz4xFTKeG2Kswwkg9QRs/yXmmUSS4iFi
xwQpn1BrLiKkDPLVmGoQb6W+LwM7bzp/6Fn0Qfw8IuhNjQVX3p3NPKHF/6F+dW846WtWym10bxYT
ftEK1b1Lpt+VFc8Tn4KlarCXd4/6fYqYmK1Kzc7QGPlIFuqcJlwPzuXkC6yqykbDYR+tjvyyAP+u
0YQ5QUh4BCz1aGh4vFAoZUdjrgnAOHoxBregOGkvIPRMntZyMTy8069M1rQRUsvZe65rqqYkswv0
/175hHfKU7tlbMWDoIR8xWtiLrg2qRpCo+TB9+w/WvrDQD672I5j0pRKsAji9dOdzTUCd/XJy7Zk
tU8Sv5pw3tvyvUpCfQRcIykC/39XiZAgBxH3J25VflCV+700DqD515ViMO5lAGqwqI0+oph/34F4
ydZ4GFUSIx5joGr//uETpiZaR7azmuvsLEZCgUURCRwOqn9FozoT20vTWr1NX20o/zdBKX6LYAZS
n19GzpXD+YuDHvvIBk8pEBWN1Zrx1VrqrCN3Xt1I8446r3xu5M+Vs7MOh3hpt9F6V7Lj08mTzM8d
LFt+GTUPFexsQjJ/TKlOMZB/TLRDNwYRowzzOz66S83n03DID0rcx6tpVbZtk1dItruXXy5OvCkA
ed16tNQGgJhgt2SoNENfatp1WjDUs3ahAPdhOvvMl/YqgChz0ul4tcCnAu62t8cxdOPzAa2Zo/oO
hZTRQ1CqJxUNNJQGUJgjOL4gU501kD1VZQmYwlrrUeyjTL+bo3IsMs/95vSfbCgSf6jwQt/hJXrC
bUWzyyzXyGSi3Kd34/D5X0YAecm/QzMi4WHfoEXOl3yjRpZ/nAg6SgX+ZsMyLDlOBxueoUXziz1K
WzS25nF2ySasMrwpWzCA9S2t0IngGOMuMhhmYpl9FuLdCNVwxjt5ICgeD62Y9EFltud23MMABqyz
3rPfKcmH3pvEfanESsjJh6/pUJk+CrV9RdM0Ae2TeVlIRMI2J8xm88aMvbLoWWrc5UcpFGC56KKJ
T+woGugl6/cxHFXES11qSg/VIHUVmVe4xmjDr11jZBeMQaYSaid9C9KGkL8BhyBntDMX++80Lwoq
THs4cPPlW/4nk4r7XEwzO/S5pYHiHUPr/ckP7LEHPRdbzDlcojKYAOIHDYvue+PMw87ObdPyRF7c
QTnl7OcULUlsDkpHs2a+3VTHp6CTYk9OhxQUwgb1xfhU8p6/5w76EtAbM2Vd4KZG/gmOUP5Hh0C8
Xgizntr/oq86FeBxm2MqdtxTfXGX6AOfzGUHyLiDYQLqUKJl5LwiOvXjwvyoJofkcqbwQwzP7ZbZ
Mn+cK/v6cyeZeMQJT+aAp9wZ48sSzvdf+gNTcaTKOHR607WQphoVMCBEmDVtMo9cyOFtJpn8etyA
g5zWv2/vjyUDHSgdMcV4QyUgX+fMY5y2JyK/4WNIyEmi0pVSY6BnGurfY0i+Kn2N2NbEtHJokj9V
26fQ8h4Ia56dm268lxOL60192cynAFbWALkwmJ744oaOHmNvgZyIQbYwPLPe8jU/+J6YEomijzkg
KH+5b+apUQrBPrmk8zo51NntcM8rWgMv6KGyYS2sEbD5QfwfEv7qL08jqMayxUesyFuXyJtDoyq7
N+vDo/rJ3RlELQrKWkMNaCypfs+/IGVA9zMB15oiDZTlUNRej1vxxiqSwXElbDmg1/9Zt1Q/eeyo
QCvebVaf9zrZGVR0PmcGdUPLSs4cfMiEyQGky64SChKBI+hB5dD7UWSk3pbVciVhmPM0p680kxO4
xXS5r7QWT072TPkE0HBhc++orIIaaaKA2frMUjpPmwtTe2uA7tM48Kg2D1fjwONGzyLX3CYfEE1f
rqZ/k9B+qbphD+scaSwPi00701INwPe03jRbABnGII1np2sBKEj9EWlJ6fc+UurktQa0leo/lbr7
Q7PfRmujbD+02IXgbgB5FJAbMUddWEd/3hWMtzP94VL+UC4dRAaNF/ij9XB0CUXk6PpotJt2Va+L
SdSDcQo3zob2+QXnQb9BxdMzJbWseKY/fD46WMw0Ac/VXrvBdqVueEjkVf1QdIY9wtQWT4PU3wfC
WnW2AL5mF9/Qw6kkGUZIT1VCE3WuwygcZZdqRSG9tLdFa5vLKFoOXXOPCSqkMB/0lNNNJg74dQde
YBvY3RsOVv3L4QI/hvJZHmxxaFKuBzkHT24oi3JyuekBtZaUbu6vBhZzTh40hdVWLes8rcT913o+
AgCzmfYVdGq56lDFEtnPKOIbzwS9eF9qBRMqpUpZo8krCZtgAsHsSB+AmcMipeBkGbF50BU8cBqd
OJ6wOlGZ5Chi1TJc5vHTVoi6UrJhLZoXAGKe0mkMY/L1xezP1ed7vqLKuldqD0c0O3C0eHmQ1n2k
cX6MiIPnhlQv0LQayNQ6lqPixM3zPyeffjAR6KAhdLGC9sMo98TzmkwNGni2PqPywoZZEAnXq7ed
fCxE34ThW0gDhvZX9JvLRwkIIsyTPoqdR94+4wm5GjsJvGYr3cqAiKS+Y9un7Ijsy8wvKHEH8lFL
Xq6cgjbkhGG/eHsRnnR1Bvb4vRwSU6CaDapMC0oAct9mN+E6K+zCIO6z8B4H+FS1bpZGCsPJHIlM
3bT0drTok+GjDxTLC59y1WSvqG5+l7ST1s0GVQjnjtK2sRk2JRMQ9BYrVV/wK+zlkakZElpc8HNH
oAAKK1v4VDs960dn2PIOZ7mJGKeh3VxeB+bTa9KqV0kx1PsTqr9ehcBU8ubfGfG5RDTAoCi+kc7W
OX6PQVQHDUWVkwqBLWb6elooiEPTiD68g6uoid4D6tAU5tsE2uUTz313g0yVAkZg/ClwtXQfsr6p
SSxQQWQJ+zgjUwqAZE6u0/hjEX72cAw1U2C9mbqjZyiujBSRGonsl3cXmPUg1NOx880t2vAaJ468
r3gM+t2MtlsNR8sVkcW4LvLJhneg9g8CehLfpdPhN0Lk52r9jWbcWNOpXbasZ1+ZwxNZMRT+nSpc
8fSs+d9GJ/JmdKr7l19bGLNVF1mcYsm02oji1Z+b/F0c49ijvQWxuzwIiRkd1esDkHEKhOV+IgsL
WhdUAkgH5ABRD3/OJ2Ad+ci5zprHwR5JIkvWKNtYWvUrNL/nCqHfm4s21LQuUUaZM5TLSjegYEee
dts8HtQTPNdAukiEG0iTYa9uqIpOM5Van1uEXmVADAkOLe1PnDrBZ/sOQUjxU/J4cLX1fyskKi5F
9xQz6Eh66BsXbWuy3x2kiO8KtbBFKC7cZ/f+w0iQ/f+AUJLbke/cDHwtdIur/NiOdYw3+i3yVguZ
xeAaDBLmXWTmS9LHoBvuaTUsQ3IQyoyXNHNEjmHN3uTlRpS+771WtLt7TiNHyxZ80It29tETjBPU
+ge36eo+dMItG7JWXoLo19H5ILXBpLt4bySlaiNieCBITUbPcVVO6rdE6Fbik5/UpojoBLjhooWO
tN2hjpyTkeMvQ2bwTiZCVEsGcZ7ALh5YXhPadNbNwm+4pbQqwhVrd5WNrwTKy4giefDUpnOB61ZA
V4eh8ZlYZ5xjgKWDNPUBLU/7Y/JxhdKNyCj5i7dRMZPFmHH0VDkCEagvLxD9Q04NYaVHzJ25kjRg
AEQsWRpP8qA0w0Qv/O/fh4Ri1i/oqgd/E9VKwznJF6emEaNMZAEFWLgIpq+FAFCV0QDDG+HORhvF
/NU2sHniKkKvQ9lvs9prV3fD4H5Rjol26WgDwnjtkVSnKUPFnYuPVXtPgmtw2SvPjvDodHzx/ovm
CYD5aFct4ByZH+SfJJK3ErVKMoIXXcRRUG0J6dMvajNJiVaM8ciq9OuFXuN/KfXlzXAPhjOBsKK5
Lemcf1BOTI8nkLPgQUb9LVisrhviVneDjllXvrl6QJrTgHPlu+ChmMcrX0S6Yu+8QzFF0Ww0qtW6
muyEUFtRN2dTmEC6xVU97MnxqDI+PqSLRzTxzSlkiofPLp0+vi0BkbM0DWv2788Sczq359cJvRSb
1/EGoHEULjQbKfUbAVkp/EYbYEci6xolwCEolUz5HXr25Ft1trXhI30h105fnkJUlV+bXvX3nJZQ
FGssiNU6Wdi1Nuh5WZVCT2vg5jao2am7u24yUnEHHwEW5gtP76m2wjeqIUSTOr9r24eTnPpjsBbQ
ukyNXS7uNkcKEYZGEmPIZmLLW98ZX/Sz3nYLVwrQ/vzFqoOJhvDrNFajQx+XZAptgsg3wIDtwZjJ
KuM+rJ1HHhVp/SaJGs+uluhoPMdm+H9j+EPkQxiMoF1lBvsyLAqPf2kMFONcK3NXtM138UYh/tBC
m8WzqForntQL5zit3/PC/XMr7J6yTQ9qUjA/mGzhi4321ynu4/JbrecY2JlGwyhqkpuu32D3LFJE
6+qSCqI0m4/wQlOtCzPF7oSTRf0bNnbCAGKUBU9lypXjmG87kvV2Wa+S1tdNLXCjveUu/neXBLK3
D/+BwvcG9ZSWhz07cssffjKGMWMJTIL1VnEHFjrYRuOTzagxZ3rRLZUSXtJyDR4gkQ4nmh9ZtftE
rw3axaXu+UsJpt6IFYFIdl/XkcU3Z83k4zuNgtWPBPBILIt/LvtiZ09B2+KXZhNqNaoTWXIa/2C5
K3SI+oGKLyFF3FS1PA0drGcWCfqHQOCn6qm8PN4fE+Oa/Kft/KyBmOAO4MwQWk/QVy1Kg6Y7ui8K
iq1N9sVWchAvjyAqdE3JSSE9Djd029EkdmB6vAIWVdFnr3N/bb3+vrjspEDSujiNyR7F+2WH8+Qp
r53N5qFxQXFplZwFS8+/9DJtEWIPjWrIlLfdZ4/MxuV3oNSlgseXG/F3Oc+P5ysUCpuu06GNESml
dqE5DxYBD6+XbqfP/M/Y3L6WVDtT1SCozVYnPQgg15Bt+JfHcr4EI7wISSRmNK5I+ZwGnuMAP+v0
fzgiFqLaeP2daftfaeouIDANTGPlSfpoIUNTizzBtTgAIn6AOtyufOuQTbDSSSmnG29BypVVdWjn
g8TiXCeoZlVcaqy+nVZyaImHHL1xcSjX7pnZqJtgOT4VOe2FpTvPsXneUnGPBZZMwJb0EZ/q/nHh
NkKL8UZIc3aRcKxYnOVaX0G/hFrDIM3OGHvYjlgS+Amx2O4TNWlgdQH3FfjZqRErWL9kMBZTJoMN
DnChEMOgIgdCNmyQKYB9zWQAR0AZhmR+JG9sQPsQC3EPvylbGx5ZyAqz5zULkAgo/AO+J/iNr4so
pO2sCJEHYaCGJPcuTV3Sz5+UCGxX8wPYtTHjogcYyIDfItmAYxBFrTGzjbYkF67OnH40WLSwPGGc
93C2ajXNk3yHonPuxS7yRDKw1MUmwLRkfulrBoTOaWkYK8JS5gD29Y8MjLi02mG6fTdCNg3ylJTT
/zQERDStNqbKsVq3luCtyGep6D7/RsB6PXQisEqp7YPtm0LTaLzi/mXABmM+nR+oz13BnzsnC/EE
en9R/mjm/1AdADIfeiceoOzV9kVTq9KOSWZ3Tg+yLvnMgBi11VKbFlv+azC7vbVCn4TnAaKPiB1E
o5ly5neDLjXfhEGzQ0aAPllK8eFDG5Bi0fkVv5qPAyQzsn3kFA07i3w/1xEOwitLx46zfaDxM8Lr
9NZd3DYdtF0907O/ccB+fkbkgqFWU93/WQ1qkJPdDqSyzjQjtRjwcszd8P+ot3pKoKJMPb6FRF3s
v4xPHD+kvHXC9BF2C7jKFA6aO3MYthe1ISAuKsHZ4eSq6mm3HOPVt4dyl57IQV5S1xNJSSNaK7mH
T5N7bXAN0Zvtf4Cb/wRrRiCPWiiUFd3dwk8ez4MFogvGlH3YLP1+40otTmbPun2UzOdj7GG7o4it
guxYM+NY+xHMt2leoM23Ggk4nIyfbXp9Cfq7q2D5TRSVwcx02gX9efIL86u181l4m50PEZeT8DZC
3YQWkh1drHsx4hZDYVrEJyeEpdhZpyeF2dYTDpr3SiiMdF7MYeqFPN9upLmbYnE8Bv/qnZhBDr4B
SEDYD/zdnmi857iaKKHb/DENjugsITk4vYhEf+r5Vo75flGaFgVI0swCeYY5TN58Ut05ZxLTUhAa
HqEjaaty57yAc1dTvsnEVOKAUj/MofhfsG7I3bExP1QIc4VUVTlO1Ujur645ONazscoA+ceGMyNo
erx6jEkh/FgYkA5abIovoduGBXTGZ7/nMU8TvIOv3LADyVAKBuBgnUrg4ZvUPsNMHLc9gAPz3u9o
UJYe3Ap876uMnr3aGsNs6ywixR1Qh9pu7CaDYA1gIMX9/upCuviDpZsYxVFyBfGtDsEXJT4nx1P1
rspM9sMqHvphKUaZpTE1dvwSqUa7xjZdYaUhcvjNnHZrfuosA0XtHQE51k8ZP7RgRaHWcHzGCfYM
h80WKXRQfSXxbk4UGbkcaD2V6axTQ9YgnEPZNm7N9G436cHVqBIpKLQc03WS1qRC2SLuuNe54LvB
8zeMrYEpgJlJlexB2q+luBK7O12nog5R4hMIXax5qFkO8rM6DSZPqPvO4nKc92YqSXO+4yyEMvVZ
DvRcSx4G7UGFg0o1dor8jHwlw9MEdJaMwcb6SSBR2gbqaN78iabD7q+rHZE8Dp5NmCPF7qodb+vw
fa3qNd4mBRqExpkDyv2cNcd9W4FsZjVhSBy1rZi5HBRSHaCEJj5XBPLfYyDlGawhsij9/OqlXQRY
zKne5yS/ZkKocOtk3f6dZ6kKa0vvxV7WudeIQK+GWzJ3Au+8OLGX2la1m5+dQWQ2M66zPn5n1Rnk
qrGoxlTsAV078DvVM33jIeQXQywCngioKZEP0HZ+WxwKMRFDDI+96XsLv5YfhjDxQ0ex5oHLkRkp
x7ssS60tcXwuPyp1fKRFC4a3f77XImHFneE7ZT1qLcuvGH1UnSGEjSKXsvBQDFx6Iyu8O6F6+yEY
ybjib08wy+BIvfm2pI+pCtyGhPTUPj8hFYXU0y9d9VK/fyvI4GS1dIlPljmQ0OprX4N2fW8edv9O
AReQ8IPBeE8q7hRAR8wEJ72SYxpmrLbDVVe8G+tc9b52CxiXvegdfATickBXzBGtFA7crz6LQRan
DL2me1EXDqre/Ws+Dbq1X4p/78hUCdqyX9BqGpG9W/DoLB5AT2sTs5dsnCTB0n8y8v8cn347Ljmq
ahLL075kCfBaoAJNVZPCz1614qGp491hx7lHaveRlg41+2WBoy65JQEAKecabrr2drMIOSnqO2BQ
Qz7HCN+oTAhrKUsCqWDtg6lSIL4CCOpwLPwlmnmlW/pfWiY5Rh23fCg4J2FGqgIQH35M2/HWYHFj
yUe7PgKhLq7oPwQKZClb8wN76Fb542TJ8+o3zVBH21A7Qye3HCLD1akFsTKOz3LRcSsZRcIG7IXy
Z9U36mSHbC/fo+wgyhsdXFKck5QdW1JcmHUMaXHwE0aTnth2VRlN2bHniFmVns90JNf6DTteSvNL
MqeM6zox8dQKlpRjzzey0jkgdLpvdHuGxxJMwOYsH87CKF+pVNSZTbZNK7DDJC8ISjrR60XidgON
kMv1mF7sUG55bhkYWBM6KuBWtFlvfw27tKoFi5H0tdKtnKQVw6U3I4baYU1fh6KMoiwwMfUBFsQW
qtnA5MpQ0XfrgZ9xeCENMGulw+opMyfX6qC9oO34yKda16HCK+BbnYfsCfQ3pYu5Y4oFvNzY1RNS
ZtiY8XelofIZW9MQFaMi10TzwTTAQttIRuIdyhTU04Be/x4Isa5cunpJ2RJspbDBs+rlcWioV20M
sSEE5pbeYofUo4P6t1NeTVwoxY470C6aDwbhZXTpCQKPAbFsM6BppIaePfTA7u87ORDGeRkpguqi
qSqCFjlFj65VHeMX4C4mr1Xofb+dbSIQMRQJg6MjRbo4K+prBewyb6szuJmpg81M+VMpogg/rcKN
P0zGz4rUwCQKdRriRIIxa0xocJa+HXeEEZgjsg2a758PaPrm6R7hSzDLINXlD3uobSWX9hWbZQsD
UPQU1sBmj6aoXBe3v0iZ/F4JjCXP1cfYe2Bb7L79fKfMdxNRbsNZfO5DcQ/3qP7Nu7EDpo+XBSG1
7cNC528gwA7UXpVJI3gk4UqyR/pg73EZD7+YFjxExhw5HgKXb68aZhh9P6ivCob89TduzFW3keL7
4dwx8LCcVYE9ea55Vq3BHn27qTIZs/JtDjnrj2YIHfcXwOeSNCaZoS7E4K4bzU4r731zdcMkq3qe
VU0qQgexh6xgm4EEFhuwIPDsSKOqvgiph4AfENTvWRGJ5F9RVlcKDO6VdYjHTY9FQdm+ZkRuh5NT
ZBAPFn6RJ2+ZN9N46vLJbeCpid5QptDqO6V1z7EzTQjmc3lqzLYuLkQKqzdZNeukBXk5eXPDMlL2
3mXZN7QemM2HSmPZhK278EmNpvsyjIFl1G/q+lsCDGLtEvAzEFgUV4rZq/067M3XigignuHJp5hd
aCTYBezB0RLwkS5uKOKO1hDR9CU6TYOBwSJq9f3rNUq+XMPu28Us7dL7mUXnyvjj5QlrHeWoWm9f
UREpdgsti2/4HYjsJVd7EYS4bvq2f7fJgZDpgJ3TRwZNXPuPrdirTiUE3z88vdOY6doT2tqvFmxy
pClu2BjJrQMzQBwPUcBRT0kWRJ4lHwZy+S/RtlzwGmjiF/LFhzrmxzLyh23Nuc61VdL/uAFBr/VA
BaXjgrI+4vzjUZ50pbVu5T1DBSg5bgETHL7fSFHwQ2v8kBWgQP/B1dryvwW88F+nwNv4RI8Z+tjY
XmSmXGpHtduLk74CjgpWqF+rnNZa2tSSGcdiFCk5rwLcD7tJO0IvVlI+jkxXNxsfYrK8Ur/IESR2
eYMqTnMVwOh16sFsYa4xe81oWLHMVisi7fnheBr2n6OhDnA9NZzIKpv6LrtOYn5+0lHrRjucMIUi
CPcb16TtGPx22sH95MxmE5eeLCwjtWWkHCWf4cy395eP07iIkQ6bIbIPleGyPfYXaJ43AiygACO8
Ag7g59hm76cxYVJ7XRWeIzr3UrAfVjL2j/QqOAVjfbFAuXNxy+dGL8PL/tVjNW8gTJTQHjFotBIw
sMqQ/5eMnw5eOvNSeE1r8RRvlhdcC/ViKMP6D6nkcR6XKrAYxVrxdmBdj1lgn+R2x2vcvHRQNzOq
llJk/7YjJHd9g28pn3eJctGifT2xFS4zz7pTu45awDGtskc0Q3sWVyrXypQpPWtaafUVpNHidX4i
AqWRgAhlXjyk5lHIaX3dm/JL/iBxq5yZpO+OXhg4FU3QPM3KPjhi9Yxp9DFU5agUgb9PfYaO8sMK
Nt3p3alkmlWf5IRAROnoJd+YqDDGE4dlFKs9U2NgeWsU7u3+mt9XRR/vEVzGEwdZ6jauSod0VDcW
k5LhzuWlUd8b5T4RAkaZtXFtqAHu59ktiXzEVtmE957knzPvLKKDTNDizZoDD5aB4cseTHIUnMs0
yhCv+KgjyZaxhh0hec9iw6p/QLUUyonCbJcBVqN95O7lhcvz3kMZfjIuNm+C05quY4VuC/+cXhp/
qLTAIegTX6+iEr9pfG9q0AlZ+sK7DzphtNmf65lZLDH5duPFk7mayhChWk5nIVzIJPMUIhn1vGOi
zU1+Lmo/I1l5qGNvrnV/SjT0+s7Iwjq0W42tLbYJwUVUGJF/I7PeXTAeOaAqUXGGCvCO4GcONXj8
TWVY0hP+2IGxaL94kxuWe53VZCw8zRYvhhDiGncfATzZFJQwtGk4pWdXBv/7vhuTHZsGhGWk0kxb
JCI+jpKEGeWa+lbmFXowyn/GYg7RpyCfCxljPU9eOk/SB4d9i3YTYiXLN0qMhFuy402WXgko0A5L
ZB4L1PGLeJbxXCZGVCqdQrYw8x8NQ609kKG4TkwUyCW0CYWlNqfyP2b0ZoENlcobSPGcLqRn1bJB
zbZJzP1ACh7uxpWoKuatTqHY8jywKo+N4r/wBwk92xR2PuIu/W13FEUv/1eHIgBmePFoSIoS5pxo
nwaHdJTb8ndjQaQqVqSk/lDWvmyGr+DO06AS3DM238VG3Hq+Lo+wEXyYMGrvowMvVRO/8N0PRtlc
cFefkAjLENUqIAHcycBnTe5g/ZT2ZNiKEGceio2siKcG1jFbMgDdXgn4CRQcSdAd/7zu4y7v8YBw
mCcgB8ZLBOco1QlrlPL3PyIP7qGfLR4fmhzC959e5rCCAyrREx8KgxF+IzJlAI3HmRObhjURCrQy
1lFB97ihavvpKNeQnI7djpTuUhB/v1B5QfAIUMhLxmh4modqJG5pT+3Jr9RD0IfEzMf/ZJISVufW
NKfPQVGdhnOJKkY8JQ5xhbWLiE4XXjh7SC6bWGIBUJkkAqRhpvhnMIKCyegpOIJQPwj+JHX2rC21
NG7InTl71w52UUM8k6kl7SGK9rqZagxLZtyrAF9c65Gr3BlKy1aykOP18FPyx52zbxWX+kyaJgbJ
qMqlsy753npfFN/VTyTKWAyIWfLp44f7tbeIAjRWV4ojEN8UBxy100cwaSBp9I+oX3TyUd8pPP3u
j3moOl21v4KoP/ETTYlkc3eB+cpP2JJIeqvkyutedFCZZPLCO3VFHiewpe7+sBOfU0MaGGp5Mtse
sVJF4aEBztR549Djj/LxJneXK+EMV4ve7A6CWsRJpXzWZ7xT0jjMfPobpel3LN+1Eyz1x4rO7pfT
yD0qiPu8UP/9kwDY9JxDHKDJXrFzEBLIUQHFv6py4VvuH9UZFEcz5f36NCGBDSR/m5iaEz5xMol7
UnLC/CMTo0Egf8lcwpluxr88eUwwLe9O78l/Cm1+kUp7HShD7jKXQCh1VtI3SOQYoH70RSRxktvE
ruL2v70npAk3HYBkJE2FA46poRGqlsWWXFyGDjVkpx4ysVjdd19wrIjPH+wYHfuVNqbnkETB4CpR
L74nD30TpYCtB9nJPUMcS1YLO8nxKiYuXx2pP96ppET0/pISQsnXiMZITqCyzeXL7rvTM3MdDsZf
jwyYj/55bFCh4gWDK6t7SNOdJk+bk8Ix0TpQCeR6N+RxaioJyfGpEgfRs+NZfO1ktuQano1bzsZc
/yaJW89BOFrZzG6DRmpVBIT3wf9VMTOBUUduP8rE3h595+rUwtDLefeQjpndgMOaOTDBrDIMuYHK
2DZq4jBSDtN20nD9lIV6uSt/AmdghnVArGq5PdRMXwpHIVnSis8eW8YXWn3mf52LUjzJN85BPPtn
BKWDHA57ZFyC/DfZ5q6g/g4msyfmvHviBqyY4dGBJSNc+h3KfHF+zIEQNJ6llmT8hqqkGQgF63P6
rKqMsDDF3b9YPumgHgsto5Z80vUlVNDvg/vj1W4bSjdNVgAX2f/C/Omb6uiD0TPkzvJqLiEFT6lH
cqa8U00CZxcl6aUKIvMCaz1IlmxMcpqUgD6Kb+YWKE6rKAJF5KbHN0wJWAFTIBnggMlIjZm0Z7jO
Ljy/8SQS7V5LHmId78vhLohlARd06mXDJk+3Tz+gSJ73SFByjjKRFJInUiwUSoGgt1sqHM7xLY/P
6/J6e4QbT7dmMK7iy08oiWIiKmGKtI/Vsq8OPgQTfYNLc7phfRp7mQKwZdIn1FNzuGGPkAF7O7Lj
U3O+fr+sGL3VBkL+WDL+eUPJs+u+QG5aTViG7b0VveFY0P6CQwk6uI8WepKvDjr8RdkEn6kQBHPO
HIF3D/T+3y82aNDROyvWVjCkkX90OQPERdgcjTUetEuRgOyegOfj9AUOOIXE2aZQUkwjLetnIKV0
EW82sunqK/BGcnN152N6RmIiH3kON3TiFBuCIPPHgaKMOMAGiGHMiUMCS6AQo716l0Uv91asrs9c
bBdhczQDYWRXGWxwtpH1HCf3HeB47GSs7e00tYRTSzew6BEe10fb+ysX2om6Kd0F7N9lDe3zsQ2k
gnS4wvID8j7puxZ4WpDPVl2gAHhT7hzjek7yXD/84VXXttVi0b6nKDvZiPrU3wW8xUqTH6mqZhNF
S1l1MWQChqD5hN03AdfE6BUnpne+nbZbCgaRQdyeDO4fFPZeXoCnR19t5LOFpah70Gfj+WeCJ087
QZydEiYiZMxal1czIcoKwb03+/0cnbDGABAXArGCmVMrOHBEk5dQkLlsZlZ0ZOChF1Q/kXQAwMYB
N6jafRrw0g1i6tCqW8wTj9uddUFKzEadZaC3wUWXnU3nwWsJUOkU5/d0JJ2fZ6vJbudPXIZSzYuW
mJxayDtoBCFWlSiIv4eCh4ZGZlsJtcTVw+GSCzkpgjOFHAmSdKerh5RMzX3k0EFCR0K3rGu+C8LF
V8yXpNLQ72lxWYDl0Mq0PdzKrw4D0Myv9/2QHxZZU+KFa/FjCxDBnPFHyaVd3NSSkN12ySX13Wsl
9vBbk3l7BVq/UG3XVcwZdhNPgjmXXG8VGwDiBc5NW2o6GOpriWFwuG/hncjibFds24oDc+wWbBlf
Fv8G4l4N2ghar6KtaM/GpCCjfp0RMamUuX8Oc4cCe5h7ExsrhcaL/UDo9ifvgOuMOS+vt5aUPjpw
tFZQ8FqoiPhj5NfnJo22of8tMBHG8RyX3vd2PVVXHVW8maqMpWUUsFbcfUb3zZ2PLSBJ4Eb7vHtb
9LdwMIXfnXE3Q2GR4ZNaYb0plu1qALB8n8CUAFol9CTbDi+B9aenodKmJul2atoTqE6OZVNbem9f
WfJr21hpszEFw1P7PNB/wpfJ66gp7cfsvYHQRtupnzOWJJmxIikeCVWIJBH0StQWatOPk1oHJomV
TCwvB+DTcVHCKMVfkTU033ZFVfWD0f7cI4N/4DXVyhD6DrwoJrKM/FeH71+OrjrF6sy+fuPPFo5Z
iDmKtdIuSdBoCcztMIEQR3Eozb0dp5M+Jf1fisgRKYSfikFNbCm+WPlwcnpHrV5pbUgohAZBpQye
R2LyKELBpPHfekYIXZ8/6L/Ds3eXhRXuWhpqoJzwwH679rOhNVkJWsmLheQCIN6/Kp5rDYPGQF0r
CnO8OiXLTro7f7ZaX4Zzg+F+HBgwr2AFYIV7b5uPMDhT/o+5KqbE5RJe+A+GbT1yio3NjxqfS9dv
cLNiB635G+cAMrzRssbKG0730rqkuacBQdaEhWw0A0VNvuV4ZSX418tx6J9An5NPwUct6mTpLXWx
3uDpUJxZA59q2M8heOoUX/i0TTZ13jKwLz4mYMbYJgFqTcMakMPCkfoEJCQ7cIvb966rXEvwWhHQ
UClctd5GwmcsMvUTgEtm4+U+XhuZXzRGDe/xP4isK4sitFbsoCAr3tyVOoAtbsqbvvbg09W8A73M
WtKtEx0HfHsfRVg2v/iFdMIez0WxeWKVprddujWaXSIQ4TEw9vKu3oWX6wzInstul/Gl9ABB8cyM
69NleTFvArz5jby3tGF3qfXWrwuviWtuYbzbfAUpaj9AZCJbO+pTPhPl75Ak7PlvkdWYyhlInwkA
r83iEl+tWzPchlqt/kA1f/QTm1Sv3nWn9JcKXYZuLM3X68mowHb4O5Xo7sTNaMkusY6h834xK4uZ
Of6ObweqZwEho0QsBiTKSReowoHl+150tkdz2HVqG45KqyYH5gXStyqBhoKq5HTeaCM5MWjo/HZG
DtWR4soeX1tshAL4nFMaYsbLq9prHVFOKpVWj+EQCfwJHd2btjA6gp+F7C78Fj1ilRoohepX2AZi
hfIzETmNhJ5QlyDD5/WqLqhVmp0spKyVw4s/LEaClKUo60WCOzUALH5lFXIJsBqjCffG+iosSqfh
0A/E2irVxTOLp4G8ewdjp5OO2Kh2dki68jj3U0ztiGTLVtIOBKRumYn/1pA2bd2Oyi3HenwsIEdm
l0QKnFA1OZtzV37h5v07FpbF/dXpY6V35XxEa3pFHc0ZQvXwnUMQ688oJ0HZs+5XAVSYCXOUsVcL
N9fVVsBPMy22gRYCsZbkvdNemyalNHlhgWzwqPyVtH0Y/pVgRRJ/0GZPYSvyDHGEkdOvguiWnHE2
i1rFNZI8ANluNMkqWxBqrJHfW11EtrwM8PKr54TZg8w2n8esnHKlSlP4RWJzYzfxxoVUV/DMfLs5
tVCdOtsWYgCUWNiBac9cSXwSMf3lvPvmOz7HT2gjckDb+/YmwbSbN8Ht75OkU3qKe3iUOEwOGjX4
cgo+KUwNTI+Q18GI5hzCojzy+cS1zOERRKmx0zuVw0bv4dZctN93KjmZiOK9saeds33Mvjt5oId8
oipyZL+FRMByC3krD6WJ/ARYGfZktb0xCwlrSOI6J6GImljhmsgT/ss60X2ZSX+eFjxjvYSnQm1D
IuzpSs9dvUkb5c/l/4w9UvcX8boX3vLLDMc889DL0lou0f7MqakrkoVmsSOe5ermH9/BQOHjV1DZ
3EVyVXZt/7Ez9WLSQJbgMX+Huy4uEu/RpGWhqKJO8PQk8LBitwEUmP5XVcLwPJOV51mLVajxeCVh
JmekjK0WMH3qzowB5zUO0NQVOJuCaR5r0cP5mwSE3vrud4BrlYI9L24rh0hT0wUIi/12ICxttRB8
gtRgbRo0VRsUnbYF7TlwJ5BFEoJblgeX4raC2LHHIL5JcToz6EJHvYFDXzyCoqr83mk3PO9ubMYu
AbHvGelOWRUpdF5dPDtelMkhshGjdNJcxIf+3SX8GyD1Ni/T9+bnXOGzYkijKZyEEogaO9YMKRXn
lFhR0Z05zL75ovSRFW0DAiZY+mEMJXY7Mso13esyZebSonsgMHV+gDRSBnAgbEQDlJ4gc0UdTz5H
6yYxiZGIxa9J+Qf3Km9jPrM1qDlwsTuFvQ6ATm/OQPxXJJH0AsfHiA6385OVBY2a28yYK5nBZemW
YbUIVmfZ/CvXD43mEOrLpqcZa9ejNSVnmfbVwGljm2/CWVBkx2urqXYG/nnUn2++O6KSf0QIsyLW
87E+rGUpvTqBAEUyORo8HzLv/WlHRGxHGZmX9CF3ZQ+t1WafDbEEW65K+2gS9EggSyVVHECgAMpm
TMNBA9ftggbod6LDoMrffucGwxS8QnXa64p+mnxwDN/jqDoFS+E7Bitt2XKRuFhfv6YwXAvsBeSp
KHr8myLt5UOC41JFhKO2Zyl8Z1PSLEDvoHN4dhc0E5AYCEiQlAqsB0qq5HIhZoPiwLjeTG9yr81e
dy13PjrsoAdUnAU+Unr7rCTORUTajKlUC2ys2pDnM5IXyUKk2q4DntoXClg8GUubI2QZMoYQZ1xH
JelUDGFJrz7ffysHGuBnGs216PZrynZV2b8Io4aEZqUyen95WtMrhUTKBqUPDAR0jfwMoWQ1x2Nm
l+UZZnXzhd3i9dlWPU/LUhWFn5zcO75JFqPew9FRs9KCmO7xuR6WKojhmfdUqqkKBmfotkazWrsH
qzsi+V6bzeU//rhkQy3oQ/Eejy3BvS2vnOXwhRIiTLpyK9fM6PC3DRZzzMcfKkeepwYq4KIm/cUT
MOvQHPdB7DISFi1gNob2lOAItH+dkWBgNNZT3N3ERPBnEFtMTrtNLHf3sikFda2EmFw87yEve8eh
2OLqU4LO7DGgnnRInXPBapD8EO58VWrfhOgz7VVItoNt09T5A4JzI3vmosizzd1OPdZ6ESZJbpbN
vscPbfWLAQbahmA5KhA/cLEaGy+wJ8kANtivt4uNnVIj5HFEzq2QbMSavF40vW2bkNCpvf69+fFA
fPywn+f16Bp6b1HDRDyUcO6Us7ek7IQAkhg9dSeXTlf+ouUQ6W39ImmPqdAoy1fs+gancS/GBQ/Q
rfIXEGuWP9ePaEr73q6zQ8sbWIZvHTRGVps0bWg8C175p0cv2a9989l93tgiqclZuI0bgEOYBAFq
jjJKKxbY9KaKM0k81O54TQWBh2LTrfTZvtr8sgJQuFG1s7wPo91iem1oqjvHicyWkPrlDkOwU3a+
J7EV82ErU+92kRPf/ClmWja5W3ed44zt/msJsI6fyUfHCtOeUOQs+R/rPkbVGhkNcoSwtGn1soIC
xzfEQNmdPJjO8VPgubsZU0/3goJdhMMbLSgxeTeHH/sIjC0+3ricyiaIcKRLAf7ROvNvEbueFffs
a8VdviHaLfe6RhOYJi6hHZlJT4ZHNRs95yX90ZBnJCFf1X3dhmGNJKv8X9ItLwcfHcxx+UUWYEHB
J6wBzyTIhI7MqGpjfmAjZKh0Dru6wPPpBcVB8O/2TS1ZT2/1Mh8ThrmeK/MJUc64gnNbXHK5zvqM
apuBJ4rwnvvFTXouGdLLcX6DPFpFfTBkzoIbnD9r7O8cYgSMR7I7MeRIl+TbiIPPFNiZwOogGZ96
qXltJo9ApKlhacwGmSPHpYMZsl7Z076uHWY9lISmYRKnLIFrpDBsKvnVmuZUPDzID5Fp/Ieahuvd
Elor7+wyhtsqFD9YxrP0xdzMWvddCqxeTpS4svPKshHcqWOBzTL9UDWEwc60foBFAIWQtpQdLsYP
OA7ZF36D7zw57jZrI15Y3MSSiOXgviA8FKfv2VhA/YlfsENkDJ/ZUDESOGDWtiT+pYrX7MRc+0+y
kj+8iFPhhv4NxCaldIQJ0GiPSp02Q88EZGXARZsQu2Nu0Z87OFTuzhw9g41IOifXMF8Prp0Tn27h
Jl/mstJmrhK2l8ZiYqPbRgnlvyGN+V5XePCBPi8DAEwD3skAWh/xNHoqSM3uxssJalZdUdvjotM4
t83/s2kBBbtfkXdt7i4cPefEIffRzsvpIrXYNNfREcwE5BjXzoxr2DQgH81G7oZ5u2O2+gjy4pXU
lV/HIRk4RZeKS1jldQe6cBBEGQ1GycNouxRfiBR9uqZyZwO8It5b2SyZ6UaWSXoysdqi+L54nKTW
aE9VTRy/SC4sLrC7kf2Yh8nD44GfnPPvBeVDInL3QvsfjpEPs9Zbvz2QnLOzrRzFRpG/oUnbX8nb
8FcLkQ+REJKqm85638FCDy0VQBj641MJSrrHju5V6Nef08AP7naoQxzRqAFIy+wkyo+ePlPaV82B
9IXXdc6uyxc6H/7H549IjDVh6BeP+pysPPV2SVgrwDQ701Owi4c/XJJSQq99q+I0LPqcU8ZUQs/k
iUhUz8xjh6vY9QADVFX9YxnOdmvieipWAuHwTGRpXtKjDB3OQlajm/NVupyKzbzz/hwIovsgDCfG
qtRYkxyA/Vw9xkFdSIlNWph6mtoqzv7RC2CbEV9dsMqPlaGwbkWFeEX5zPeS+qYCY43ah/ar/srx
72Cj2HH90QAp3hjJTqycB2lOywP2YIEO9QJndR4+cE7Q1pETpinzBzYbjC5sXj42JUdp2vIYOLlS
x1YxxVaOnCmBsT/HMnVNhx//Ngq4yra9T5hnSLrmGIYUoXPZfSb0xDWxT5Rpj89buhBcEUFIDRi0
7ZGHu863D3M5GGunhwxAlgRxqlbPfOwTXBGkotyH6kkYnhyliVbBOpIoG65A/7p0r1ItSyTFl0Wl
XHLuywyi3RgJgi4aZcYYVtPLcwvdt74e575rnYNDlH0jMpvm5vIOTucgWOZWObS+Vb2SBBWmAU5N
UMk7F+ld65dUNTrvgXKg12WZ31GL2/8GG1auzDoMQqZaIpj5IhfZXU9bKOtjuoHzmj9pnIRbsSkG
+nTivnCqDqhrit1IKankEKoSoLO8YjLOyuDcms4rtZDGdL+jlWcirnl4YQEkjBZnzccqTtnJ7eBs
apfMYr2eDwQ1Vq64cRkVBY82cAyK2KUMcHtVnmJYnMvoZ3N3bv4NsfsIb2J54BcjKSd5ZD9EgVnl
4D0upvIJvBd0IvwentO8vypur3G5Q5Fj2r7W//pGMWVu6iFNYJvdarHEbn4zfeGwHCqLLZdyR/cm
kux2rv6sCtDMSZUiwB1VD3yKZ5/RbqSVIsVSPJGtERiWrvea96plFRV8+lWz6y+x78kFf4n/jOsM
pJwWfZS3a4ANKL0MLesXtG7/2pl8TKysVSyGhjcPbIkNDv1nPJ1G7NDmOqBF6C+nmqpOQErYTFLY
F7zLzDwoya8Dy1sEhNWB+DCygJ/0/biBT6Ey0hhMWQoMYVSkJA9+LS6faVRk06Yun0LjR86eCa3c
gJGmeSJNrwNQUn/U9Uuacwv6hCJn9shq5lNn3o+tgi2u0GyyPW+GI2BHJEzd+NW6M7IqYp7ij/Uf
CdQQgYINGv33yWJIbSMg5iLXz0YTJqGmaIfXsJkResFYq9BylceHrVbJufUTscGIyR5c2wUHzojH
tJTICRYQ8NUCVn2Qs+eqyN/bEsCFMFnGpe9RAg5sIClcNHi/VAUrMgHFX0GGC2O+0IdBcrERKqRG
9z8RdMlqT5CbbCE9BFCLZCQ0ew/+FkRdhXlWZNj0Gm7CVLAOrdIJzvBLvah6OKLvfKsJoMy9gvv9
SYFpbq2ljh5zUjrNON0+BTn0xBs4FhWiHf+ee1pqrB4kErwKSmqpVEs7GpPRJPuVkEo+VyeA/RGu
E/OncmgK02whLLze3VR3W8VWmrzEwyUm0B5Tk+tRZhfvZLsWhVYpn7R/SzKBvwo+LRndfrO/Vhfm
JuP5yf6nqCYRUI1AFbmJTSTvNmJK+TOe29o+VJCv0IW2HMFoy49P8QULabeGBTwLRhWGIfPnkCQm
MpSxj2SUr/Jr9xykxkIUNjDRuY115S0NKRLN5F5iiscX+UV4tUuK2h759EFMFOn9yS5orCSgOsIy
T0FNQzjLBFOoHKrFJ+CkR57eBNU/HyoSHQ2lN3Ht469wvPmafuRxfSh9/iZmTQsykelimnaLM8RS
6jtDV2OWN2BPluITskWsTgHu/wnR3YwcZukh+T0+PqIqPLmj95q4qxjlnedgisnPOo8cNRqiXlbB
zgMVCQoCXOVYGjsqc100oyuiYuMj8S7VrV0pEcSYtk+CbCaqzWTe9QKHlSRYAskmXVKth+fuOBoY
hXHEPkcHMxB1qZqel3lOheykY20NnQnxCsXrpnA1YdQhpg9UAH+xBmv+EG/q9vH8Bh4pKG8VU/eV
BXh/PAEuwyJ5N6z9jAcyWEQyOHgYpGMLOCl+tXZNt162bbgiEjDzParA5hsXL2AyZyvWvdALEhu9
Bu6ATBt1Sy3w/YlZCR5VOn9KW+mAqVt8oeN+Dh5Y0zuCyZhqJ3yA8plC0ALxDvnivQeQKWeC28+b
wOKiai1CEPeRhkJpXKmjmdxTpG8TWCZxI5F3ngmTf+GsOIWNdluM3o6WDcd7rVZZJkdIxIcNu48P
YTBvxADNYcS8mipcc5KLoqa9qdVNhrq50J0qDvkVq9ZUf5Z5BtOaHCO2ulVYgQruXZzlG5JFvt2z
vVSP5vp4V7sCY65RIKWL+cr5xcoh1gXhMJSo/NVhaatUbwyEJR3YTCfR4gopsPj9NhZ8cUogSS4Z
b9rhngNnX/UFPSilbXqRwbRptTdfnPqfU1ZN28tv8PvfdNLqgH/uoncCWPSZRVdbzzFTVpV8MVe+
R4hwhhXY8qhI+g5tBbvAPpsreyO+jRn3RroG3JQnGadoV6hAMsvgaLY0SK8mFX/UfGFDgMPKbUf8
0M3c2dA8w3pY/GFd+EW9AgbWC6H5JeJk8lKzIEr7BIVJj5ohftVGSg8g/ClfrnlwCdeMg/EAtbiF
lyfOkj8MgWaUwZpOKKXmohse7w8N2WKEjDSy2VJYkZ0ZiHVPkKpxJex+/dwXB8pN5Pwv8c9QD//O
uxgYGhA2+LnK29j7RDEhnh6+LjzW6iTCQBcootNw0HUI1DLsC452WcU7ZFHJbt7hgtWVlmWUCNwk
P1VaMJxHjKYTgxom39QpXrSFP3mJU17S3RTZd4WEcieba/I4Yzh4TnB+v/8JYbbDtstBdykjOU9J
NTM+TVDh2agnbGqyVdftwOExzL7M6YeXGCj04eLn/z+ZLZooaj5OYRr2AReUN82/jLA4vscbIWRM
55AC4+S2tf//oFjrzZjY9sYcLkuM1XK1m5U4+2lfTChvCecgaDu4cp6zfDf/ehYyrpYw8ysZGaZn
fc2FVj8OaSHDNqkEPGt4doge/iwogwVgAdiOHjbxp5TdhzC2H3GbO8xv19fk/wm4oNpS0wyq63YP
oSi+aXR0WJExKyoezhfWVMs2B/EKQfx1IpeHMjfGXA+vkFjQajW5zb24+NSubr50fxYB8vMsUkeH
puns0QPthCcUwpaoktBWBNes3rOYQ9vH1a2k143IHByopIXoCBe7icpAEVf9/eSdHH3CsbTMSCGn
QyS4U/IB4Wl8R9DrGOcD3BpFdQUQDYO5DOiEcBa9NnwglfJLj2W9w8GsCYxiSBdHqHd6wmmTmA58
A2UrZcMY5vCLTcFn6Iq6tKTqhIQyD3zm/A8gRCU7N3CLJHnn0uibpqXgabXwQxBkFBEVikSat7j0
XAdnbb/nbbGA6UtsMTn5ValpEsGiFkx2Y5ltAOfRwwfXSAjByQ0Ul4H3Bmz9gRjaVWPuQx48Dzn8
EQ69DwKtdQQczAe/yzytM00PIVjPQc2IXF70QIAcsrtTbuBqWd6m0IYV+srmMqMs8Pq2AgGylrfm
U62rXCEOdh9TGxv7JtAqxBJK++9Orfsdp1qMxMLEfWeBP3fk150KXI1yfPbMoFL6wLQT5MKXuqfP
RjufDy3QyC1kraR2GWL4EuhzUKAk7bI9mAU7e0ToszkqJ+pi19mZuV2R0jucKxHza6OM3SsBdoXp
Flj4YrOLOInDAlVPHZG8plPyO3C8XJN0Ckt4PfAo2yF7wmpRAMJ137qDDlwIWPCcg5DqC2qrsFHA
r8p0NHZ9jRPifPqME51JeC9xPsod0zq6mCZNKy2H345OE1ATpT/RCuIb3b4TinuD+yQzS4yUPexc
htFLdIwZlFoJN5Ik5INE05OyYA/KSQhJV5wU1M+XnOQvdTUXXsemtqxhPhLqbfUU6YMrBB0nJRkv
2o63qEH30rZiafbS6KpQzKPA8GImz0gRuR6iH/YBut1Y+ZnQVR98C23azcCJWLoG/JrsYMOmq2If
9AO40gfPG2e+sFlzY20WmyxtS3N1NIktozE7+grDwuZeFTOJdXuzrl6i9F3kH8HBSXSjBrwh7U5S
szxFsHncdblTorkh0oB9F5W7aweD51OlEjYYxdtzTOC3tfjLMwmLY09EnGhKOK5s/MnKPS/aCQjB
9hZDRWRIgyg0113vQS8agTjwnTHJObnkh1bm3vr45SqMopb2+RlFkPvKBTq/FXlGxKBC5z4SaHXS
axmDvzOrxbK6wEULz/OUFVljAGPlH58ZWO9NooHW2Ti+ajy1N7eYlwgPYBoMIgOuBmfzYO0cwC/j
D6I0vLSOkWV/Ffl/WP3wjZ8Yt8iCeNriJ7pJILvDLHpWRuRABone07njD5yE05tuljnAmP3kaCek
Bob6N+lxdTdAuuBrRVQx39dRItk6uVjRXMmfo9mc2KcgeJuUDMQM/mItSF4oHVsOF99fTBu8xUdk
m3DCQpOrd43MdY01RisgBAHIo1xpat94X7vxaWr9sUNFyVg033R5xcirbH9O09e4UpUSsUyvDXlT
9SMaJhjAXyOLFrmW5utLZzKFGKSqYyD7GLeGFbDc/F2IFKGIG9hJXRmGn1w14T6EZpfwxirQ5LcK
xAUO9JSP0cubYXQ9w9j8ASbyuO5zhv8R/z5i98x6R2eRZI/GEK8IGE1D8xPAvsqOx5jjN6n+uBEZ
1RYyS/LzTTAYEjZmJfl5GWZ4TUlO/EEnZfNGtSOO+KFWesVhidiczXry1f2avhqSDuqG6Heuuk6g
ZtV5HAXoNwUG7sih084Lou3PHhdMYxsgs+vpJHgMnjy7nwTO/bmSbexho27mGW2cBZVoJ78npxUa
GS1KnrK+FyFvOtKP8vQi8RzxhvRz4WypieSsH4WcWFxKl93E5b5cO457ZMBlOAfe+LSOrzwPrQxJ
UCSLjUnpPCMkLZUhPN3vUFytUGgZ6e/sOvEXXP6ofqKRbxumdqVcKpTuZEwkDEtbZHPXs/hiYEUN
NAqen3UH/C81HCLRt+E9Mx4WpgvpcxU8YwiChmTTHpGJ+7TowaC7WQrKAngCHxCxyiBP0mYTZbsF
tvhZtpoFHMT0jvzWLgDrV4d1Ig2wy/gXyoYzfyLz2pS/zXVSHbnhDCqg4tCt/xr1DeUzGnqlOWxw
7zt85nUgOKMspmrBZAPXqviiFHYLn62CkOsYoqaw3zHnjEVMBcinkKgsGTwmgOErv2HVD7+d1xLX
sRiVB9RnxzscALeboN2dIrvYlYYAJiec7pdO9A4Q5EOJeXclcFOiT2BVVp+pQXEQA0APcJO2NRdq
HgnA4Akv475NAJJLT9LzL5QVuAhPLfVz6ZQjtm4bUxtlpF9UIYau0CnJXfYvwIRgiRCY1wy7Zmij
IuLtUocs7qdfQDkFRqQkSQivNtHpjlSPTMDBeRkeDjO4NpZVkVo3kZDf8D7KacKJURN6VudB524B
2aXzrnTHVX89/cBu6ooxpFPpm+aogkRNWee3aADlrraERs0CumL8BUss1UmErK17cXAIYLw4NoTb
MxvJQ34xnOUuxWvgB6Y+TYY5enHShnveWffv2WnswsuMneZ74Ko4D4D2bM2FH8C1wGOpDp/640Yi
tnjYGw4vgMsLAEgP+UVTDO0QC2A7c0ByB1K6XCs/AF7FZN8UBylYCldWbTiEDZA5e1iXgLTYnlf1
jmun84EW1U2Vup4RPYtlVkde1PJwqYykprm6bCaoxjFM8nG+2cTWWFThZqOHlZFHjVFmfcNBv0gB
Q+eEb2wUzf1Ax40mgQj35a7E3v9pKMCtIbqj4SHuVoo57hzktgnfs7wyly10oJySeN9I7CICHJHM
/egOgMWoXt9QeMHf1fBehr9GXpCODSobU8oENGUDuo3G7zPPiNW6mS0u6zLPBiGU4DU2EpJczGqj
gc326uOso9w/cncYU0zkCmFIjjBjomVE1gfs2uXUcZ21WwG2GyO+PvNSqc26gG/55LmXxla5Uc6M
LAZJ8fAhtSgYDaZ3oK8v5FCoDZYmKYPnfP1sUerUry/a2CHNdZa5XkbQpEDSdqXG3SwE3BGjXKna
jL20l5onhQHeShruZA21Rh4w2Mkgx31pJssKwi5Q/7H0Co1JSQln3RmTy55ZSpRDV6XcdAamMxdQ
mF2l9HLjB2f+LzDMBVrhr0vuP6nWbenY7WYv/zFOXz7qroXDnEaqJaAqwgU6vhJQ36Jy7hBtxc23
uXyg1KbvtBiD5LzM0Pc/bZ0JmFzwh4Ds3R3qyYKqO9sYRwLy96SxdNc/Vh/WiSqfKHeohfQLdeh/
r+Fm/vspleuqGQaA0g2WznXkQZpwEp9EtgG3PZkn40F3NrUld+jVBCE/BJbM0P4rJV/iFQ/8/Rke
gVTCzNIl2kqsvNZcltxcmcEG3O9YPWpqfkUUk6UYL0XcTy4pB5mXcWrgyUrRuH/KQG3tsbr3KGee
rkxSpllI3BDBwSXadjtPOJ+f/HK2JMr3DKFAXOsKkBuQIsIrMWuPbDPzqgaGZuqZx31Ae2i4Gec0
SeiyZEtTGiEYv/tUSKHVPbyR35a2Qnq1v65yv2VSj6z4K/LbhXSrpNFh8Gq5TbLUhxtyGmq2ZcAh
/oaZH/JXzkVgWNG5kPkdWPD80TDayZGtRXOiXINiYWU5uhHzkjVYD898vU4yyBv3NX4dZ7YinaoI
LU6cdjXpBeEz+3nTNA4csOR3doFkPrBjjA/+RsAnz04Pr0BEVBpssUcL2cwEcKk/EHujTPmVrjek
IMMIUF7w4tkbWZ3AZg22ksZqsVW9hzrXp5Wb/Kn73Tg6dlCHlSmItZGDDt5YO3Ddm8QT7cpLgiy5
oIMTWnJH1MfY2/1me7Z9bvGeFSp9ZxJisQ87gyw/GjdbxKYYI1+wLWpbJ6DFy3RcyKEVuFIqUzC9
Ll/hGXkLmi/yfSOLd6vGj0F4ZPN0vUJAmvICTPLMsmN7cuYX9rA3HGDSFzCsCqHcsQEbv1dlgZ6D
ZnStFbc7wUI3k4UqNnqodLTC0Dac1wl20Mtr1b1Wlo5ArVgkZck36IzIIHBFjjapQGULGBGWhmpv
sek3Qj0+HiuhkPNAVdlgd45d5vaAtIRIdF571RURkcPRSu9LDGj7zS3Hm0ASjEy8SBSONiKIViEy
uIxhp6ci3LoSdTN1I2Z1hKMXhZHGxUN+iG+I44WADYUv4y8lXoLw5W5AngeCRs8ZUfGEcNmi1lYf
B0Ujy4U4NIBTBANOJKTR0VuO6M1VTVfBthRF45975gqr9pnxqvtSiIUSzQQHOqTDQrfU+IjhVY3T
BHMJffi9gHwHYJexsE1yBT8hEBikN556AlJZQhlNHs28gwM9RB/GtmYaiwy1qit6QK1sTFekWbpA
hq2IZa/Gz3WcyLMWVYlhKHwjgLOBhUynAzrCSTuXoK4v4IfW1VrozrfKLudOEbdvDnEE7PtsTVyZ
1qe1ef7cZzCC8k+cSMtbp48qLMnjZHGE4NP2Ndrjacd0Fh8NjL+XtI2Ing/gEf1QlfPXIes6Rdf9
QWM3x4CGcVgQPInQdIYFSYr662/FAsLmN3i7hz4UJCJ9TRUo6zmMFFb0wQoLlpZnST6q2qJIQrw/
3FiZtprleUh4ek3QPj9m4g5jxZHt4/8Ni1abFuqAPezCkvPnlzpvRe5oMnJdK3rFwkPJFDll3ORL
jAN4kAyKHPhhdIe/Sx9DIey+U0rXBOW89iX15MwqjohEja9Z5450jfB8fLBnJv3DjAwXHai4uIvA
hjlEel+zlPBB/Fn0YcZU+aKHcJQ3R/OGzjjmmXyLDcmPRrzalf/P4TuSnvnhbqAyxEXk7RzgQT+I
TFaGunaQYc8iWqzCi6z32ERfW9lpkA4gidjPp1e1p0RF3Xq7JnOZ04E67Ha8MFdY0zeYG4UvZh0D
WnZYZRd/J0/UYyIjf852FcRA+ASe11mwdDD7DOAuFVX0uybWjhSKGkv+/D3ZmxURwlq6Xsx5fwx+
rmyW9nm7WKlxCV13RPe/wAOKOpb+tD3T6e7OHDbgWhneabRlVsIHSGeF0pREz3C1K/8bJ0/l+IRH
v/PDWbWPNRGFOAH47/3avVQeZnsG7k7Y34cjKpG0xFwSFVLKvwvcX+BijnKalSQfH7o+6i/We9f7
wJL7Hhgo1g0ImlybrXJKzbMAZa77+qRrEItZyrg2Gy2nedvusG+kEb9tvF3+yepJczptM+BCQNER
gVKfGL+4X7F3NhG9i0KUmijTVI8+zjWLEgEO4dey4BNZKuqzjiTQhcxCo9ijBJBEpZh274Rhxx72
EZISNzbFOrD8iZcMeOPSxy/q1LnEhoAXo0zcHllMe4IO5UU2Xm5/k12XX388zRtaYgp+aiDCxPnk
+Xt5b+9IMJYbMH7hfvDKaobk9e9O7cJZHP2OqbRSUOMVmyhFykQklcP0s+IzNRq2eUjtKM6PpeF0
3qiZDbmKGBid2jkOx/eIn239EGcvhg98NitjijssV3VvauJnv8Ub3uPAYFKsLAi1zVCq44TgnHLc
yzoQOwlSM4Dy+uP6Dk5eaWZcZY7nIIYZtjD8wNxxfpHobeonGKuuto6l/r/YIQs3Adab0BjBUCXM
72D7wuSf6XzY/H+hQO1HO97WePGeBkSKdOYonhljDvXkHN4fTMg+X1Mvuoe+2biKQrt+JFEpB08F
vR6AnCeKwDFlH0XOq4hKB3RiKwcWXsLOK6MKGEphV4LvjPd8h1pgt3dIa4owlFgKy0VuQzsMPH9C
5r3htlMRNTzQa/urZ5E6OroyDHNob/N4Q/FKeDoGTRys9AY3TX+X0YgBBlGgPS0lyAfqSObkLmAW
czDty7LTZfk2IGj8dOEM7SRXVwe75K/Huv15VuqXTE6+JDKpZ43oqUGxRx5msWWUZ69r4PSDMEIC
mNzga2cLpO+1OYfgfqDa/Dp9hrjzDuk+NOw+hfW7/MV4iONI7NC3a7WRCpalzf1hS9H9vTH/cOYd
Kts7AkVrg9X46NaF4kVJt15hNtvT1a9LnlXZ99+bMo7EN/Cwh/T56IQEI3Bh1dilyMFl1HDWlgGb
zkx+tRbb114isKMKa8tUHvDhYSKXP4VWJ9B/0K3pIlVp+T9534EvFqFZyU1EKwK+59bElJuDmdI1
kLm+RxyAyu600sciUJGDZzu4CtZOI4TFqIpEHF4tKUCPVh5qn25ILSFkzgu/lF+SZp8MqB8NT2+B
W1Q0dOXgsQ/wgpqvw0TLp2cow7+2XeYp0XGeikrmw11tTnw7nYixrJlHjp7dJalBghTzba2f3+Sc
l34+WJGfLMACr7UzLkWVzM52Ek/qV9JqBT/fMTo05uoWA5w04/2uJYxv4ePkLrGUu4yPsAobsPA/
i4VmgdgsdvWnWwBKE6v5CU7S6kaglZhlsJd3gbFQVtCSg/q6RkT2StYQphPRUfTNB6s8O3MV7Tgv
g04ZOzUyyuogOFc7EK44HZsRuCk1TKN6TmG4j6h91c61dtHn9EeCE5dyyBTbzS/WuT5wvJpvIfaL
xn02zkW5iTL0mo78iPAeSvGo5AhVt0Dc13N3hgaTsEpon+vGUHWCzJpel+7P0dvkook4ReBYzJcR
es9rGx8SijWUZxFRjLy2Lx6XQXyZBwwy1MfnEK7CGoLnXC6//Gi30Oy3prQsUj72YPFY/37mYczq
54NK7X2Gv3dVOe8KDmqWHWPdONKteDsSPgEPsoO5liyeA28vtf9k9mgwpEgJ1eEyKxfwXeiztuvV
7MT42EkGRv4QFSLjPVMPlsuBxYATwouqcH19QpIfdjwa6Obt0JCXENIuCoEOyW+qTKUNpm2Gu606
afvXfI6G/P6vNP4teqh3VYsXtdDeVXeeOfL8cJPvg4nZb281vrqcXtksQck+EIMD0aeOb8bDeFs8
pYOJqsynDodhvxLHnJb08WPLgg4OAyQ0RZ/yoq3TEVajfM02qSm/sNiX8KvDC4S4e+/Yj30Q+H/O
JusfW9C2+ApqZ2cT1w51tpYbLOG+TVwRTLOrejmD8w1JJiXRMz5E5XmMawP/a13Lq8DY7K+jJBtz
Pxb467RX2FOFiaV0oUygdLJYEoyXhM1ZAMp1Ql6Sf/NliI3vf/leBTDcke7swslyskqAXmS6HAJy
BMISMOE9+rYmVaojZLMM9+qF0/CWuXQu+AVJCG47IE2FhkhKh7HgdQWiHCABWdDBB5srhYb+/zuS
hJ/mibnqY+DJwFfcGgpdpHF7xgxd+3M7cNE82j4K/B8Q8SkJWD4RJzgYAm83wDRSnw1LRRQ9c6mc
poV3Wos3svTc9YxvrliCPHG8eYZIcP1PkoouzxS56v+6/IgdrGY9mEQdxIaeNGTzTbXEsDncKXJw
bn5XkW/lSsVnVlGI9atWCehf2oetOFhWmyja6bFmBjaszqcduajxQNO4bnDmc0+JYBzEKUIrJfiB
/R+nrWOwydrYrRIsDfDdzw/20G1bpdfOjU7LOoPJNn+8IfrZlCd3SRZpz9hkYKFCKBLic/2mEBBd
KUgBDg0nzptGGHZp2wPc9t1sfSL2z0IowE4TWmxxjEXa05U0+neihMk09lJgqS0rvN3HF8YrtFTB
SprDzRPdN/RQpBJFVWrRm1FxvdyASq3v3eaJYNy+KoIJIr3BLg2iFMuUphEfyGwfSOSWfwU0vRqH
kDtyzWNsXl24DbzgOYPmwBSb7bEP5ki0xnO63SBdDEkOIfiF8GagMQh8sO47QNLAFLbGCaXO/YXx
U7TEEbGoU3bgsye+mlVkaCOOyL3HkLhvMF2zptPlWnQFvWnN4TxjRMqhvP3APiGAyV4URZjZ5fUJ
KADfFkAlEJq93sL+4mSYyLkBIb5IcDnwzMMAvOYutu8UPBDY7PuW9FK6mU0t/69Qq4sBjw+UGKFA
ox6IMUeQiY1rWwsIPmK5umWslDBPIJpLh32WTGBlvumKsDh6qnFYlGiUCxX9dZFp1CYUW0oDdSfy
5f2yny9abpX9yl86WEwOrNS2VpKSPW1M6HLACK8t3MSlZFXoug8jpyBN/SrDKxbHGjua3QQXLdOv
olVBp/QAkYt9x8+W8Wsxr9HFs3V1jxm2nVfFblkjzJA+I8CnzEuyVOUWojHWo5slIOKfGOM3Kwnq
+YP/HTs52QQy7m2dIEsAKOEJk5Jgh7zYWnvE8slDN6KlROg3QoDhCJvmmSujRW80f3tC0osbb3vS
d3LufhVFFfKrZkxtiHpeX/Eqggr6BYiKnA4vYQWcQD+SDx7oISgLRPUsMCsfIag5v+xV/GOUfJ0U
h9/hEgxBTkh2cfegRGZIz6w7uODq9woRrEQOYEx00Izo9AZiN32VHHOsSVKw/uWoItIuf/v0oP3s
wUcXCwLx4v+SGAaFMAr2aUREP66jDa/7OyjDBhotAZMOXM4Ob2VPUGqs0vECu7h3P+5181APlFmr
QJ3mOu6uw8UUMKZa8UOIE7x+mOMdvmvcnDUCvY8/yM8QwNBR4civ6jYxpT845wFW2+Q/sr0CK7Pu
uXV3yz3o0ZW3Ga8llLXxQ7eBI2s5panp+2Jfp8j8BjJIw2wJvSnuBM4PpQf8rOohusolHHbE6yuE
4qVsDbreTFdplbESTBP5XdDIK7CaYjVObrwrQx+1XWeI5kzu0yBLTAkY+NSb/i9BhObLjcB/UT8B
p8RWl0FP0Z2dCHbmvsxk5rVa5cdKjZuDr0MAlenHWVXqeB0pUVHsCKscrN0n3f4TyHa3YNQB4XXs
K3xXEKTYdeMXW+qHun8REGCfo6842b0TUxqWZnBBkLpS4y9Pe4OmsMB6K++PMoycDf6UvTwZHXGq
+wi2Q9hdrXHwL3jnOAaszD2qUEMMN1BAuBKryVvyqSYeoAeXhLzc0SybR2aniq6YHKxJiBE/EXzM
x1zLOz4lCzjG3nmBcyrGLLigmBzMhjEHOH0fUZ/K338Ozb4E1E8mM1UuB8jNtU9L3YTZhUxXa7ri
4Y25kklFN1ZFRbjL8cqg2SZt21nRoKGStbu1V5pLf0mlGL8lZLzddgc5hgiHYRZVoB4RCWgQBeVu
+oCdH6Eb22mX0/vSfsZUROtjSOzU5ces5Uwe0OB9Ry7Zjvw2BoaVd7vauxT6QPmt9yXGkrU0icZq
Puf4K9Lkcb9JBpwWi4ZmkRHxYWKCQlQEHziJYfRfrAvV0ige0/f6DqL/KTqFgQOR3JwfhM1rz/wE
SREX68X8mWs47vXLqCZH1+4Z1VonNduYduzm4kDpx3y6IS07rhTUAu2HWjxFkSpDsUEsvqKgEQ0A
6IgN0I+KnxQeHs/sWWhD7vzKZ1Xc/x9rsAYhTW34LNa9ff/NrveogGSrWadkGCnwgf1P3LI/UiYo
vFt4xKO7YZHm2Ir08HTiWp29ezsBrWlfYsfu4FW4QMo6kOqBuqo2BPJJgsk3W6YM8jkcbCHd1X1S
zDLLBR2rwa1A4hjvgFwwa82UgEweuIu3RGEvHuBquXMZPR8nSXoSB5VKg/xmYACku2jNauKCrhJV
U8JM6WjcKT8T4xoAzaes4nmtnSWfVF7zrFLEFpB5lXs5hx2odoNYN/1+rAN82/tBSBLE5yR/4mQc
T6aWanV+wAwXXvEJ52jpTpdDTMNEgXdj3o+hFG4p09AoZvsh3e610OwzExLvv2tmVaek9/PSmn4b
63V5qAEF+h5GAPML8xd+PWk3zpho2MCN1Ne0rjEkVYtOMevRdibex1olQ7HGmGcTiVFaNJPADF1i
WcZiXZc1jr5Uwltv3XlUGSOx0l/ZooSM+kVagvE5m7eu+jUKUC1dvORaHv19sV3TiFy/HZAgBOPy
9yyLmQUakTJRbI0oNB9ns+GqhUBfcoeKVXOuxfsEATP8jS7Mw6/rSCaJl//s0w4YFwQE0r1BzdQa
E8A4upySBBMqjs17lZI5nW41LHAhq+/BiORdvYb3bH3u40qF1+4oc7+k9VWfbrLf/BGrvxGmBUeZ
JHKiNSSm4cr99WlpJOBPUmyenCqocHXTQU4KQ9dtxnarIKoEu8JMDgn4wOTFmuRAMDdaUZ84B9Fn
pYRtMCRMr4SwtIdGa0WiLeRMrQIkAxAqr2X5KGiXPtgeGheYpyStY3cn0EFKLvLrnaZC1osyC/UL
FB3xoHRVDte51LkYJEgCqJVPMveLnNHl7/v4foLhQkznI4lQp7OtzDa7y1ulYwuW99pLIArvB4Gz
L2RoAH2aFXltXO3KJLgEn0MQJLaz7AfMtMFlpP6vicpXyJvFjzfjsb2Bhpu3NUDBov8rX5s4EIky
CCibyKOMnXY5plUOShqfHLidaWGrhW6W1Va2MdC47m9yU5JYN5nHB1IJbICP7GkYbdOYm330jqf7
GIk9xzWmzVcXZslxVIHozhytMj/Q0eqAXfPrP8UgLR5mua4GlKN53xEJuGG4c8PudbiEKuX1b2N5
ODxL607xJgmaz9nQu6+GAlq2W7QxJ5cDioOXGrZWwUO/fOTbIT+Sf+9XJTm0/msN0bd6vV6MrCLR
FotH6rEexBddpQMs1CvsBGBsXQroa8wCCqhrShwYvfXYJt9kQVpDUxtBWcMv37T7XiGMux2jlERQ
riQa69xqe3n/R0/miw1mjeYdPe+0IYu4X4MwLAVSdF5EhUuIv/AV37wINGJjOp296S+WhJCkLkvM
hiVidADuLKpTexvxqUui7RvQKgvbkrQpB3/AUxlHjUmFc3Ln06Z4Wk3q3nXhDs/sZ4wqYMxFPaIM
lH5VFQSr/wk/SGNUcaeKVLnhnLMOCsF41tNuW+jPCwOSUklIMUMbWdq8PEf5EFKbRUWpJXRs6ryZ
tdONFBb8kleHyOp/TiPP5ldaI+Cx6AmgdJdyZqF/yuChjE+/zUIdSdK6rxo6yKzMVSEr0sC8HnEh
5svA9BL94QHnTQECzQswaMlQH60Ux0vRtNRemtLxgAhY3KdFka3SCPmcpL+ByyqGQyitd466Ncza
0VDOyUiaPV+mEmasHnPC3MyRVUH7LwpeweG9SFLO+WUtkA+R/9HyZil2FIWFr5gxRuZCUa4mKb3Z
ASkF3CUsdGORErt4DpZWlEEEHN5EC+Kx7vhGt8+b2rc3vhPxHSMm2phNDAkhJwe+bH9Dol3A/def
uNwsC66poielTZjTtSmvmf3mes1I2CBrh8xw7ya/cP0JOP1LuIapacHLlf52Ng5nGdG9tvEyw1O+
Ae8UUIqwpyJhmxBeEwTKTkPfjGXJduMmFJFKsZvV4GTuZKTB5GmcxM6cVPjqT3udjNGWHUxGw8NF
OaK4rW7e4xDa9gCY5UOAKV/PCFZpTn00irvXaQrNvr3vvjF5/+vHMU86aallMaH6+CmNHCjH5Igk
NrlmRtTblnon0N3Ntc7Kc2f8baM5I/QWfIsUs/9jK+xmDFid5XXP8XzGA8+JpdP/ty7pWVJC30sR
x/u68o9zTkEPrVrz/RzT5veg85b0lYa0atDOf3q+JTcWIAJv7vVmxhh4XwuN0W+kQBxrB2CwPMHB
q8RhZ8knsr7lQ/U6o0eLwITm1BHDZTwUfAuqANL1IHngciFb+jtV4+hOJgwzGh9KgNWxx2cOScik
vB9aCXMR5BVb9id2IyCWC08A2UhZw0KGGcJ4V++YBdZJSl58HsaRmxhYaPSVUPQM365gISreA7ME
pdnm59gz+/9X6zJO4mDKwnRqHhcI66spVSglA6w/kRomePtjZPh04Csp5ESAj5s0hMjhvbzLEF9o
Ug6IKLXGkhSUAoNGjKunwFimBxULChq1Mhq2HhovYLZhwdgxIr7z1Th3D64DaZB1gaCwMPpzu4bv
eHcevilw4CehsSH4SlzlTzRgPq5LXh9Kp+x3IR9s6ylFRklwsHmRmRBpnnG2hyRjdzGI8qzknEVF
mzAAogUfYscV8UNQ/8ILa0yvMkiRPb2luDs0PKyDlhHrVHAvE5c/1WRJhf9qkp775KCSsOOJcZLL
kcdhG9LXEy+3oQVSQMj/grzXiN9PD3AqpD21P9kPOevKzXuY7zqHC5dNAEsoKH4Hidu6L1ds1yv6
L6JyKkv9H9Q09tyrKxDBf1Pd96UkfT9f/sSvzNcgw8z9V77Sw9JhkuN078zEN8BsbLiRy6rMc6jT
EWVgseJg/ixlJvkkHNjsh+CC0SrDqBmdlAyNspTauCOukiL6u2zMbqkXALI4znMD5USjGVQlltQt
6xJckkTVORdk823p1R8TXwlnF5Po31NrpV1VbqnbOCwboKTFhLopmOnzN8dSwksL0+KLCJGwAlPv
PzgcoF1iPA32gkQkx9CM6jQ7IMQHZEwRoY925x+wmdcm413JZh3U1Ol1ITtXlfPYcIUSqFOvDun9
CPGjxYfHhFNjs8zPUU6szFwYwSWVttaGzO+6Gqz5KZ/iElT/3Pv5cZ7+xKcDdNxdcci+y2EfSe7u
eJOl0KKuD/vDX8L//TwgQAgoN/OY8c0OHseiRA/n7m3Q6Uoh9hF+i+3MWy2xOfcc8KxRatHlmY/v
mic/JBopmIf6YskxR4A5c8J5fLf+7RB69PEHDU0NvXh6li3JxMUBcIJ78oqkKaKBUuQ9bEr9c+Bv
DRNLK7dpImTGP7dk0p2AJhVh0zpM+h2KsuJf6u4e76NidkdzunYRZ0zUh33627i1CJWrdZ7El5b+
xv+UT5v9UoNPqqhMIQdSgsTU6lNMpbKJMS03WCqIRz5Ccj6CxWcRaURD5D6/hFvuS8IZ0weshfw2
ZR35Er2dQAXbaZP7fJtb4/JBibIAtWQ0ob4BJfwkIbQtx8Tq8LJ3KGdDOBOQ2tTj3PeEz9PBx8Af
Yr96p7Wp7hy9yiPKoJLOBomh/Ncy4fLg8BKqhwpt4ozGv7sDdSM9dJcpuqOhl7glKMJvPUY0B5+q
AGfchuHiqiwfYNAx3WSzgdekDGUNkiVtiKXxjqgf72D5oxeil1fVSaAqESEiNKH1lktxLM+jKOqG
COsVv+K6GY46Iz4h9KP9Vhpqe7W441Vo98/VZ16e7f/3FB8AmNdBzpNmH7LXu1JkES5j3doeqFEG
Ok1oWS1hjXHwPREZcbAls32vxj3RRJLZhku2oZ8As3M1SWLOFNMeyzcFgBQwyVH9BAiJYucIs0bU
nCFscyFHjzJ3ZsLg+ZsoiIMQZg7sWdekVtDAKjx1Rwf6KjOPTjANdCnQDyxyr3IpANcSK+UlZJLs
e9Mx/1ffdNmbjxnHaM4hGacFLA29ObUrLWnqBtg3xGy50SiTvO8Dgf7j295jCwtOGYzMgWreYOox
gnXN/vMKEUnYnHxLR+snvfJxzyZFaVE3AnanbfCEh9q4Pb1n3MVbTn+/RHqNLA7p7Jsp0RGsHQhK
zBLaEUZm2sy+3dTtd0cQ5I7Ez+YSZkGHQ00A78UiKj8R2+bmN+bn8l2P2MIckThp24gK3fEiFoVv
bPpVW/dTgasXR5teFogSsLh2LEKJ9YFitXZ5S39AvKNPw4e/AeuBBpDXpzhCmxobGdho91uyKDmj
riqM2aO96l4o+UYM330TxwJfs+2q21YesGP16deUPRQSNuaftUHNzR0bJbk1bbo80TwTtD4vacs2
vhdEMmMVL41HNuZsjCu9AK0tU7zvLBSUO3S9yNoQbf9knqH5NmwBH9FnZVNVTRXSPxCIku9BAgMj
GF5YqVtAmktRlakxff/mKf2DQTYUrPQJ5zgtNOeyigUBjA5joz9f1ZBmdNjYIJKPwqs+JgFIKeDS
Mz+pkiMj3GgeAYe9DOLvylsLmBGA+/vnTK7wOx3fNm+n3OcJW0zDT3C5OcXsJ1D03kWiYn+VoK/8
p+bU0rEpgMA5SG9oul+DxjFNNVlNybVt+cWQLihC9aNNX/9tIedznmohvDvnmoYBYt+s3sly8XpS
JEBd5mv7oh+NMdiRG1Jv4yhuG8iwHueL/uBKrpLnxiHCBQ7UB2DxbbCvQwllxiAuCsIqWOvgrmUd
Mg7x7j/JXW3CX3Yidr9+s3/ZylfxwCDE1KFIafZZ9788GAWSnm+YD84YtAXEG9W+3aV+ZRg8sPOO
oWScc6LYnxtWeHTlHn/TDRrw9AmprfDJoBf5w0Av0OCFWrpkaZ2aYnM+7OSO2WcxFXLnNOLl4dt9
H0xkjn6/8sfzLK0DoWOTlNRWwo0BY9e0NNxe8UqvpLb/iXZCSMkqYF2IDNhfdIuUHuVZ74MKFd0C
6ntKuGfOdUlWoDpIU+y+KU2aAWw9HckOfWbkMtR3tGKzuMkQAR+/NCq7OOI6WJATAxDztSbqENzY
44F+feRzlNiH3380N6wgpogyKFumcWuCDPqSFxcQ2ONVsgm5Z+hH/hHE0GppwwKC+w+EGhNZUU6c
SucAIsYCM5zDOAi9cz0PqnBkC80402wd3wboZNU2ZZMr8+rBqOxMBYdKmRN02vCbzt4/0pCaDdgU
47rVUfd1Wq5//3IeopA8xTMqa8zTJRalRO2XTxD8dUQ+c0GRGKmgHlW/fxKyiI7LtSCaAsfRE1EM
qnIjtASoJsS4fKUSJFslfLvDIwKOkCma0Ve25VsoAsO3hL15vb5xt/dr2L7nFckKvP+NgsNTU7Tu
w8bcIxGkf5d4xiXLiqfOcNY5+U4PgCeqb6IArXBV9ZsbZwLAmvzwhtjNB0qRpsVVmG4cm/1C66lv
0gLdK8hm/mX9NIMU7iRs1mn77f8le+Wm2/ruFMXtsSyzGt+mwsgG/5gpB2/mX90rWYchKQDnC7at
r0lQRgEel7d3Ge01H/e2mlRClusbNP40TfZZ6VpEkJsU773GJY36jeDoBDr9hQqV887BPxi74Z/O
AQw/trrDjqnUS69ePGWULSd/wzs99r7kDj1FY2P3ih20FRldzCO/cK1Er59IBUA+Yw/Plg9NqA5a
O2BoJHCql6wMNdNyaA6OrOTorQZZw80bsOzo2ssMUur0E9HIgv76KDn7eXvylDL1WWUR62hZgwG+
5fMVtM5NVUTvtF85E+uva03I/8vZXT84K/RlhBs4da72322kvyDzoxh7Eayjc5tHD6/M3+N3iVn2
I4G60A9+syIKTczcvZDRrmrcjPQcDTceF3xIBNNbX02SlSRdRIECZFXE8N6U6OMFjY9Tkdn9/vrw
sh5ASXPuUF6cSiYk9fBRFUOuJhVfT9vWyfo2nQAxVXIFj1qqkqUw5xwHYhVXvTaXjM4F+Z6bkPgQ
OSp59sYI9l4xxTKy4fApx9ScLD12D+CluFtUTKKbqMiCHuv1ieBG0w+h4f3iyRFj50jlv5mz9cKK
n+mKv3Vw+YqmLYdE+MQTZJCiAV6oEoOCHN6T+nWi4NC6WJXIjXvaLSAR8EzQUxr+RAxuEEZg8HF/
4QDfESgpTe2Z20OurNrXx+xmbRdGRm+cZPLodvmMB0LLJL2DB9171bnISDlbnS9o5p8q6u0ht3Av
TxeHJoWYFGVBoSuBWogXB+RGpbdTlzR4VWpwkgDPdC0FyNCytkya0xulN73dDh9r8gG6EoledFoj
cjLSwmcvRoSm2ZOsX3J9fAer3m1VtuJm+ykSQlNqJvSr6ivsmOY7ROCsL2XVvcba8+zWyQRyoSIw
kK9Lv/HuPcI0V+0aUfremJ6vUHmf0gPN6A+o3O6i7q/OVYtkKtwG1ne/vqoZ4Y8O5DA25GZQ/mGY
j7Dt53w0VoIOyUKXj3CC3886bcbOPWFGIuPCr9SVcZRqLiAU2mTUUPtgq34ZX1+wWeBohrJJ1G9v
oU+K6WhV59Jmr6611k//fAfLZIfkQ1Jn+Lf4Q7uF/v3sUdwoWbu3q/Sbxirp9miraP9B2zLVUHSK
Og2cs0bo5sv4yYLnpho5ZmaRUMx3RuojY7Nc+9pPVATac2HdPZh0U1LbwplFKfvn0Dk4pmxDOnOm
991zVyUSW3XSc/S1GuvXkd+GGHUW5FOvXiswkJe56tpVMewt4kWsj+DQ+ZFRl6b3F6sa9rJmDYkU
wiEwJAhx9ELapDkUI2EkhjSXJx8R4z6SM5+uRIf+F0UtcM8syFuGjQukaQpGdgSCcwxPAhSXC5HC
bpVVK/xw+hf+afZR74UEro1IH8FmyIMZ3yOGWx7b2P9eRHc4bg6z9Y6lZjW/OeRswD+LRMSkWFKP
0gPaxfyONNe7xR3XTwWUztfA///dPeNP41BhiuMdbCJTXo57I19DkI/tn3FGD534ZKSaPNFFd8Mp
LJK/WjqHdcmwaMzwfhj2vCciR/VpsXFpK1ZfeFe1nvpgVIU46jBhbjN86cJiBEFkoMc/vX7CeVrz
MSBvnqMnsRnQB1RYJYtUh+99YQ+fOFQ/C5sy+tg5AZxEqE3bH54HNxjOMsNQJRVByYMlkjF5aO3H
jNu6xHF7ZEo/2MJW2VP+gj1EjYPYxuE7nLvRgEVhayeWAki9qOH3gAmi7/uFX90z/ptwtCAs94r+
8QY2gHLsr5z8O95edj8cfG5nmPcRTQxA1tjkYJBHyb7PADwiRjsfWFq1HYgPJtGHoGGL5MmkWXYj
sJRCE+hkUxAJfognOekxzXw3ka4jjG87YmKLrFEdDehFi/DS82Hq4TA5T5iOcL3yu5emF0f9tJ4B
rHro5RMbHCxGF+XnIM7zXs0rmwJRYLL3k4Y67oh95q4oXv97tEev5d4SHPskslnK1C/HFuIoQoNV
0fZmuuA82v/94ZZxxZqrObih/jXxWBz0nQ7SLKzz8sFVocWti8jmPtqARPd9BQukgWAXv9MqoZcf
ybZQ6JbtjJmRpq4OOYHI6f0XxseLs4l8R9+H6FYZstMbtraV/YGH+Nuu6ATWh7Ec6EDE6BEqoIv9
TDiOuEotYgh1jcvPGh2kOPouB6aD/75CdcS1+l0X0LyF+avd1gtboVWdrcnCQfig33hdKzSmKXym
6vWUCIz3PQ65gR+liKjitImHoj69GywU2HzOoU42FikRTs1ktwtnOlLV9RbWKFAnlamRI79+NluZ
LAzJ2moZW0AC7RHCMVtj/JD6cRcwZyBg2N0NfICbxts7ivxYpGvt4NF957Op9Re5+YpPXnKBYs+6
3vNWLgMXqfmWKRGHIn/zpjAGXf2Sb+FnITGTKlKsrjNn1JkO9VC1jcJKqDMwCpxO+WccTepj5i4q
cR49Csg+6XmvIRdQMDRvF6YL8eHHvFSqOPV8POGtOpB6IEkl10NfQB2MjOKhBBBuDds/3WvjJKyH
/kwqrFz4+fivTN2fLgB1EEg1OSRz83tBYzmzb2+5k04FWIRGqJAOBv86i9DPj22QC+CZ4K0VNl2s
NbVV+pMQool8sZ9KpwyXcU3DmaibI1rs7vdA7ieq9Kgu1+WeaEUA1FV6v/V25rtubWrd0L3sTi1f
ZwyiScyn/Wmofj9R3LflavPN5je7Enbg8K8JFI8AKxja3BVq1kkIUM6BtQq5e3KFfNmbkmyreEdX
miiWSBvilyMBRnvGiNG9+v5Qow6+wJD8rl+CyCJDe/xzSGsZ22Fxet1lFUz0h5tGyxEpOb2ox22i
lGyJk4uSBj80uP3b6f7nLQETOo3lkeRD/YK8T9eT/vR/wBjng5PsRWbSTV1ppWoZYy3kfnxakHoo
OI3a7m6o2rbZV/fJiCrTnd2PVdvLpMhP+atVowM0xydx3INKz3HtHUj3PZRIhKdpc6Fp8woTVuDU
CQI37nRAGkm5BpvtonMNAJjz5WVYns96Kmde046g2gANHCNQirwVyLZzsfbZZslcte92KYwMrktv
Rq8LB2HvPm9ao0E3QffZVaMI+s1oTF0W0AHxilCNh7Ry8laOizjtVTPxMlYfKpWJI4axZwot4kgc
sUYrf1zC+rEGfgGLTOav6Z2fnNKV9ILo3Tam1hA+zhkUIT+bgIq+zRafTvt1RbEXpiW/95FuS0mB
D1BqiFlSFFEsw5vb6Ox7AajQgFRF6Ja+kqksweroFFdfZBvxJ8oYmpawHtmGYnfgjSYIYxlKQJ0U
5J5R03Wm32mqnbfzVybDOxl/To9i1g+xNbaNTrCnrwohmAzlqKLio1MTw0EjzY8sznN4jP5HfbQW
xn9iBvGYIa/+2Zw5d9i74SqhulTqRcQqE6FGWYCENMcTPQXYxp/06SXosmywpBRXHFFURhmnWeq4
p+WV9+G9+IvFDYRiduPEx4rKPFERD07u3MuUziPnIsKbck75ykgggMEvVvhoRn7pE3lu3eb6RLCy
5Wx6LxNV7iKbkXoOT2jFebXINeywJvEtMKji2CNTxeaZ28sML9z/Ehr4r2S/H0hVXu1gB0cXEzM7
8Yevo9J2qHSbHPv9pFwYjRgi17jL1lK9oniDwz1Xk1dqc7O9T6QheOjEh1XOSXbKVQjsyNRD6bAj
PqWkTicDXC55wKyf5G1tFyuSUg41wD01xCCQ6Rdd4rSY9zpE7AORG7OuZsHvTdmu8IU8X0BFrJQw
6xEKA4TD09l/EUMfxSFXem23F4NzQkcAKv/9R3f5CD9ljaxHvanVEXBxxY/jd0vizc4r5barwcWA
o2ooC9hWtBCC0Cl3INA+bk+x+V6EzeXiKjbZ+ePuxDdkfMP/6jT5iOw3462aVAwThwXBh3cUjPFr
BowHixrhtjigfDA0Wusp9EY4jyv28JzUHrlPCe5+NTdXOPlQ7CCrFMZg6KAXNceMFXZiXaN8z8BA
8az82W6i+RClSIu20qvGILO7tN1dnTsAJ6ht74c6Ig/1q81i3KgIc0mZvuCNAxJ9fStBcTdUByTX
QPzfkv+HCDAjJtfFptnnnrSJorlPlX8fJl8cE9u4318Y0UVOEbyZ8nkFRrZavdI9Cp3HiGm9n9G4
yEkFZil80jIP5TvaHYXRzqar3pseECskSjZnyTmYCNY2Gb8/bE3vJ0g/3ChYcwHZaN5M79icIeMx
zrxoUrzb7bxBHTvxSmJBZs9IEDfKF+5LtuS08BRbfeFUBRO/d/QvF9zHVWCa8OTeKbjxirhS6RLp
l5aP9bYywmQA26BGHtLPGC+XTSTnFktU9NylZvdGLZKFDPEWsOnDAVY1togn4OheYl3N1cUt+6R5
mrMT4BRpqZd/J9AoivmFnMK6lwMJQfwNZRqJJf0MJdtfKpcPgoe+5EBmLikITy5hGuY92tn1YUhc
9xlayMbN/dRiEAs2cYqvEK+pd5635EaaIejxzx/TC+fKnTTYakJX2vj5x/n4U3pkFEqoR07Icjpm
JrkaeJOWru8Kf7B4XsyWIUxIHUxbpf0zCxK7katWx+80MYKw/6lPr5akVoQBNYtAG4/9a8aSdV5M
k+ypqfeKEn6QScURNP068JcaxLpaqdErULx+CVogfN5Id8dF3WU9/OCXevMBubVh3UjSjvKBVd1L
Q0DH/CfIco2CyuaiSdehHF+z0IneoXV0doepDna2gi9DDNRz0tsAWPWjYzMiWi4o77Ewy1BxK6PO
qU6VKCAbomtug0B4sw6IiFaEL+dyPFWCmqPVUgykrRFqxXMaIDMiEYZqWgqdD14CGug7ieJ5dSo6
iO4P7JlcPOmOrJ82Y+bKF1wiEh43HMsEwLX8XlU5xOv3GHgfI7KBQjMXkj/4zd0UIkLhRqrz+Iin
dYR5Xq+b8OKKTx0tj/SsH4zB2GFjeehf8h9pZmO98QHWoXTNGLLL43RFt4z8crwg2yWzakgzGNBz
4G1ghs5s3a6+lE1UGRW6kowwA1jsIkaFrkUM/EV6WD7msxGfz1Vx2gLUhmPufACgzZ4we/pqYB4V
Vpal8r2Lis2o324l6Z5b8vAJopHaUEPYDaFIlmL4S+/p/66hIl/umfV+1mTkR0Vxw84/AVcKreLC
/JchMa499Otkj/HPRxPpw/gx9VTmB0ITMfR2U5EPdiL8ziX9LXdx4GNm68oezNA98fq2hjctzXWo
y6KNQvwV2cqb7ugzCD5EsbH+fqNJX6KbWx0Gzltbc2vewgv8q2EVZAtvBrDXCoLNAJRTeSahmUUc
tTZtt8iutbThMZAGOdCLf22Y03E9dexQGl25W81nYRNulJjTP0W2pC2Lf7SqW0K9PFHkPe5I4n7Z
bxpIrnhF68H3CLbIsXoNR071eyWrpgEXTAXbDwtmDceHdv+rnTFeZaP7GQ5OLzZzNgOMxZW3wT6U
xn9uC45E/5kogJ4uf/shh2AYhycTzYFG5QHt0Aoa6x1ceqm9HKlVEgxzf5E1FDlmB9HzFMlwhV2A
I85iwL2jBVe31LS6XEl8euwpzJne9Gl1efEI1tYb4lD5eGStTiVoslUK3yMi8u+lkS+peN5pqjh7
KQxE0Pln9Hs4khGiErqI2YoazHfihEjnDZRONCwg77wju24OdIZvAKG7jUtE0OhOXgkMzBBx/ndU
4sDDnsfQB3S3CzxxsTKekQatT1ACnKrC4HIfealRqKNW+Kj+Nqv4ELzrGSLKGORnbyAnLZ8z+Dg1
xwg8ejFUcuDe1gh4TWjPaeWk2ZJhTtkLo0G95tmMNF16yhj0mzDzGrJdbqiAJwFaiuDqA4DONEeG
IREhOJtPL2l5shpoMgfDKBHImLT8HqemA+P5bjxEaB9iaG2hexXlGpbFiEyrhh6rijqLr+wmUggC
D2xCmC4lEGrIRNT+wrAHAPolPgCsK9F4LaqeDBf6nJJaVTyXi77JMzGTsJ6yBsfrwr8ifgGUGK1v
k0o7E3Wkuw6k+RmEVXJK9ikLYIu70JIfvwCkFlhKi/CQKH3AisxgZABGEoFWdsBzXp0FoBYzhfE+
y0SCSIVunPzwVIy2JDH5jNzUC9O+Vfg7PljFqUwgwbHt3/G6owfz1gw4Sb/ivGqXdSFGHr7zHlXp
S4UtEulDMZR2EaFnP/uRdY5WggQ/Is7m/81NWcVZtSYYupedLTvLRSacQFHnpB9HHbyQFWlt8Pk6
l0Q5Ts8ixYnLV3vl3EPKOE7+ptEkA82TzVf1SongcFNMDGs/7Vp/WJztBCbx4Btzq2+5acLZrJWG
Alu7SDpWCeSe/k1pOf4R28sOaV0wsqTqVU1wXqF0pjaV0PdaGYQo/zj4WjJE+akwW6+7yrZ4ON1X
w9NzKCTgG72ggTwJC0QiVbPw/9LXfm1wQfxSvNZwfnxe39DKX239s5Hx90e9DUyw8XMVxDeaT2+f
JmGiUfJhF+uGM3ncOfgETJ+JgJbvUrcacC7wte3FGTV76nttbjqpMiatNu+2OkpU2wylK4PZjwod
P4J7ZQTPYKNkhzZ6W7HU3s5T3CSY4DofmCUwhcYgk3VkndtHIadxsrdFCqL3tMQGSQNh/CcRvp4i
hsbzbcQX3inLZ3/NbP3eZAsvg0C8Ql7A4Vm50HlEfxQYet9eAbkEl8ihXL64jdKYZMLz437EPIs7
UO9DyzGsDYPJy6VLdDfJBPGNtdr7SbdW1zyX7Vu/yRcFfQQviwDqqXKWjioI1mxtFJBTKftkngdY
gpzmh1Hi/jK5Sb5EybvW+iVRccg0r4RKBMeMMK2IswxTeqT3NBMHxc4qOhi4toNxzQ70N1wivbgH
cUgHAQwpB5DvCgjDr3IGNztxmQP0/yYBqzRM5hUTlGPPMTYtqhrNoSFhgSn4+IdLWqRRvkBz3maG
djSMahyN1QqB0RhIMjFEYz2M6Poi78vopeS0nX5tggHacvITOq+A4V6+PzoSr0dbfQz15sqGS4sv
eO0A+0zZwruGBsJPy8PnCnYhJcsylNf+qDRIdRt6MW9CFNv3TWqs101aEGtbVxWIn6Od8Dm8TUm1
h515widxdjlfF6MAOYcGPVadKfCONJjAM0OuBTUTSZcc3eFlUpV0MKYT5xDUiWvwlcOiZPIDABtV
tkZwM9DP5F64Qy0K69pEb6vp6Lc7NyHMNMmRyuYdq0gdk5CPX8DGP4JDTpyLg1YVzKwYAbsQLoPs
71HqjAQsZPmxgyWdEAOL/+fuO6hEHMklzrKdmYghX+4mtIUV3AXS561xXZyv4zFZ6AH/isZocpsc
MMu/D5SYPEEX618bx16o0yYTOvDF/xgBPydbHF77zr1NjHS4KLW+DIu/4HC7zDkRsya7SdPj4vta
7pkEEks9vu5Mt5eob+ryNUVkEFMqeS151VuLsgeWWpt4J/C4HPuzEAVwYrTDeu+8zbUktSGKC2uZ
U3hEedDk1c9Kow8t7j18qsplG1OaQc/ztgXcDsmX9RuCCIzm50huT22rI8evQkRHj1jIc0XTr43e
xkEJqTm4JWlA6J4Q4gVgeWX/4ETYotwGWyxIeZe0o1+qxyjE8MjvyMeZ700O3GW7W9eezi9773jd
Bc/qMDUPAzSkll6SCrwOy+C9FnzMeJc6jBCGnfmdqbiqiPgCpnZ7fKLHzATUD8w75Y2qPMcmCNq8
8bUjC/8XGhNU5JPirLL/O71NhFMF/7gltc1aBMxISqgrEMtYTu6la/Pient4dUANbLKrhG1rgRxN
FnDJyhuRtXVThAM9bl0Z0cKuWgjR71eN8Z55/XyuEH8NctnuGC8bgBE/h1UDPcs/P5mksvdjmH+D
D6e2ZBz9ldxZutIxmjYBrn22VZU4M/Dk1NuhiY64sE1XXeF84yHmwpJBCYt6ay6q39M+G/Y16TYx
eiQgDEWmkBwWEnI/o7nIsJHV4TFZD6bF9V+DXU+zmLdGXpTFoIDXt9ccdYl9nL5zQrVrdi7/ByjQ
bW/CUpV4xt/aL59V8uKhnLoiO0qSoL9Apm5P8HmgAUDnogt4LAugcCgy6unWWnfIcs+/6dw0O3cz
dQkA3cP6yluhJJCKWJGQ1Dnly/6epqEajwt4DiUjEBLkWvIT47L1f6g8ikFaqNNWPnP6P9F4le0G
Pcu7jgcgMlg4uojQUJ7ExuXcMiFwCtmaKqh0mUsXu8SibUw9aETk84hF2wY5IPdQqqQyQdVX3PQL
cAFpdKHfM6fkGCh9ngQB1IZaYrzBwv6MysVMg4qKauQFHxMarKiZg7/xab/R5hRLun5jh+WHuwQJ
63IO3nX1wJvm++GA+6POAEkffOMyDTT2nsveUGuVCvyEW1j7Q/Islc9KgItIz+yY79+4ftNzD7c4
EkKV2ycMZ8XKgmdagVag3UID6D1eFe5AIC2R5Bd0LYtW0Hi6ynQuoDnv19IJI0Hux5Hv/NvFzB5Q
04RhGgQrXjOFDMeVZ5Cgpn1bSSXduELXU7v64AtlNl/gVkbrvcgFMh1IMUyJNgQIOBrN+08LpyTS
zMLq8NPy38twSOQNk6nh2EsNsgCbnJId45R186dsR8VmJEdNp3GW9V4xIffBP8oHl+BXc9hhURas
BrrWxoRg1SEsqjWHuG24BbspGB2NEGSV8M3jIhvA1IemFmMqzx5mG8XozwUKoMi7zvz8I2/EVsFu
KhTmYC2kF4At2lLFTiSGOH5QlaMaiaqbe27Z09lOIM1VHTHkPXDfFYxtQhDblbRBCQxauXAEHHTK
5RYaMk0TbpS3pIgHkImCybgmLqqell8jGttVPh3HcQbslQTHD8kmBuoQWBJGDT9n+dgI5YA6yizR
xCEwk4NI7ne8TuFuICrHFDjoaxAxQGZQH4lxXAPagFPVfRo2n4I0DYjnfoL0/fVCHt4OSF4QFoWf
yWQgdpq0ssb3P01/eV0p717ziaoHl8S/orjO6tjONMKbEEGT/sdfqQzyjEf4LmCP8RsORzg3Vgyl
DmEQg2Qnabk1rmMwzEBNIbyZ9a8smrXS6qoUCRhpqoS4du2ZY91w/uz6OwZDnK6FT/m1o1U5IZI5
qTfidydDzGR879vAxX/OqZ4rcYFKjTkDs42vzK9j0cy18BQI4FrM5cb/8M98M9siC+Erg4cxpOWY
qek+2TzxJlVLrZinKmj47GC0w7A+kYw/NP6q8qIWwuBOlft1h+sSX1u/iXdoTlhfeKct9/4H2gCM
MRKDawDoBfLZ7/wiMPpGxgGnKt1CcJxUpNMW2ro9VGj3ZA7Gbv/NrTkKaGwvXGsrL8Mnel2ZItJW
HLcSeElQASw9oeC8VdU6kwaQNTzKKLYtq4m0qOzR8unRBbwXaBxgSroHADxCu3H/9W6junQHjNOt
hYtK0g9+kJjqcU69dN5z/bHH4NZPEaRVzlTVfx7q9h5W5O3HJ96TvjWtulwwSc4hrl3B4BXkfRDf
gQmJUsCl7sAYhXro5ItQEA8y+igrKeLAn2MCgiLUvROirp6RBLwc3WvsFGgCzAUnM2EEpq4xQVFD
V7n9Au29y4iDQf1JjNHWi06hbrASPCgm0lsE03joBnhRYa3wkqnnJ4RbAzCr4O2s5hHwTDWjysuo
OQOw4NDBs76XPx/eVwEfWIzygLPbWvUdb8Kzk6U7JXLNnvMdJsgoz1WW7azsdLKgJV7gcRJLZ5zh
dATYNdTDmcKlz4UB5CMdtOOs4Bmw3h0ok7BiDLSxcuIHRATFuymtJx+WXN4i/G/BQRka03p/ifHs
+uVzkSkno15FIkUuh7x4VXJKq8NZZSGipTTxv9imeRrDlcmtIkjSlEXcD0R0dGHwckoIcXbq0Drb
CFdOM3ODYi1ZSTauznOe2w9j6jvB4DFwZNqyq7E0zseTVfXvqy5mx4b2WmGbrYKNrFrsO4ZOlklQ
uM3+HzW+IaFIQ7dYFsCBoSocIbTlWXAQO29o9OnZ8EtW/xVyiO6Ktw/yTXHX1CDnKR0Wy0T/cr2h
6qa6pFO9g1qHql+Un9fKAAMdL1APx4GhbmMMopPaQ+1GF2IRe5k+2Hit6Z1svKYg/zFz7LCeNZ5g
nEpQm9IOumzxxffQGwN01o2s1RxQP/TGNuhuxxeEE6rJUlxg+4LBT6e+/RMYrF3c4N8t92Si4Mdr
OUNHSrMngJUYo5t6j/rATd+X+r/af0hjHApMbp5DzQ7obZjbb9OS6Y8VTjLaIgPN8xnT4URl9GFc
lY8mPl0xP/vu4Q3tyqSRw8kuvZVK9E7z7p20s6253+rvxFHcwVpQqTgMRTQcruEbj7+uvQ5+ZJ5/
RNQWzKFcp665aPCJNz47aCUabf9ojJxwj9sJSU9zbwVvuabVsKP7p4pyioOmKyVTBl/JMnt8s8ya
bS9ztpuG940Vu7zsFn6Bnz2eVkkxNZoNUg/iWam7setigaR7XaLycUKvKMb7LRWn5Ekq0ibTYJWG
uZRJ+oAf0nSXNtJ/kTmRw5xmeAITzHmJz1wF52k7TeRCiwogLRdRJlSFljUni21sWQKDEMc5YNL4
8B+Rn8yXUUBAakU33oYHSPsSDOYuaik2to/vhMWL8rmnZeAaTKgg0w99tdi6RAED+dNDvJmVVYY2
oAW/uTNqywFG1JC3l0Icvk5Sv1KJRt4RO7AM1ZHVeO+RtT59FNzW+eUwPJB2/fJabRzCfbTIMDOE
8gcFnpEwEwo9xh7eYI/U+22Iqdji1QoAhbzhPSA3TUIkD1BGsMSFRNQPEGHySdnjxW3xI1MQwVJP
GKLATtwYT9B6qrz8pHTX5ztAGUYAf3Cp766yMyqlyhryyv++aC6vQP0bO+3NXMG8FsrKbETbaVWo
5uKWe9PBpTdBweFXXapHOaAa9VeTi+3XqX1Pt6sBoE31Uq0A3geNNHGdMqr9n285nuLkBM2oaVQk
Kk8dYm8HmDk9eWhQzTgjP926VvbmPfOzrsLk6BReN5kEC+V1xFGiQgP1AD/Puhw0oobnRN1g6PzY
v/XTrC3naMpT6jyj1ZlqvptWE8Z4YhSqEDnHj3mRiUMLopHW6FmotIcfpYAC6q6or7NnSAm0M3VF
IoQ5bYd0ZNLuqal0j4chrr6xV+guwS3HzFpgK2o9S2wN1gJrkvuTXyFHBZuO8RcQoPOYVw6ImCWY
R/HQE9EEUhy2ykBQpGk0icvgtZo2FMNvVT6PA2/kGmx2MPDBgItQ9iKwy6ofpMIE8aGjmG4YKk5H
4TvkDM1CWRwH+J88dxQ019/UYM9nnkoQ9f0V605x9vQ104M/L8rjo53VEw7ex3m92wMnYABixYVU
74vYMw+HVVJAuu49pwa6MrRGWHvK6byHkl2yZVyQ3DzBdX0Jp83miESanl7pXs8yQWUaORgA6FiH
O2WbHXhDUQzN3PrSA04QEbPC1SXikK6TdvJOA3aIZCHUk/1RHvjxkrEX0LgHN4De7aM3uSMWyKBK
2GuCjoVOoiGyr60reqHepgwIviyihiZksIP3hfhWbBAOJKZ0cMVdj3wpWXrS0X6dMjEA3FDl61jg
2l8VRUJTWoUfZyoNljcoWpSzslwqZ1He/3QDS6RBpbxgzyBYjsvvuKIgEpUxFV701CZlMjoPefxU
khbLDG+H4LZY8Zph/9EGSkIabV1QSHLkEMh194vJ2dfg8u5yNkneYS4sYHmA+xv+ATd/thSSSfyR
Lhukt05XE6NSXH3BfSowC079Y8Yd7tmVaCcpy/0pW2LrD5wH5EmLXuCkcUqepcsYlXihbsn3/Up9
rz3/1+6PBFj0Tn6Zcvt68QcmSDnqw7i3CgSZeHetR5lmDTbRfLAILQvQ5O3+/0XyqN+cwl6203is
3NTCAIz1mqotaut65gfH2l78932Eoypgvpo0kGN8YvpSxKpL57vEJNje8FwvCPG8Pe4IvbVslVRC
MSjI0TvKVPwZXXGhADWCaxD6ZRdKp0S1aAfTX76AUOR9wuPPWs2F+WfxS1oojW8cMNFZZS5O+Qbg
a3PVIUxeqDJsZdx6D9ZHMLwignRL0BItoNM5TTb8cKtUhfQYHCRGeiXbIDVvDCgGJhSrWKvO2KvA
uwc59eFhx9k1C7+B6XaJ1P7PuBexbkyIVAO09/3ibXM80+0iF5xRUMyKxsIXY4DfoDfVGh+Ae5fL
lROqaPN0H6bQjbUC8j2rzOdMTVxRUys5hgz+/EexVCTyrM7JX5y0wCTmKI6iWInNj8IrCfPMcn1y
vcSqWSojPjBRdMd6/0fMD0iNpJW5tal79xRQcy+7PC+rQqsvGvF/oI+HvY9Eg5bkCT2lG4UDXHvx
eP2WRd6UFIb5gvIMlPd/QxG0/VIr0hOSdNaSNAgLnmMEdr6aH+wawOO+7PyT0qvBdnf126uEDf45
Shs/4tq9UoFgWoYBmSC2AwBeUhAvtNh/n3jhrGWASFJHBK1w3EiyfriZQjqPtkFieS/UYdVvxWHk
q22kmTRH0DEzST2sdJDzUx1Fba3SXLFsdZqXqZnzxYvm0ymwmNgF0+VvBdz7AQGb9fZheMeSWmMo
6QkOGHAED037CRmcxMd4ajD2rNkUzKLHXgAuaj/odW+aR9Si/hCj9gUBIFN/vUR9vF5H8UGgibTx
+Lmq/Scttmrp0TiyIrkohpHlVgayvkRhlaXAYs4Tsvw9G6l8AJPQcyPhBBx8vGWAlUMTnWxfuj54
peKkg3bB6zoQkWMezTBGNi+W/utYhviobmoLeliriBpvMTRqQKrWmPQ5d2a829B9Hr4pcjydtUbo
yg1nFZk6NyW1l135D6Ksqwy02ZYuS3+eM+pG3YdOs6FrHMJ9Q3DJMrywhWuy0hJ5XBfaf0+yblxf
8A/ydMsQuWkOozM67ciqZ1tIRKKbT4Ruf1pxoLzQ5cXMVfymEua5oE15wbszhl94YnUEABMdGDB5
FkWOPiMGuhfJJrAd68GzklvFw9KmC+SwgvEDs1p5R0t9TsXZPx4YWnW/MldwrCh7NPf9h/duTtDt
d6z9xH6rAuXsTYj1/DA29QUSI4Uln3gJxEAVlrPOU3VznEHjs8tXN3CzjKXfTY9cUwoFc0Tx8zG8
UT6KJ6cBouGrsgzna/hmHxcfiqcF0A2VL3fsyjhkMlxoW2sq1AK/tLV4+tMMfv2Nikfokt6Fa2FI
mmDEToVY5X6bzT6x4bDaNFPpBOStfSisRLdMxoV+6VONKLvzdPhBxO/A8oLGFCqSL13mpDxhG1+W
44kN8TDqzFaKfiEHsfwoe02AGJ/t0zTQP3FmGe5sC3+3awPaqLUp28b9KRadharM3oYF/x/xKIcz
mofkw4isMYgiD9RWYj4f7QX8c+7mHYMHDTTraBYOyA0PyyiHxXBlOSJycQs10zjErkz0NXtl/MLV
9c4BTVrUuSrk1uuvC8sx13Ysq0uti4WEn7ZgXNXROs8UfF1no9/oD8W6SI78bOojmym1AF2jzyLw
LHxwcbORFsC3DOWNdMLDVeyeV4EQtrb+Aj7lQaBiAPPiX/8/BiRESJTx9myXo0gyFG4o7P2u0bXv
0tCiRB/qDZKE31q5rSJghx1vyvTWCopAmTuODlwizkatafwBy5N1UVlHW8QPjre3y+FWj/R0SsSE
uRIvG5N2JS9P5GlqUTnLZ37Fx0pfE34F/SJRjO/EpQJA9z03Ea3Bu+guhUrWyI0oUzxI2jVAiVdS
YWCjqY+ztZaM5qt58GUdy8vUbEBDpcndNUyXxdXfFKY2qS8DyTtWhih5ngWAna4f6o7yhP7/k92z
oLz+kJ67VsDuGum20GUQB0nDZL6Oq6KIyKb5Ga07/HhlzvDd2pFXvcbh3LzTgZOgA2Ya/0TcvnS1
mqft+JaD20FvJ4Yii9snC/n+iNCxWrux+v6Z+6OgXUIJww8jKjmGpBirRW6ZEmHtIuGknQL4xO56
VaR2cJrCegrV7IanghdvNMXzhM8YX27BMOoGhkzfLqTdPyvtZT7NOar9cNd1A75ROI4Gy3l1gkGf
FiSF2eEuAhVWJgTm9WQIKavSoJ45es8pHC8LrxqYY1NV69GXz+4yToCSZSIiTWGwZFqSXdrO7TU5
tYjrwwUlwmukjybx0c1sYS3jGCseo83cF8ipLSfG3eliv62sP89eN1FoMYYYgmEIQkJDZtwhyu+L
zHbO9I89NwEGljHHiiAu86DjM7HrhiJqVKN3+5u4cknoW7eCuiwaT/yShJYokoRhwLXH1msYtRxg
RCnNw6tUWd57BFf31Yp1wYUyXniwOmVL1CefT5omuFea0iFciozlNoQksd8CMH8nGaZ318XHPgKg
a/yxLz/tb++Ed9XRFHkxRqpERadIkq1SyxLB9R8lk/bXw/qFboGb6EitbJkGUb2jx9dkfmDjSdtG
n+dTMmnkaONfJ5VWYFyZ2dxR86fzp60jB1Zalk+I6oMETWw2B8xG+GuI0mitYmmRN9txmt/nICeW
0sQS8jHRhVeNW8LsJgI64JoI/m662KNldWy+E41OazIe3hNQaY9gqijE19jRMROvlt0dEbwhlKsA
UdU9QEowsS++bGtCtvYVmtM5MvxaCQ4wpoB2FM1MPScMq9UnNt4aLg0FOIMnQKaTT0tPmG/rDhxF
zRdAEwv1U+9y0ryEDsBRLGl7lA49NLWIIqRf2+xNLTvQ1PAOwKrfeax7skUTwnqg33pJUhatCBCh
nyAweUqhue39/WwOKT9mC6MSeE0YOhMTVmdvwX8Ge+Pb10mvf1o/GiUFWDXMpk1UdqwyjVQECEs7
+RuJbm3RdK+AIJ45qY8iXU4B8Ds7/duWowtLMYz27vAauMOkWPFIzGhiE/izXua28F+W2YWlE7zx
FeK9w+I/El5vvaFqWsu0ZJlb0AYEHvqhj6X/2gobgoclX7RLpAliEfT2MrplXWOw4zM8eMt3fZ/N
zYVGwnKB55HGi5dWfFH7WlVP+riDsrSc0P4TEyGzb1XyAAUdm7Y7MVr/9191MQWHbS3jBN7WLInH
qYL+rHpwiuG/+S0zwjOOKmVr1HIVE4OMgi1iI45rZ5Cio+9gBStgPsR/zpFYSbGFHvmGHA0ZM8kO
5l8pidLOuUXlugJAWf77e28lvO4oi5jTt35OdL4QsAjyPV4kJK8NNijdPGQmAC9/lG6MN9eUNq4l
IcKShfTVcJtIers7w6twZC+zXlkmHvljmM0sannBw081jog7+rxIV1IWHk+q5kGeLyss5E0tv3wK
oMDWmVngWKpYywRtgIdTk6iJRQBRoHyIJh94um1EzQBjIFA7t+1NxGbAT4zWXDlxcGDYTqQnlwmI
abpxF4LB5wkp6UU9kGXY3BEtX6sd3zMpg9O7h6wqhMz9KKMFVtzYAaxu4/Fj/4XYKBe/K0H0dyuP
B1MoWS3GEmiPye2OYImvCJP9t5sx6UzVkfW6qRcIj9woo560SrevbfakoG+rCDk3y5TyUHON9UYP
I3G59opSUSyfdQZI6BKi7dlF/7/whuW5juy5PVg+cEFVYhr6J24QhCre2DOLyGZoCKF57x9geooC
pnS28Mq4jPisS3fDT/Ab9yv9xi55Jgj6aGrGoGFAM2CDExlgoRcjmRNtE659AiJTOqkQViEBRxRW
kY7AB3Se4XGKwGhvbpsyBU6UdBOZm5LKyPwD2yQ5GG0oljZ2ryTH9b6NAeAAkO5RiqL7QxbREZL6
DA/JiZDni0T6/4OjmG6h4LoPIyRXX2ums0VoyaElfb2TmNjI2m7H7hTxSP4nPf3CkPeV7gEZ0gxy
b3wVgVXPIk/5JieSGvKPMYM8aTIAFFEAgVlw8WlZL2USj9jWk5E0rjnKN+wUzlZnZF7LPv59ozKV
S8xoTP/FDea/v/nvKQNbnkScqJHJTKQwS1Q6jShK6MeaRBeJDb7M2cxoXWQFmPo38PDGvQTKJuH2
wE6VIfouXEMK1AGqWKcLhUU3w3T+eWpfVLxk0aX4Kv+UGFITKVZZlJ33bytN2AFXlAo83xMcM090
Ha6OxMBjOXyO+g1nIs/ddmFpb9r13kx5Az//1bhFwQNO7eeyUQN8VJi5veuoNzbgQHFBKnqmCrOV
1DCzOQAkb6+8Vk2T9G3zuYniJGaKwDg/dgEHXj+Rag3Jv9iiBugXxaJhEZOJaQfW5Etmo7/dUNDH
fGg2WTR2InBLdwPFzjJwT9WBQg+VaUIW4ZoD/jPPsj18q8B9YfGNUf0f8Ed6m+9amkAB2pOd7iAc
4m3nEPT0I8BIyGTdYHAeJDeCH2JC9FafYGQ1Cr6ag6G01goL/NbMofbNRJz573EIm11mJUjM8pYz
/EyG9MTE489hDG7fRkxTOjmyKFpOuvq+Bg73NE3kKRe1DvWkuz12vLZDlhQhPWmb/+Tza1/OB6uL
kuvJFvTOOrXUe402EnQFbGJtY0xWILuIJIGoyrVJpJAYAr2RE/xKAF0Xvkml+00XJHqiyNJQ1g52
h3V6jQqSp1hOd+mbqMOUdVyKZAcktl+mKVvxYmO8NIQiYGfUlcVSBDZ7C93sEaHeziPMhPJGb0fy
hEz79EN/N9Q5cCjVpZMxIl6NXAyqoxsUvTjI2wsKxE/n4H4BAx3SF6fDJyvi2rJE2ZU60k/bjZtn
GtvQe1CG/X/Y5esBuXQNw6xwe55mH7+UxOh3o9mM1X3X9Y+EBA0PxfDpNCoDIwz/eoqUej9VsRmB
hVjSqamB1aMOOlpPe+SnjEDQp1XNTgFUl7KMmiFDnHabEDcD+JrKc4hsGnrqBrra0qfsHTeI1y9T
JLyOr2j3CzvAh1J4Wd+CURor70F+ECN5NeDGTF0nnug1WQ3yTA2N7yqnz4LaJBH6Yx5ojp//BC6M
7VuoyMijWjJRS/IM1fQdq+TVQRTdZ9aYHniFFsDvNZDbbN0+XnSa3iyIu1CyYfW7mzoY6ssvW255
VuY78fguhNErnsWDWxQAInaBUcPBe+ZCHFjH3ztffc1WBXb/wZE1XUAT1hAeMpeWPJun/M5QIxOV
0TqQREBtZB0eKQJWSBXL8OPKXojMgH1hsvVa0vgowfcPzC5gIPmKfZ+KoGD9d/moZmzpQsIM/UiS
iAsGPyHznVelaU62tXGn4EDGw7fwrLOpdtlZ4F4ZUP86GBky7BZfKQmFuembE0Zbh4T5KfhDnyI9
HjvSd+qQkAE9Rvfnw58zMJj3o80f3IWS5fsx7jsS+opFfOYYxVzqi/chdX3No7p2Q1ICB4AqSaTQ
Aknt3gxc3uJff+QEWkJsAmKdYfE3JQKw4YWh/jf7IjvDv5PXKHUq7DrRkJIMMA4NeA8ZP0z9cPIo
8PQv7b+8t3soWT7afvE4V7gyXX6Kh2So9WI0CFPUAP1WKvebmaFfy0bSBpeYJnUN2aD+TdnNDLH7
NAiq+Rlw+VrVUn7gEV/Eh0uCix+kwkr6nNJHzcddqXCmxV0JLPrV2OPzriV9RqaW7NXPpP30FX99
YwAIjywmprt41aHXL8ZtWHlxtu/SOIoMmURWievkGBAzP6dZ7wzVW5cElXtWOEUdEjFfkn3eS9Ud
GeHGDkLYCRBWinNTgnbpzBxrwEDmkQXQbd5CcijWwewrn395xeoMmS7/laE70bEJanm/8U/3UH/7
lSK0jTSF+JrVl5RrwGgqt91AGZlDILNo5+QFr1LHkSws0uuDXGzwLuXb4QqEP/drFVGOrMpM5gYK
NsVfgqCyBP2ogsRWyxOjY6RbARqhsnFCtMCU9/RxrrvGJ0q4GtTr5DOdFbanXhoNNEBupyVTNKcb
hoKlDsR7vbHTQn70pggdoBfxbtPENs9KxtGyLqg7ACQVw3QE6XJBP3LY9wwkI9I00eG35We0xxs4
Zp6nmvWYttUfBMs2mpKEX0uPBOCfiJgvPq2jzztMth9umXTXGL+j48L6OOomjLBGlQLPIDX5QnUI
huzKH6TYZoBWcRTrpRb9E6eUsIqBhQdAROekTg2rW4t2ZN0PK33jtMzz1kEJZyLH13it+BAq/eBg
zXs2WwgD7/bib/rrC2FiwTZeVIumSAoo/raLp5OBCDpQ99mdYfcaeAsms6zNwC/4c7UPMI6fKZcb
cwlm7eIR0HOfA/nFpxGZ587ScOxJsOcE+sXZVq4TKKjJxps2OgDvPuToA2T2YBF3+0OJna6IOjUG
n6jhQdqWeKOMe7SRJqxflF/mPwuMwvTi9reRuejOQRTuZf20M5FtCk5XyMcxK7rjMCdVcrTf8GKE
MlosxiClazhkApz0eAh28JkAM9g+WZhUqdfVaQJmpacL90aIX2plkBigTGZW6lkKVKV8Tg2UK4bT
GRNLBVh+A6PXDLgK4CRflMRKAu51wgsYQweN2cxGceGOovImtmPX7CUplLo5oSyMrfJFAHiFAd5E
lqI1h8041UhQuxfS5YskvUDFvWWyeILeGHaOZ420Y5r8mqSoFWm/5FXfKvPGDRz3PuUNXy8IYYei
y8pQMptmFj9tA0AH+iJSTZzdbCEKN4N0t8EWuKq03us+mDZXQDQpDSAV4XTM1b5xJYxM5ZSjqbmo
4NyLjIddWrqDDtYBPt2/aXVjO28wCLLWzIJCrlR0r4iG4DukgCfkI3RB4WUCV3zY+1BfNybB5+Xv
yOS/JzPYQZB0Di2n3KeqZ++I4qNGYeX5tTmlzFq6gu8jyn4PPrgpU1d2hp7SmsPKI2hFEkAs1rPW
i7FGEQFyB2SS/PV1o5Cnh8Wzifzq5LlwjoFBpXH4aCMcl4QKnI1pFKF3Wle0Ca3eHfXvjiriODP6
PM4wXs13eiCI7fSXT5EVGVYtABoMzH3reG0itRtvlUXIOwCIjuojmlAUFzo7IzH3kP94h8hoekEM
cFMe1sGNhr/byTZzu6Az79J+Ui0zgbegP0shXZne9WbWvx4e5WPcTcGfLlF14M5O3DkT2oRb8fFj
L1jiC2vsdtpOklOY5HRK9I/sM40lYLfjf9oUU90ndbNNCjy77AR7mVlN8G4hqutzfUPEipXformr
woDdZWmBp3S6A6IWpKWvfYRyW6ED6ToQMc5qkGxcC0keV1ke05o5mm6E11zE90RU5OSWq7s6o2pS
J1KeIIatKqWi89L+TYcehF0QtC9KdFfrxdXs3HXYTUoZxB103XysugVVvLvSOJgrVFqbylXsN2l3
+cU24Ist1TGCi6SvdQbhk9COhhCPc5cU/fZBX2BBuLAEiFHMUhG6xZSlOozicXiM7m2MevYxPbS3
Akz1OJSYwQgNCYCUyim9yOeCxLBKwUlbagzhZgb0U6msnGcEPSW465i+1nW2kwXFJR3qpSacEWom
ArMrJN2cjIwENJV5nRlIodTuUDsr4zPmd+2oCXYYazoN3pWOIlzs+IndNCb7vBVp8l7A8kxORBQx
/ubHRRYgEVZiNIKm+FXs1G6ifXpu5prbkKqKx6iK250ccePrwopTzNGBrbAeScrCo+VYRTqYHVFM
bQ0vYe6+WPP3bx6JYtk/y6bK56VvRZuCCIT1m/yIhO+sbC70GMiORMPyn2LTnXCxjEx/Dmfn5OMb
47X6u32OT86/uw1SRmv+3jEA5KUqBGNXhgFYk5RrO66m2SnO4H0wAv3+IxCHR81uvsNNxS/B5Bg1
Ku9kdkFgTNKyVdeaetXCXlx1Tn5SB5DEDOkg+HPZg+FGNsYG+FrItE94HvzkWHRnny1L6AXylUAO
FPxnSiUNxTxIH64msmgkLt/e7hcaaJjIV/9naS8XNQYLWgfJxWDJwjHE6DTCP0p+qyTht4dIgtkb
edLI5aePSeuMTpI72u1/zK33yLYKT4owjaZSul7h26WFTH/kZtJZfgsRhPKebNljnEpGNLdkp8Vl
+yGcraTh1ovAnZ54/btdXZHJ3B4RzECSXwSsnEVf7XZZFG6s+VXxSKyOCMrO5vlJUUplDQ0EgnUN
JMwg37/2LD2PZ6vyavAE0z3BRC1dUIEcoLbeYw3KtjzPl3KvTy+s48pS5Qsob/wFOMeUnL1/Mu2C
tzL92gJWZIRRBsojvF05pJuKQQWEB01QpQITXSf7BKHPzLStzf77ovF9dsxM2b4qFMhSdqIeytEV
ZKP1mOV/+hwZDYExaPcBhIjKw4DTGxM7nvNxYg32vIRZ+RpJcCymIZ8WqE58oaA1nD/O7HVVWZC+
9Iv4VQjXNxlm3eglFkOyPJzc6Cc5ZPmFwPB6ubVTdxz2hgwWMhGT+X76vwbEJGAbYQJxJTwlDFQF
vqEvLfUy3xxLZo3WY43dj3kR81MQQ61FciIOchQ7mxvt+riPyvfk5Dsh3sNVrRkth2TnsGuVIHHH
HO1XVKt9N2bp07CtU1CsvEN94yAroHVdCbXipCAn/kFuJfLOse9e5Cejo/E77o/JfSPCqIreIxn8
6wQq8g0OmFnUu9eXP5UbtczwoS26nnj49eepstoh8zPTs/aU1xXFg4xmWlXybL33LjVffMnMHnIE
mbUqSVOlEFDMaHkKr8UKusi1sVgO70i7tI98e43FiTxRQmDCejwoGpkOwurSLbCmeK9hoVa3X39c
kK+ZSbCl92REZxhU8K7s9PbIv38UeuA0RuxGy1dbfeT7ed5+FTC8tRp3GsOSdR8JSrYbDfvopEbS
qg3A4I2sqcnt1wpVk396yGDuDKy9Wn94Ow/laN7B5D41RJgiQg3dJn/QzaJuX45axER4Eqtl1HLa
z+rKbi2kpM6B/te+icWCxmAlLH8LEqFrujAh9PbcTQqUuJe2wWiXu+efPAXplIpbYwGlJokagx+I
6/PeXzrBt7Ztakc+NYneyr/x/FjtIq8v98Grqx94GsDk9FUQAKzVruAFLDUnhjzfGmHc9nLNMAdi
JFVQFUG0shjiko94nFt950BAAaQnxH2OUL9kWgEkKuPrzm8jmFCb0S01P9SslwcJ/eua+jId14y+
IQ1KPiahUU1/ek25uvJ9+L86mM/DzyVzJzgWKk5BrCjWtRays/rMsP9zAn0YZU0NdfkgUGXmeq9K
4bWcqP6h4iXlpaeK0nY8LQE/HcEopBXVfEAr6SEtpi3AanVW5u/WAQHwO2X/avgjhDlQI1E4cI65
js4A3CLfVKaaiHVH42dZGxAYSDkp0NW6FV5JJ8FIGubkQwYwuSTReT9wH1WaWSrJyA3G76yHSSy3
YxVDffG0xUB6zlc6ZOi8nWbSROnceS1BMOelxlrlovbkFpsWdzGfuqoROIGd/4MHJiflnE1UdeKo
NaqmfD16ym5YioDPjKUW6w8i1VvV5RoR7GLYS9OVoDQeYqX1r3bTxxKbiWbxlOnAwQts0gWFOBKt
wKe35zABLsDaEeV5B9fuk8f5xyih/LRkfT6g5jE0efRdixeAWwYpf7Xm/p5MlqW++iqL1PDJiEJJ
+2qi0ny52R/W6fOIMV7FaUmzCcmRq7Hs8Iz0Y+VByhb/wNMBYJ2R0d9oER6m+PyluZ8yvqgUCPGA
jWlmSE08t7kUJeXoBmXja001YKNHbF+mTlhT/MKR98y4+pI6WTfnhIlkvqGQWUMp0eqNuH6ihEfM
VxABukm5Va80267X3/MWDvXw8Cj0BiiLIV/dDwVY4bonqBrip+Q4St7P1y27UiOtI8r/8tJnoYix
nI4493vdFrttn9YfmU2ugcTcdyB4dqGBhs7yysOvWRQUgDSEvrzK0Q2lefkInQY+RrrVfXUTsdgg
1HzQDOUrsarTCfljfPG0t0ossjoQXho4OeVE9pTG7st9ZgVjtivuiVWg3Et9zTjRsYfrB3w43Xid
BZ27pehvZj1Isa6ufSmz1AedqJAv2ozTZcSsngT6kfbOatJX6uxkvit6zuU4ZbmvseVX0Lt+4VKz
f+IkGrIwO4SE6uBhuZq1gybu05ntPJgMbOJ0Dc5rfFYSTX+AVgZe2a9qzsJO+kZVCMk7/7sRrtbe
0xyFUcirxS7ncWObd3xxwdCVdxOrQfRhjxLfn1TOniT8HgiDsTXJzuu2aCtspD1sWwIPO0k3itlc
5p0tGyYocO6LefozTkh3aLC+vVH9LpfviwPaezOwOOKbTMkVYthxSYPIxagqGTxi891QS6wsEFMH
IWIPVY4ysE4dm7ezWwwl9znVsqZlkvXwKy6RN1jIt6kRMAdnB8R6+je5/Tj1DAMUi3qldysd5tz6
P3GtxT6lHf/mB9lKpkcWRkGJ3TClSnQxpjB9SFG8atCZQhAYii7M92H8u6hF/MB1XQT+mbEqaOiv
Mcc9T4fHf3HCs+G25E0NBlBbrFWf/emXXfMNTZay55GscW9ebineIbpLxyh3nbxe9rko0MWJAReM
sJ7ZvdGhyODyiuerVU4khaYMGHFVuNn4PVy51LVxf8jvlu9gCOKwbc667VthLUKZCeqfgf60CY9t
+3Id87wsAPb9K5B41FzqfbyXbTVAmcrqBRpAr/deTLlI0MUERfCvl4+4ebUsqXTSFtaWLZZxbtZF
tJrdflUFJtRMGBpyRpG0lk3Mix6YXqbeAiSlcEWT/AbHn3PkwJP0QskgrwZ3GHyATPMyJ3KK19Y1
fNkjo4AUSyXoXZRalRLjrUzTY0/Q3ajnE4kMKDbkqOCe9rEhVjHS6tnM0HAd9H2rrniWy+26FTpY
erlU6J2cVbSxDZKAjQln+iEjTbU5py4hg6FpSc3oK7kDVwky1tyiLL3Teb9kHlP8oJrYJH0Wv8mp
rVbQAgKpTtTglIc2wc/c2kWKYed7Q0uALq6PV0uEon0DUTu2bB3kRce09WW7YoTiuj2QFOeAV8K5
dGmnC7JrjRYGuFWXh4rHegncUYyK/Smda05E5ylsgrnSh0QK2Kqv6q6w/ZIkKMbimIa9Sa6fEnCU
wQs/5RZZVfDyc52yPgIu1sWUrgMY7vVFUjSgGhkZ8DWfu2/YGqClToJaS9aL3F8txPX3hXXY9QFj
Pdl7p3YaJgEy1rd/qMdDUKDXWywJlaHdJPRpaV+7VEsaQjVk/tKdM7UmjwP7ueqBvX3ZQdM/H0no
AM3RuTsfLhlAt6Ibiav2pobEoMjnTpM8TGDl3H/Ek2J/pM78x64gYPf6cshd8OnwlZuklFPQ2esa
k4tlz3aNsJX46RPW3bAhoYzvMxyvKv+wPCRRzMfKleRreREF9n3Xzu2G42Mr/ywPAcTaL4u34YBp
hPJnVzCE/rTsi4dRp9ExK8/pprD40sygxXi8ODrucNsmgCqKagnOL+r5jsU5vhlXNgc28X/lqnJf
bVM1cYjy5SpsPO4Num2TIb577e02YfT4SitZQdFcs7v5ifC6wigqSI60dySjq8fj6ZoNsHJ55USg
nSk7eNCHuCTwbyYTT7nmryDicx9MrChmQ+qSRaxcGv+1hFaGMN2Nrwybmq37MYcRAg8ifCYOZZ8o
ySK+1rLQ0DxisShphppES7vweDVPTEdS1Z57Cqfq6tl5eunAWFmL92DlKGZYPHm5ZAvgay5rDJcl
9CFk+4j9SlejArnXknajMYKGIJ82MutA6m9kHnnZIHHYH+YOM9HAI5DF3LpI+u3CVDxCovnTFx7J
g07nyYEm6AMkXcxRqNTIJjyQxurs6LcPoy73Z/mOnistmxrTpyr79JBAtmmF/khwpo5yKwaWw+5J
3umSGtjgpZbP1UR2p1QfrSq+0SDkyBPuQItH7zM7s+Joknvkhm3EUZFjPHeavTNmA5WvDQq/Axe2
3cSm5QMnu1+iiAU0+kWRefVy5M/OwuwGaTUMtn5T51/ePOtU8FO2CSLobibgtW5FOIDEtq5dgV0b
vm1YbEOFnIcrjyZo8NWjke7u2RyHAXO6zU4bU9FpC4upduKxOtn4YEqp64q7NPrNnJLCX/GdC/Kg
i4ca5kOk7AUbbzuVZDyYvukF6FwoBuN/Whw8OD1BheSH70FWFufGLbcBFsRQveTbdwdQJL0QptEV
CRGL7KyJfQSrrmOTrdUj76SqyluXq4cD7liVe1YBUzXOJ15R3ugSbEgw7q8/GLma+BgWYIj4ZFwC
p+b4swcBKYrmXZIF9WWeAlZJXjieQX95rA0jzNGL4fnsdB9F3i4AAg7tQgRW/ucp/NEB42K6wvUl
L49Fw9GQ9LKCkB1VmjBMAqbUXxccaDCKc6jGLZiVNr9JbW6oArdlXyP4kIvPP4v4IrGuIoRNMQHS
Js5o9N9WV5yzjCxzoUVE7R5ue6gZY4gjsYYnRG/UeX2hHq+GutZaMzIFEBf1yzkwyYVs170snggu
gQX0j1eTsgIMxxJMgVUy9Zx7RiH23Ekr4yj9Hjuk5toW2K7yzB5OiLgqysmLvMRVTi75m0bWJkNc
pVDpjacUydx0NYrgcRKFsfWVpGQmhvR2c6SJ86VS18FA56FXiMEUQM641qxDEx7HxhNnAFFMcftn
NeSgAXNRivzaS9wGzOiEbcOaPQe3ZNjYHp5kwOlcI6OIE10sOhHZYQ0/kLrIaCqeygnXkt+uzGSe
Mws3Ts2Erm06xkruhiKXlK4aExPt5W3K9cJVlJHKSN5CqmEEzIIvyYC3yCBIpr+PRlAWigkxqFdS
SdmTvSE++eUgxNyyeLmOZbBYNu49iQRMK9vEYGOD8CS6Gg8a1hd1CQE6DL62jW51shxyXUJS/CUc
t+/hM07sOZj1Eu2DJWCYqb8GozPSr11rrqhWAOdwsQRrgIr2u4TA/wM2lSZHw3s7L3fLi18Wlx3a
PlGeBRRMK0ZFzp4RxNdj2bw34Y3G0tW9swauABFSXmAQupbXADFvON8b4hRoHBUP5FH8mzVtW334
1rEkR4CVsaeJgc5p8ONJuUaNNUbIstHbd7NqSh95BYEbfymRY/dsXZhi80abkSR+qO94i44GXyPA
7Yurhld/Iu8XAistJejxRp8ol4Y0r2GQVAndhHTHAiOYleD6agjVTm/8bl/q7Ck4aOJjW8RAaZLQ
jpiS/OWPGsBO1xm8ubm911XyEL7j0+JY9fZwPfidap843FBZJDeQOPLzxrIQgmH7xsz5YgFxJrht
JDgqpm2skM7ReNqS/SGGGnUpxASDEoz8mluH/qkC8ZOAEsLd0VYMXHQB88M1dRpdeKgtQKePtG/C
DzmRVagENFFFaZDwTu0rttzeiWQVHYgfoM8G6ELJ6UGv02D7oPLScV8+6uxdW8c/XjHdXQL0oSOj
lkGCrm3vhbN7ioj8318qk1DJO6epVIQ9350zgsVL+TzD82n29xLBA7WKFi/gv03rrA806BrPZfUc
arLPNjm3CRem1R4DaSXrsx9BoEiYPlRgd3GCHJfINYraVr9vfqqEzko9osDfIvLHs01pX04hnxMq
muccisB+z/5sjyVSWlEfIRcehA3Apm0xaD4iX7OlMyzBRdD2yLgMC/z6HCcyEoMhr1G9Ty89ylTj
aFtcWFnkZBOLKqDaosOKhelRjDMNNlcqfbF7ycXZU3ny4KnwIGLYZQCTd2s9JOpbA9GcVhhKvZPN
ucSAaPVqz/67hSBwqAM43whUeP/Uf18eTJUag4wEfONYVj0N2jbtDx4Rw+NqELDV1EJAPZpqnA5g
8UOO9s6zL/ep/hBJn+LuwORIXHSdJTT84TJDrlgF6qz4K127A7wYVtHlFaePXWdZCtNN9vAQQpyU
zmMsEJUJyF7k1RKfXZX5cLhDUfUPO9SPbajao951sQpknP+BtLApyRcLdsx+E4nhlLS8VA8sA393
ecxUtXgkd9bEBcWWWhu553PcSGH9IGQLAJtzb94avLKd0fzPkhBfE88FOsoc/Mx1K8wt+U5Wu8mP
GNu4XMA76KwJZV99mChpS8XjTjtZVzQJalX9EcJuStNY+GX1eM0LrME1eY90L4j4bbipN9Ohe6os
4z619zKbkcw14Q3jMY/8vAyglpEE+F0qJv1IoqfRd4irpKkfD2gEe7OBCa03jX6KH2SUbmIdEgO9
kz1aO3+rKakcpuJ2UcXI1bS2XO1wfd1uSyPkjnDgBtkMW57oR4EqEfNqFyiKrkSVPNz77M7/MQtp
u49H/Wjkph3nx8R0J+KGgd1d9yDrW84aIPa+2f6lgkR2MeH+UUuHjOkDlPuRc4+6IzAsZj6P3VvF
2ywkN7jjVOUiNen94rwEVBkowFBC5O8Q7IVKIBjpLvSxFlEmnwOe/5xI8bTLNCeaC264bauFOczx
R56368ODW/fg8IZ9suRBoICKNhdfjFHDqKkrkpWhVKkUh+VD51Hc9dGl10OfP6Qt0hJE1kmBcuOH
A+YqgQCjAiH+WMs8gVWL+XWxufcMyuvdg0HAkAadrbMGw78zJPK5L/0dP5T75pYye3PLPI6EvnIG
s0Dhlk3lP54q82CtL2vKatGiHrHUQpRQSvWes+6bQpPPn50tCCbyK/IhY6ozeFo9n+tU/DJ0IoaH
0wSJQrv8zrWSzmGa081zDI2LhMk6dxxk23+dMPfee2dbHpzgAKI5TUca6wYema/dKnqpYV/FepXM
fXxZ9VGOb3n//lzLai1+9BjtlUz4HBHnLNsNALvl+NdV6TlW4SNiB/rmuC6sqDq5i12dXPi5LAgr
2LqaDEPuI/v62usYGcOxPoLOfjfgZxEv+TvKBfB2HvEFzAdHogIYo1l0q+bpcazQmtZQzR642Vga
60oM3ljWPMvb/a1klDqGRFg/0yfxzRqpWRWdrTr+PHuzEMpcbx58LSxcsIPFjAFq9CF147tJBxsU
85put6iTvoXxywbCCKmgW+YTmGDwn7TC+zlpulCvjIUPGug2yhIFRlIic0438NnX34sA0S+tYRCU
CNTm/q9LxfKkquYRCu+KkP/Amcjege2l/lqTbwCGlQh0pCqjIlHpgFzj/HoKzdnHNvKeLQL0IRpc
pnXrEi2LkbQ/VmW2OF7kHZJIz6R2N2pmG/+uq7wUwM6s30zMkL6f/iR3qrCq8ej7yOsfnCDyzDye
j091r+sBYyCcXiLki8m3ogZ+qFxcxz8DtS1n06YwqSsOZ9du3wcQ9OldoKT1Rb4cUQ9EpB+VQB8z
XX3XuHtdx3IdhplBhVku2pbl308htfTk/kJ97qaiTo5mJTDmjTsY31BYYVLheOrKOBO0Wm6bCrTG
M9S0/GrBqiOWzRXEITdV2blCIufA+EBnu7aGbSaG3Do15iVPVhZNyJJwncMkD+iQtS/vizeDAAcA
IyK2BBYHw4h3zG0nYgRfqhlyH8ameph9ZW44wk5z6ndoJ0Z0CVvRO9YjuwO8DqUBTQUOOMMqCtQc
83AX5l0S1sfsqWaZBHpAXkZpe34w3dHVrO7LSkoSinUWoQ5n6tbNohjPdta5v0LbkKo9fcS6JnnL
PnVIwd36e8VlxSZp1MHvlh7mvRIXzlwlnA8lYaNc7vuhdlJf6GHWkHSO1nGxNV3a0MjW9izPj0i0
KuCeBz32V4XRWD5ZJwLYp3zj4okmrWt/mnwM+kKrfRsswYi3kah2c8FbXoLVt+E67uFoMWv7CiJu
PtCKTQIDhTlJOpMB0XfHAzXonwUGWujICfhDMYKo3XdIXxqwZpK7JrsmmMiQms2UwuAb1uE/swMH
u1L85Gmw0Azfy0pgwSzcE/NCJasemn0tA6IjeUH2S2ncV5fMOfkblueBqo+NikvV2NdH7e8DVGmu
D4ooM0sHPTi7jtGbx7RtbDX/EJ/Y0pxJv+7+lrsiQpa/nF4eGRi41JnUOgpHu40Rdo402eu+XE3R
nvzoWSJgcOk9FZ6D0MNrBTkGLyViEZd9AfCJJSgz7izVefadNzeDC+jdYGKVUnPoIS60GOpiM0zM
264a3yTZY67ap27kQaxhB11DLTKr74ncT7yonR5WRV1jVu8Eh69DRMBa1Swc2KsSmSbfrD5UzeYi
M41ADzqDFUrJdjQFrtGjJYXeIvyWjWIWJg0+IDLKEyHBXzeQlzFhyyva8E3Wl00BQdtIEX8d/+Ld
5si0yqJ01mKzuCeKkquPAcz1DvtjlVVeRUkctoGl072qs9qiajWbJMm5ACos3mHsEhNgIDwnCIkr
7+PSnXK0nCJN/XzQAjqoZNaC9S30rRrdHeW3SGHX1Z1rRqbOm6jy9shSXd6jj/ho4+u7f0HXCnbj
3oRKVDoEMXmtn4lhbyQXyGhir0mjwzWtTriHk1jGHUhv9dhvkTpTlJB2dxYloBIUUHg0mK0NXvLm
/hJ595siyCTHCVCW6Aw6SlxZFl+SFEosr7rHKYd+q8v7xkaLaaPeNiEZXT5VOiFmn+Q7ni1wnH5m
Km4X2bIc5z9PNFC79ri3aGXyY0S7IRjU/zeevJ5L0OwVdKdjttlcZxd8XlstDk93CUbrOHxrS0nB
vdTZbV6y2Yas0IakArsan2gQiD0N/mV+ED19U3aFAIh5I/wA0pO3F1g6kRZkSioPEJaeAUElLSzC
j/vQxnwz3s96kohEY+uKkaU22YzCrx8uWuep1If4td/Pk4BF0sgvHLidZBQ2liYrGhG13E7BCNMW
HOuPcrxYk+2VbgtfVxJkz+kOyV6WSdwBcI0IRkbfEXn2wM7EVAzqdAsRFGCo+Rhm0x+k8Tctgk/j
6BtuqCOjwcFj4u7hjQiRc9bNwPxlLwVqqSJtt860DxS+yz71Za6a/VvgSuaf2FCAEgCU2SLTuTj0
YMt0WfT2EkhgAPoRi3jpdKjtSyHXrfSeGHYcn+3NYrh9FEIDCWeFzlUSvXohc61gXu5M+5dZ1AaV
HO8EBbWsbV8p1EZzItodO4tJlN5Cl7aHeKnd0JyPhe+4/G09zQJNuIZjSsZOjKQ0gveU4Y7D6dav
RvFl6RS2vOThwNubqrIucDIMYEHKnUu+lgtfw2MEnEGZQNeE3LhgeGb87KjzsrNHxdq7d6AGHQhG
uB6cgPOGjlByWukj5d2hKVG27Wh9YQBvPuDSwehsqGQimPc3NpDWPJdtkInUqR8lH2Vs4deCOSB5
aw/W4uK4SwTBBJMKPup+DeS4cgcGCkaRUegnStPk4p2/UsuIyr2xuBRNcqf8osAWPFbEBUKydqH6
iztquRR2JPVceL1++wH+4MxhHHP8kBWeUcF+URCH0HUSKaudtT1gfVziriuKxDnt2op56mhcX0Zh
lwmll7m61QkZrzr+T3TT0GcKq6W/JwmRbUmtnGgGKSQZuNwDvRaXh7YVkc6NT446wuNnbq0Nx4cZ
h4w7UDnFLhpXPRHIVplc9Ty4tHdWXycGQCTbJZNERTwc7fMnpicdW3cPdo1RNHiqgH+VTTAkf/jY
A2oumkw5U07tXfZupNskSS88z3/WkvqLx43cByHe/pSfz9or/D5jvbI6gaTSIbrc9DSnYi7fZyEy
Q4FjgaLEM0ue/Q9EBxlhfgwnzOvs7KcGpE89pPMpG+jyn0Bt+D9IO0LPwtkBH2jcNDDXB/LQSosd
OHsrbl5jcIHSv6jVLIR86eudm2qcAXmIyZHFPuVkxSZ6mD+Eym60T9MZMZWAors0/c2tZCf/INSw
E0pWB0KSIVRqZ/KMw/oI2aLfx+KXa/5hKIjJuUfDLb1CtDi0PUkLEukPGKypmtp6frpS/dEe+xp6
Qy42fcuQb0uu3vPGUE/FOSpj4EA3sm+xJA491PRUANF1DefWzaasX7SQtECmT16k3tiN8gKcJE4Z
0r4vvutUN8eElkoBPbVKqLAlOknrJSBFD0zcj8ENZkjtgEqEjc25/iA4rmqd5Q8PQ4W66o+QLW/a
XWGgcZKvA44eZKfaA4jKepPS7Nr6L0ZbLTBL92LLHES8LuhtxSoE9HzZ9mk8iajk64cIAcamhhIH
iNfs4IYX4mKEyuqBzijO0nXc59RowUoeOG0jI+3NUEEkBOaO6I+mbH5frXHXP7bNvdcieBesXyOY
l0V50qJi8htEK2zv0Vm6lPPCRdTEOzil71SY3RZRwuNM/tYjSiAmO6v5KFSXgrEnolkoD++dV2rA
mRl8TqN8d3F7R1vNQITqx9/VXgLxlVrcof31+DxUhE2PaAHrah1cRcTb5t4WIGI6F3ridpTqE3IR
5qlvsGa0AVvoj4wj5h/rtyyMzfKqOEUGb9wSIQKtIAOb3oqGzyeU4OYEVvHzYj34+YC22Wz0yx+n
mnzE7yU5vp1G9ppjZH25R+FeOMIUwJXVpaMFMRBc9LmmJuoI7X+zzcQbPmlL4bBvaYfO4pbssjQD
+8BT0wjG11i+wB5vYAX1vQso7ujA4VfDhxqfc8ihf/yOSue1QcYkt7pOlxw1Mg9CfaMDc8r8iCLO
zfBFzKLr/9pxCDa0eCmnxdKp3eB33NcmqovJ+WRlcFJm0Kd237oHBr+R3uy6RrY3I87Er7srkjzx
wHnvzLw+TfVY5hXB6Sq9wy3NeDAbchzdJN1bMMd3dERNtSxYOPeRBFtYD4hVJqDNZ2r2IHCv1QS0
V/ex9K+urfGPoL/tWHBD6v2FXdQwXu1Lrdp+0Bg2+sQ2gpNIqk4Sfr+ChyaK66umdzlaTi4ivIvT
cE6H5iniS+O2qHi76v2F2Rzr3A6Xy9NMaRGZo0ZO+VJg+t0ijApeNKpAw6+jhBBiAq1o2FRkfJKQ
coW5MFzL0qKocMsrO4/lj7BMiJS9BYwMzOLeAHH8uqXLrcYxCwHYrezhT9IKzmqOAXDz/+n4BKtW
d8nwT9EgCBKuXEqjjs4bhjrgzc4fkVHm72pFRbmV3v+Y5ZzHJ4Sr/GA+3wMTqpaoDbZIZ5WP0QJ6
sbv9TmeLM2RIZ+xPFM4gL5hyetN9otZBkib3JQnBxTixhWygS5RMnVy2LUC2Q6Wp6Pt0nlxypwYC
PhlqbRdsJgb8WAjpcWoWfb8QPG0XxX6NzbqVvLP5HZGSDVvYM4Hc7Lv+r8fhV6KavQhvJWjK5V5J
04dFH+O1ilQLhaGYZsQjPVF+n2QwyiNZ7Fp/UZXQRVGNFDQOiPvQu4E0PI3sWnEBO2pjqBxQD3pW
CfLRmOsGe5MZWA0qfBl/ber21sN90BxTrHPZxjcw9pHI2y2Z8iWQ8rUS0vWqHvCEIPJ9CJv7oPQh
KRrs/Ppvcu8BcMhBFZcJDhP7o6va+ympTToIQtekwdQPMvLjDz/wOc7LzpKYPlaqrpnJwvKEf4xA
5v2r/lMC4JT7k7bCiGueW2MWL8MRcvN0Q+QtQXPbqOg3lAHN3vkHquC/TIdCfjpUioEX4bsFPuQP
43NdIf1e+tgHKdM4CtSkzWtRvaqyYMjdpXcu1e1vjkh5+xhCEPMrQd4jZA+96IVyoh+hoAG4+Gpc
A81Bx1mfPYqYoJwvwOML0yEblS3Rqj5L9cwlNDdiJ75DhIMX8yf6BnhDK63032sg9KvXxX5HgNuW
czIKcW7dz8eIln1kmDGkiBDJT4ptAq1aIQon4IbIn7CMUvvylnq17ee3JZcVIvS7PZHYth4yZWbP
B+J0mQhTA4AneXUS+RgFf+TkInweD/CeC+CftrlAqEBlCxwGd/jVQGNx9KOWuzZ83npfbHTXd/Ra
IY3pkWHDBQq2MIeXC6DqWqmOdawKNtEjQicLEmvS3Fp9orqL6rmkrhQ4FYgCOmgCHBR/VyUX14Cp
kiiJ6jn+eRwhAmzow64KEJLstDGte6VKWty9L+e0j9/UVknSxccphmsxKPfNzCxBFA95jzT6OCie
3yWCbTx8s9E79sb0Q6g8Phhc5wnkFvJGS6aILcaFVWH7FJIWhazt75DwiydiMhfugk4ibEBiPiYO
YIAzZuNckE0zyEJtmkavort3kvE+92TV/56L32ongZHI/kbvcduyE6uJ3Q9iarKGu3LJLvFokmfl
RMEjoh4ZV9N+Ec4cDm+1tEpQSzj5Bj5657asQOA2CFHfySq0vaHzJrvzOZcljTSfB3JJWwslOoQD
9268VocUJVwcI8aPHvYKGXvl8tyH5FkltmIPDcM2V0iwhaFNHnbZxQRWU4ZK16kPzNa3VP7uVtmv
lHHIMsoml9+zbuv+AP4BAT8ZRMkysocdDgLLgny0t8qu4hR5pZv4Tpr2Udf2OTFWesQsLvYIVtV3
WrAfiqq3CVPVn/tE5XMu2y9xHTrLxqVpGvTIU3ZXqrveqoVyNvrUqZTqJgPb8+2ujv9BD70kmQGv
dhrgtvnbXUPHayh2+S6jyzqXCMVTWDnmwaGsob/Jd7Wsp5whW9iQS2nlBTkOam/L2GAzMIKRG754
oKMspSEe2L8W2OcdbKKefxROzSBa27rWBZZHVC9/sRzKML7xVNbY9EGP5SVmNc0yxVPNwQsZdTy4
/YNwW5egT9kuotMLJt/LqVdcA2bUDdUJQmSX2ywET3uresv9fNDLd8pqAoWHaJOjbl/+9ymH6cDj
BcZPoGgbe9+cAv57BqZclaItJm7v9hqHFz9/o3sNhIYf/IgNJRwaI4gaW7uEdszeO0CZ8GTsw8/0
mcvDB9BFcOg9Gw3TNCrs6D1I81MHjgJOFGwVHjo4sXQunQzq/9PDIk3wky+5fvkdWl1F5DjXydZa
DmoI8FWNhGt0ewDtjKTDkKhcvXIhQzBg0zk2VKd3VdZONWjyicyyIu0amIrUSetQ4NZt8kdbN9/T
PO3R0zjdi8y09kS4VutNbgP1BgU5WC9IQn88Wzcrc3PCMv40HT7phN2IZoI/Md22F5DbAOQSIdF4
Rj1w88p88EtzB0J5bTzfGFPip3EXNceQyKl7onjubpcb6Ncl1XpuoSMtcj+dhgKD0/KVBGAupdGN
9BFbXumWpGXWoZL2Jfm9vgUittZ+dluyA6djYAhb78GDh0DXcVF4wO+3LzM8SxG2ggECeQJ8PjnP
OOT3Lrs0Ofhl5wqNoQ240L3gYwx+M5h3A45ejoYxghCNC74irkD17FnJFDhW44HuB3x9V88t59sH
VJQ9fQ+uMb505gjsJJLqL3r1KL/citSIg1UbuSs4uEqg69an8vZm/xxnpFFMMHy4/gqyshT0XGHf
7CUiPYr37bs/Dxznz4eQZyfIRro45KUAyKY9a9rBcewxJY3GcxNCoD+JHbALGPk6NvEvfx+yc/Jh
PjSYvHO0kJKWaW2QTHZXRPrR91BWrRBFr6O8MSqJfs8I3Nf1qHKJzCufOLmDU/aNISQmXg0ORmL7
E4Ps4HFnMsvDwOSrvj30mNnaD2oC6umYutNtYgWAvc9+zMe0laLKi+lt3QNcZ/sxEsB7NgQtiFS2
Fm6J/IM7kITeKN9IRV5lp/8tyAJz2QzWF4gxMFAlBvaiH2BkNX5fpno97Atdo7CHgNSm/VH6Vmku
w0ixgYMiJ37qttNUN9OtnipXt7VLJm42zDiuTU3+gD+V4HeRnhYGSJ56C/ShbnEeMcgtyzvHkfQe
+y8m1eZH7jgvWNjV2cJHB0ZxR6x0JYV27NVDeobZI7IrJBRAUmryE1i4i7bj0TtHqY+PN86JDGc3
ZQ6lO9L+fyDFyKLI3ib60OfAbXfXlp2hLWsLrEuhFi2xzAdsYAXP/8RSxxcHL+B97kP4krqbvE/Z
SX3B1aeNnmxjD5Kx3x0wUAJMPsvSL/aqir5ELWQjvE7k8PVF2bbH0vWj0EID7Q0gwXzI4E7I8swx
KO/I+Rc3smQPHkKAarfEoo0+kegtuT6qqRCRrJp6nfu7XSGFgkfR0Gss1HpqqW8kYTJYSHQldEmd
6TXQ3n380QjzcPL1dMEkKSlfqPDkiL8bqlHbr7qIiyo3Ao2n2kH7ssRCKt6fITy3avan12/YIdBK
ccggjLOcnOTCLnYn8OhSELYzwfcWDM+mE3qeMDsbOGcCcwVmHgUmJPNeYOEQc0Jtwo15sbtPO0Vt
kOhBlL3QKITdsHQax7cLS5zPm9caJ44ISkBoJm0u1PfNRJf75xjUbGkbNYL6b2igCotsRHuTjXu2
SMaqP6FQmSQ0cilOpK+7Txg0Uk7eD9JzOu4XWCI3ohLiZkXjKxvPvOgCPT/2Dd9Z+hHxleTWFrlO
ytKVKtXXrZuhp0GaYHbWi0LjljjMWx6n3Zyfjh9zXf2hk3wY+Uuf7YsMZWT+6RClVxpxeFJqHfGZ
WuqOlR0pc1VJLVnnKPQB48X2IJYFjS/VrcNH5ERqejrt1HfFigR45fzE5AL+aLn/D578vybh8YMs
OMggM78dYWYh5hupfz5Nbfiodf3X0k52GpEUCIXhGdT1TFgVy4HltCJYi5KJxLtHcTtAr3l+wKdG
eHADZY5Cm8r9LqUh2z4P66heZGhlwWkwgACuI6BSfhOb7enPsMNrCQln1GRuSbvRjSAj4fEkIe6S
TpeUWZ2ufUwT7lZUwDy8ZPZCAltJTT+818rtndlEFSJ7zN+DbHSQpCP1thiU4Yat83bY2DAh8UUp
JTQLQIoRdwd/Li48/Na4JVkx9DIm539xe1Ze7puKl460fR/YOModqS2+IQ7M6CB1KV4PuT+madVI
qSsRiPGLNiMbiPfF52lV5u4Jo7AHvgAFzqfFyn/4JEbnM4ZscIQCgnqIKuSi/rprWs4goCfyYJRf
uwVnGyuesgj1EfI2Xdp5UyAJ6jJGPshTI3bpqf3bCcqRc+SeHZ9PJKVsuLLFrnXhtVyZcv3vCgqz
TbQxgLlF7i5Cn7ph3SjG7CC2C6LxF5lUmGp1Nx3mkpeZGyRLvpsmG8uttUms2M7K7NU4WhPzXOO0
2KExN018iXJaKboYbIeBh1To+8ub0xmBho3fTG6rn6RwyJplpd3mXIUqJRAm8uYT4vTWpM2MtbHC
pK2U1GtJGkR3RdH2dHqIfCDKe8pgA/PB6URGKZssl6PqEHn3NQmTO5nJPU1q8o6dkQzO/42l0Dx/
jQAGFlgVxy/ivfpFrwt26WOLOKUWRD2CKLVUvKtQdtLAWMe5w8RA5Vc/htE2OY5C9UFyIE1nuLN7
Oh9LCn46ZWIEshoEU174JQTNJQ/d+JHBAvYuTV098oRWHpeJ222WK9PPxLwkuoi/pRUQ6LggT5vO
uguV4m221faV56Z3CsHTfx8ifcW3FuBRuG+L0NC2B1z9QBhROMTXtPyo0EuPvaPusi+ueENd53iJ
stza1WOIyrTLNQ6GmtGewUVqG1eLpMsdeID3oRrpaD90M0Gmfkz4drc/HyJJXBQTcS9Xtbrxnedb
FrKG8Qt2ZpP47L8nFCmN+4V+ZSP59iwZQJsxf5zdu/nFLVbUNOa3mXogr78odJep32ggth3/wdmm
oE4s8+K2o7GxK/56I1QWwDcrgR89Z7vqC9PXao1qnabjV3zVuU3tFniiPBP0rBwC5JIEHZs20Acd
WvQw5ey8gpLA81IcbgJvqpYf0hXo0trLR5+ga7aImmoBNtHif/Namk0vGhZU/emrwaq8G7/qfrBU
IxgVwtcyl3zudLyZbMH9D3soJUWPpaYPfjVbc8iVOtsVbPUGpezqo0KacqKJD/r7wuvbbVHhTPIK
f47rVkE7Fy/jy7iPdwvjzXXYYkqTMAWa6c/z7V8poW9j5ib3S/aE+TtoHz2GD+bOPUQuJgeQqUzX
dAhb4DjZX0WhEajq+dxTzJZJ+Lt8JSSB40fWACk3HtZ22i55BD8hcgUi/V9Uy3ivjPWfhIMp01HE
kzyS14P9qC82FQg5bPlOKCdreAT5quQLB0OMLld7t9uPgK3TWZ3m4amlrTPA3IAPLcjekQz4Lz7q
bE8cttSveX8gsHOVFqY6MfbSr9HVXzbVvytsLE4aP38KEtXR/aDXTK7cEObYT+Mv07j+HJL6xFdT
JjIYN5/aHEGXWh6HJudCKclPTPxEEWnNAGIopRVqTMZeWGXFfQP92vnp/mr45XrKIyQcar1mneoA
wBbUm0c+GxDaAOg6nY4FQo8eGdoND7stjU+D6QYjo1prIZ1rrtuC/sVCvbaEdVi9Ck3kE2xkUdMw
KOqO1SI076SqvLy46jpAGIt8n3BZCOlwQn0SNXS9LIXN7n8cynbPItaXej3m/e3nhY4UMbIsz5bd
xAL/9fL8xiT5y9/NEilKqjqpMyS7PunrWPlINhAnYi13bssedz2Vg+vh9j7xfcfr6MHJAsx3eVgn
2Fugpv1nsTIrtE9CUkvmoHeR/2CBCtd0EsA3CVxDKcLKwBU/wpxWEHXfJw0Q4bPDRd9d6GnrvBme
+9bHRnFedLjeFKJhFvFR8FHPp8G7nNZ+xtFCFa5CHKPsatQxdL2laTwUoXk+JpB3aPvx6WFzSnn6
qcKhmBNNu/4NSzjlDClSwVMLVIrcnE1jTqUGTJ396tHra7+qLsvqPF4LWBFv04IBRiyzHAmuEXkm
0lrUNWSe4gyk26/Ygi4ISCGDZhDoe6JhQEt2e7NJ/Q9AS4HQiJIxsPQPA73NH1HBBnI4vQiN1oe4
V1CDHm1bmZcdC2btyzPfXW/YKk9A/BikA3cCT4Ghl+NbKEhGw4Ny7XyTdqYHnAOye6qvjSU8PvOB
KsUppAUhp+fcd5+RVgULkrDTbdXbUtOUCAQn7Lp3Qyi0knGbA72oAOcpZqAF2iTRXEdXrmpw1PMZ
ekkNL2wZA56Uyg6eL3+q6JcNWOoVvmMnmsDqJHQIAVdPHnDOGacgGgWfLuSdotDE1gl4PcKUSE1V
fcIhtsuovIjQezAFUWSD/41qHESPul4Nw0pS5X6p71rz9jz8l3LNE4T7kao4TiXznKPy/vnmkpI1
/WrHJX03mjMivo1TsEmEXKbQG+apF0QU5W/VCqGCB3Zv1omXn5sZenYTu5rfTLq8k0RH5iRs0fNH
0Iiln84kPjzpWFXcpgQ6tG7EonRGSwONZO2nBIJNg/FwNYSOlnpdgCHK5wfkUiD5XciAG2fUDbRK
fSibcz45KvznTUp0/VR/1VQb5M9dNZ3nF3KalF7hwgtztiXYKUFK1kkX0s8N+arB9jIOk6gApiNZ
oOYoauedo4hWgbhtEd5zuk5qpWrM02ePbD0eOKPEgp1MkBCX5N3Fj0YM7a0C1qDMSbdhqieBx2Lk
708lX5UPwE8VoZ4riP6nhI9r6mATXNkW7XW562DyReCxd7sVfAQJf5eRRFbERaS/S1i4xUgVjrbF
BWs0xyZZnw/b99hSQGomGP20QQ0NxD74ri11JJfaZv9wuzH0DBd2YH3KfKeWqo8r2N2tp0K160DL
eQvmfJK1AmcMkxbCTvC3McAxYOnVhjEguoFUMyeYzwwKDGzMqtMBMJO42skSh/tBRwC9LMCJvBG2
QGx/6MTLa80sFAUJXNJuHr082pSMgZQaunQib9+gRskWeL8TxSFh/FEaDcqZbHm7hxnGMxD5Dmuz
znjw8nUlykKUAVxITPfEfmplhdVqtS1cIA8HxgFSbzLm9XAxXxa3vzdE8c6rG+IVhSpEPHMIvo53
qcHf7GDec4XE47uPFmMofneKExKG4n2EbsWGb2G1qfojOcO1uysZb0XF9BB/2m+xryH3CxUy/t98
kHXbKDNHS12WaxXwFoQjxJ1YhYa33ZWhgXpqX0Q7SFRIO/t28zm+uonJLHCflt9HQr0g9LQRbvmb
8iOw2HYJGE0RPXu1ATuT4ICNAIC4MFYW2WtjAERR/uMMJBeccvNgH1aRzeS29P1Ue1aUJJQJGsZN
XIiMdIJS2St8tyKbZciPQSLyqOfotAMnNfiGA4BRrPda7Rmmt094wHERVPvMgetbmBXEpK4oYFJf
4L+sMDu9RzhQvhTM91AEUzGTs4I6GG79fIvoearyOAjSW+wFW1psmkKWbmkh2uvaMA/TAAcGhu1o
KkPNDpUyIQywCZKocoFBiAP+RQsgaU2T1d5fZnaoJhFkmhXigq7eTr2TUDP3zxI0dCgYYS0bZI00
XUFAlgbiT7OCQqNxim4Hsan/9MJuaGCCQY8t/C+eAREj1piErRrg3gZ6p9uQOBBn9CnSfBJ0kXxr
KtVttM9mfUCPjdMO9B9uw0Ae4YAM+tczgDVwLYS1WUNxTfbLKBYKnTn7P30eU/2kjEY4b1jz7yBo
pimL+QjRdkc/Gj3yKNK+bQjKhc6Kj0ixX9kfGDxKYHB94kbeDqfU1JfjA/Ua821AsNcy4y/HBw6H
7kjA+heAAeS/JZxziThyNRvI2DkFbIroiT4Xf7tWroZIWD9UYJsyu485wvln/XJEqYY3ueFJHCh1
suUgv9ij7EnUKnEJ1FeK836xGtF/7PMS8LH1h2L1r05QuVNABOGnUY0CswzMbikXOJ7h1dRyHwpu
bVOhG8CIHknc1qgL8R1zmfVNK7rZZCbyN0fsiPC+Vl6Rv1ZBc/hjBjUNQcUpnBwhlr8kxaup403N
3CduWWBX+Qwhgc9QqX0QoEHraNgbdLPjE0HlicIZmNVhOspifxf6Wi0s9a8GDfeE578AbAaoXBDf
EM7cS/lQ3AcFLV7whd7M/XnM3bKzI2MYmf7+nKIGSvurtasywU1TsF+OAAr6ShVXEO3aSkbCSRXv
ALY9KCV2MCxoZ6967lRUS9SZz2Ay7vuZGSViDR9i5JkcrgUqvhys4Bq+hERsL9cYB4VUGSTmHnM8
mjC73DpmrXnlhaMM5yNvniCuDoQyP8G3YDT1jhhU/ySO5Vvm7d26e9hCT/r1M2K5VvFZ7mMwXm18
KZhFko7m22ope7SCSBYFb/0g4G7tEvO4UjMWhfhG+uVHYnPqiVdJs262qX5Kmw/E14TBupfJwmXU
bkcNOa40OsDb82g4VbBIcYIqYyxI0Q4S+m1gfKgHyt46WKCVvkYz6OWmVSO29rKq1rg7Pt5mNZes
yLzBExliBCscWRHfpBEpdVVinaap3XalkoPOpeatlznN3J+dq8BMI+/AUIAAPOjvqU1ZY3dPlZug
ZE8k0+TUxRbg1s3n79T6kL30oQOyrSMoT3MKie7spkWu/E/dGVJs0WkRyIiz4LVg7UdQLd9ZyVzx
bWp/kaBrUIFqTT0NdG/mk4l5jYPTTBRPwn9usz+/bYp59IBf2NLzVSpmwMagfga8X4x9wEALT9g0
FQSJpsCPWTZQr3a9yhyY3BsZWOABMN2gPF5qwJqZGWzZXWGKiOvT68kziPjzljZukIRkxT6VWaaQ
uw8sruy0ep1MFnuTnHSRmoliDL4O4B56mj2M+noLEE5HjAoC3dmdiBv5S4AAdXqpHdV3RlWMr/LU
UGquxc9cdKGZmUG5z5YN8wHnUpk4jG9j/K3okg/Kmf7aHVnYhd7ijV/5EAao5vx47l7tsj6jH4QA
gWBLICAJintE8jqNYuULQB9yZeOIqaENSPF4cvPNL7SYOh0blafVqJDeq2cz9LVfZMeW54cIq6g6
M+PjTLok5LsRAod+1IEDc4+LZrcFdfOzHJHhkyckF5WUBcp47acqe1ZujM8wO/JtfE0CYtuCTvE+
qzuMX4lVU1kvaymlyztcOL6vxovBehNk68x4gede2ON6GjoTDHtGYwu8kjr+EOhVzV5VMW8rCkTj
F1Cm7oXnGahIhl0enyHI7J+1YcRrspCu8unLcBbnC6G6hGCI5srU3LHhgmnjfapGYlrfTYHVpZoh
BUt6YwwIBxIpJL5XHRtG8p960AfTk/yFdEyZ7V8wPOok9jSLK5CsPAtJBJ2vyiNe7sKaY0cGkYoj
p8/aQ3mQ8Iy3dJ9TP3VabAyJfEupoyUaKSIKkeSP5nzCiKJrSSeMC0Cn2Ig6NEBQyrJs0wd+MMm3
EvbfzARq7wKX/qWMF2XqqKnbbocToatA3kMhKeCQRYAnfyMBo4py+0w66JdyBvGWsWGl9oNBFWjT
dhLicUms0ovMtBTfP0eLNxKEKsRjVe/WOYaJM87HNCs8h995DEBHfbuKPb4QUv/R9xOGrWmFSmSp
0e2Z1sN46JmACtP9rANmCf5Za2mClxeiiDA/2s88wamW4Qi5nO59DI3Wz4rQ1ZL5y3yLxr5z5oRK
BypEtCvK4QpSXSLMz3UDfSYt6vxvf57D1WuJevZpd6yPywUI5yPYuqerMO3cem9B02ROWimIaXUY
eE1pv0aLCpZX+Gjrcil40l3KZUmuCP1nwfqaEvzbpawwmk6qDrbBUG4dEcP18XM+S9eitUwa+Z9J
wY2zxzbv0bbwA+UqgwjnGvYX955xMWMJqX6xoej4pGrLI5C5hwIXhIetc3ti4eGEI+DDvSCoAJ1a
Ywe6ZE2xsq4+SUHVzN3K0QahWxhBQlAFu3ThVjAbMFLRsrjG8Mz9f0QheDvoVEC0PQjSzoWOZ/x9
9FEdOk0e+g9T5BKKEv2rnUWKjV6jHyCIhFA62JPGtD/tdc61adhpEhkVOUX1xwHLMuW5sAmQGx8c
9Vaw+KjTIsBh2h6XaQZpUKMNGQQhk4SCfAsx3IQJiveO5oBjZcS+0UZiCOqmWCGl33nwiAG3utOX
pA6S0pr4wYDy+4exO0omGh+EjDDtBJFq55TLduJTRr3dlY3K3SNj6eU14HP1mS25p/ciMy/7eADT
yODtB1MDc5rsqgRlKpJvWXubg4uwIyLJxh085R+OsGn6WKjHYN1K2HXpXYF5+GPa9BYKgace5w7d
wkTNUjnrkSC9lwt201nDAcri0KmBEPrbALDxRAv+ksAA2iQADmGmS3z7L+RHgZrtEWFG1gVeUZNK
Pz9qOfVriq/62Lxd6tZk99ILJELBkVRl7aauEYMaJ1RHpsFG9pfvksI9qTPhh7kUCT54IAyqwsrV
+/pka7R1YPcYWfWaWDtah8u+ASYrhmMZuwTGQHY9a443hG/kJJwotiWfLlVZoSU/NVJA+wj5+SPU
QOfpapz5Da4abAYTuxccBDAzoEbJK74sf4ojhXwJRdCwMowVtCATx4s49OIjk5w1Rsp1VqIpfxbM
hBoBr05LWpUA/BpGtaj0zUCyaMQM4FSTIsDVOMTqOoqy49WPSKz03Hx0g4ayTSsYFX/vqa/3FStb
aToiB8t7uANI3E/SlAeO51+3Zhcct9PEePbzGVkPufvfWypeurNzY+QyGZOa49XBoOipjIg67vAV
ZBslvAeX5RkNnCCMSY/9LvNbQQwcNMZASG9MZ8f4Y203BRblxL16pNNZ9r17NbzY1X/rKabYDciS
dp/SMNawyuzvO5bG69Y+VRIfK1XmECFaNlKhWJJUNX7TdbsiymrklHOyMQcLYoZlhSBA/jTp/d6j
yCO2rR0zWMkKlK4ZQYbbw6SuG4moXhU8xG9rwSL+jfgZL4zuOr/goCK45dKr75ZtQ50aeoZowfuq
cBSXM1Np4on0J9o1sR+ymEM3qlnAPw8KdS4dS34JWaoyHpyD99/r/BEvJ916q08DVV1MJfwMtltU
hYInH9mN8MuXsL+M4S2SFKZ5mOjLsXLu6lnUwGtNpS5rPyfoMwx3+aISPT8W4VenkIIOB9Z/yF+f
kw47Qr2c/S/aaeHpHvv2tQj+eYr+DMigi5ZTZ/aVpnOxqvGRsG2VRs+pn2BNEMF8JTX467gbsg2E
DgOLVLcvzPi9k79n7rPoZ2Kj87EDk+g3nTvVPG8en1LZ0xn6NKK7WOvEo5phH1RwR0nfSMb1TzvI
RMgqtfNzESSuP3oV+LahuROzGf65LQntTglBXaAPfYBI8A3kZoaGoiovOQQrR16RSe5F1bBuNnVD
iynBqwujdZMj3UgDDnka2ZPoaW/ZX4Tgw/JOYWzRbGm8dGWde6PSZZXVCTbLm43GtQpwTE1n+aG/
MO0eI8VpurEWvZKlTMZ1WiW9LYHxyO9GKJPnz2snStwer9BtDKLq/8igPhn00bIHSH2TTXmhDpeH
6EXb6NZhTqTl6/JVxwOpXz1At3/VgjO19MG3DCHhbteddeG3eVM1wjkWvXr+rZPOxg/RZRrPlfmE
4lP4POST1rwpGdZgurjwqscCUXAiFWPdZaUIseNxgmmPg5Kj0h4Ug6AHBJRAOw/8ehAhqafpLAim
ucDClrlupEVrocaBYlhyzD0sZb9OMaHS2UGt9UigNDJl0MzU1LUtURXGGAy5MyJTqUOqXU/RnY8Y
zqBTebrXSKUzhNPpy7TIeGIF2yEgKS3ti10g3LY+oMtZLPpeal1zXMxOX0VZ5YqA55vKhKGrGaCS
qNSKnvS4cVhCmDZ4FXtzIH0oDCwdI6jq1Hy7uGpNs65IL3t64yCX0esRXinYGjsBMNFTkonF1Re0
ygv+/UQpP+yAoqLRH5v0ZgFuiukBz3Kwy/JEbCHJDZGNHzxS44Jhm4PnSInQli4qEOYyiMZa069w
Qf0v6S8+WHQf+b9tVSZv1UIZtg1EeYu7Jxqi2VogOyDLYJJLIEI/aLfPUKxzspnOyKEEOGp3w7H8
+hj2Q1lTUAXLqakVsxyNCy2sfNKs96wct7U1GGyOZMsnl2rVc21t09WjhXmWCB9ImCt/48a87fYI
oAfJM7zxDSuSpAZ0ZiaMfsgW6RAXxK92gzxZlN0Pkvt8Y9Eb2m5Dwy58OHyAFPrWNao03qtWNiyp
cE1RkTl13XfZyP3qABfzIh4df09eUgHiNXZerMYUs0Xrtc9Q8FUQoBiQNTodcZlIK1dhL3u7JEWU
yl5rQA5doJ/20HGOsZ2+wziVld+s03abwN1Hx++bvwneyLqJAWR85pnjJJC6Kpol6v8bJktYPaYm
0l4A7vYQHjJTod8kpvnxbsOh1cZPW7/oSfcYAR9Lo0rQ2AGSUF9ENs/3n31B1Go0lD0e4miPLVpX
O8KEL7YZ94ZnOQ9G2DXiz3gR3Y3BfZhD2LoaYBz9rtfoZdEAMQ4DNt9J7x1NMWVxEzWQ0UcSPz8h
leZYkigjUNvrIA3UEiwSFiVX680/SsofCGb24gUNgY4la5FDOLqY7qNhbaS/98gwrxdISPsBM3WI
3tk+8eXgu5DqNlLqXMT82vlfpJucCHzBReyV9Q2YlTwEhA1fl5bs7UNSlvA/oOD1tyoKFWhXnL+g
gvBppoAEjRql1d5PnXJO0nwKnkhtv+bTGKb/5GbPiDRI/ZjUYVxTAnn5HfyJ/KKnofzkcrFNFhET
jqnoN1Yg21kMo+/kx8YmX9o1NyJQ2U2RtLzV5IjT0XD1vkv9As+1O8Du6IZIkoTapFU1W5M6Uchk
xkigWfcbY3smX0ly/AOS+cbQkNb0cdNBgFbfQhhux9uaacl6mWJqCrmc25o7S5nZtADS+3FnyX2G
MMtTdxN+82bxLi32hjUEleH/Y3wYfZDGGszhl0XdOcVAD7BfauQrZM4lzi/z51WpT8U3PPXfBG8U
uSj/F/zMoodtBaYkMlW8PrvSOtymYW1IC4tC8QRrROAKc2XvqRXOm00X/ZbH/xeVX/S3hivj0vMG
eLTcByndfmGGSE5FCmlhRT+p+DhmWYR1JVB8RPvObdND0EK34v22gnB+OH371U8EI52YEslqbZwt
JFHDutJfD1nCQRGJidI/DaEK71IICCJteR+5HZGLC5pqffdyU3RrN06xZsMsv00BM+tC6sHYzkQ7
B9vZtuLRJJJbY44PmxL6NkEE0Zs4exwU6F5RZTgxKo4Et8Okw/CQq72oN+2FAGngwUtvVz0m6icS
445j4/yqq/bnGSO/BSoet0i6SDS4KnJFXTO/m915F7QVfzny6pZ6I3e974YAFrSTIwL+Pxgar1Qx
Gmy9GeJpdJWSgY/unHqbinqhhnqdDCn66/EkF6sngNUxBVgaOIMORdNJimCqC0seF09bh7/l3vp7
LDJX6WrnAtU3E/WvXHpAmWyU0NDTqmAwJKMDYNQdlTVTjoiqUh/0jqxyE6jxn0AEbqbvEYRBCL6O
WnupK4Rppr2sses0zJU8op49fHEkSqkFc3PJsaaVYOBXUfmToFSP+ssugadqVW6cqanDIQAkDmku
3oPI2lr1N1RcGOPOjt2K1bU0i0vdeDaiLJIYjydBseXeX4Zq9kn8mcmiWMVnKGHW+PBv4VeV8U+z
qqJ5wEayBWWBZXou6LvtbAejSdpmFWdyzzNT937NgA40jcPhRaBmbaFOpfreF1ikvVm3L2URytEb
b2JV90OeQM1FB6QNvS9ZGRRNyCDIuUcA88Ri7UcQ62/f1SX8n6CPuHSPf7R7f3ISq3D9A0pPL/zO
R85VRvQ70HVvTj2b7Ms8PpzCsSGMsYUY09B8uuLP48mVwf+ocv2wVsDawndofTpCciUhdoi7crUF
v7vKobBzcdkHyoT1MODxYRpDpN5/8M8pTQE8cQpHFeSS1teAZjyD//Y9PB/00mWwZ6/RqZ6jhhhO
Fhr9xzwAL5cXxXjAORHgLGcz0JCSQAPPeJtNXbPbnr7rpxVJ8/iUacWOdD3TFDObJ1rXs3caQgMj
j9PpRdMlNmgLpEmINzhYENlMea554a+xeq7wAfD//TF6gdrL1bPGlQaV1Li1uTNffr6CWXzkYuJt
KPuVAV8HzxoaMxpQ+15ae84isCX04+uIVnfNnggUylaQAv1GcMPrx2EpOVPkM2evMgXFpDKODG0O
S+zJxPtdlosu9cUIz70vMhZRGOdLLX3jWmtkETnwvgmCue8BjsxBwodRb3uJ/CKOmED8vDmpfCXw
aBeyLegq1a+WwMG3KmhqwCKdWZEcgT7GXyV5OGuWEcmJLbTKFRj6NvWq8uV+dRFGTjYpXRk+IDpt
FOZFOrpXK/CKa+DRZgiL/5udG6osQ3IUUtuXCrYHLHGnJIR8SbhQpaD55HY69FAsV0hqvyWzsz1Q
7oLpvmx0BGmC6qQZvIE3rTrYWFtHrkNcasWreVecIJ29CB7/W6Se+HfxDZOI57bV0SXyQJXFIFYS
ADgkmZ2gXNz1vAIKYAG3rCTijxIiGsL3RryfFg59CvfkQBROJr00O3gdMyyluz3LJXvQFjtg/H0w
BpSXN5pFrPdT9PeRfe9WGyTYBKy+8rb16OARQeKsC7EtmzlfPzV13+dwHOnhUwCson1ZGqyB8pmw
phXTAiC9+SNE50E/GxRxT0RGu2Wp4UJryBaaigG91KDnnXJbNOCNiAM9kdUwxa+gomVGVzdWau+7
VMMb6YXY9OgCjWDL4xOZvuvAgTc3J9MRKndfZzooGEGoBAZFGtpqTaD6hVxaBMRokLkgUQHaAH3i
jOg/ghk1Ih2ekNqPHWTkQKVZiDOfOPbh1cdkTkhNFnsOeREC6WrZaPzXNlns+4yXBEHVuo+xQwEv
us3AP7htZW0eo2U3ieW/d1QFScwTossw7S7lY8hoZvDtlpEdT+IovkQOD05kJ7ydJ7TttqlMsrc4
BwGyyj6X5WoeoxfNm+wYbuOe0XdNhXqrgCyREGVi84qkm3EUs8BZyTc55KqLdrjS1upuGK/n6BcI
X4Jlp/hDNlE4aZRboHWQ86XIRunV/wyMlw3JpY8JLeZUOmHRFxXVawpDQh8m3EF84NfoNbMnOCo0
m5lf/yN1OvFYjFceqB4wvdQVF6P1fnx3E7zLuMyOyQnWA0cCxa0SZ3VaYdngjnpI4FOis3CvPMEU
YgxucwTwrQqDi46nc7NKJVtfwlK3vAh56w8g3jUEVArZEj9yFT15UB4z+IbPyUILjnIdSYDS9ST9
VRUV7ZGONFAUpbDNgnfzZ9bdO4V9ZMu1H8jYr1tKm7XCfUiAhV5Lo2dz323qLQxcrv7ZXqak4wt0
C6k4oNFz/WtfbzBP3pfPrWrBmQ8Gi3eeI9k78q8UGTkSGPrajb1ti91PbAoY6mnIaB1aEYRjGw5u
yxAtEpBMEB55V2Go4ST2paEHViinZqVeyJ0gwNmiCLSwMa6jszvAUXGWuE8oYp1KRrVTr2CVkViC
frtquPO7QjXhEGHWG/JLyUBu0c82LskamqGhLvbXdohn+6G7212UGb3XNp9tE3RGw6CFyEfQ2nG2
AvMEa0nnd94lKiodfV2ldu5JsCW4CCAhdlOWCPdV3bffXrEWHTP1RO176NUcAsjBsjPsLwQEj4MU
NpbjXr3wYmaK3mJTr9g9WZ3h9FTjQbQ63xcgbgfDuTFN7e874D4R5OfSV8siDnFraoMO4Ddom+at
C4FOphMibIYZr4dukGJANv4DMjWjZkizq9IgriDzNRIxzVW+6rtbQcayYj+VxjdclDZ/kOCICakx
hcTQGla/zj1f5LH3BCuKW4IAfNqlwoM0HhgShhdRVzShF5LDaxLY4J1LU6DRdfmqyXB9OIbZV6Me
RdGCTmkrHwG+48QlWrhRkHLuANcySKUNX/dztiDcQs2Pqh5C7ZKqR78CvPYQsKmI3BQK68sodvxs
E0/pff51dTtG6ToYQhM3yZ0jCiWLzynh456lYD54tx/ThqoZCGJZvSbi3bbHL2+y3KXJfuE8tK0S
VWZRBiVOabfEvVFiwGTz5LFA4cRefpbgEMGFwGMY7n9qvj5qRP+5L3dHGovqXGjVW3VmjiZ+Uyrb
injDeZfFgD7pFza3rfievrzVJOUs38q+ODaofhEbS46YQg/dCco7o4TgOxt+VooP2BAFzYE7zLxO
LOVsbmBl8Anp9wwn8mFswIClFzGXlDM7Nsu6lU4WcGSf4MaZdZPPbJKFVM6htPORux4MZtxau7rt
7/ejGKE4uUO2nw7sh4AAjXNmraTZ0qnCop6hB/kUTbJknX1mGo1ZAv1PR/8tABaBnlhGczs24i/U
/HpxjK173CdPeBfKnV6wxfUjhJY5th7QIQIPAPTZm8Y200uuPffZ+LiAZxE0yvAgnNp9AN2JKV1E
/LOIP38Cu+oZ/2Ab12f6te6TgD8rqWlHCR2wyQjGg9cQkPsvjtIYkswSRHjOX5WXFwRrH75FM1Sx
PwXS2V9uAzmL7pO04lkrsKSM/b639CY4VoV9ejqUJ6rAklTataKIoFXuQ1CsiE6PP0SIZeYv+HSD
jzhEDCaoSHqGk2Mf5CMTm0oYzs1iDYTZzBOpeOXaFWsTX5jrbc5cYXTpX1moQABUZ4hz0Ofylhjl
7hV/MIvP1ut/qw+zKVpJAN2DnU5jLw+YLNkjmk3E/V1eYSiXIgud+DNNfAQDpqIPwhgvgsiypzFb
MK9oR9+RkV0o/0Yk1OiKO/FLtzzDKOLyyHLmfOXcQPaUSCSXJwDS41c+i1Gczoh+PqCFi340LzLi
btreIqZbUYmXVfX9A2cLPRsb0v6WNlaYeyj656GiJitTBIWYoCqhmV+hakv64QRpnASrTk3tQi/1
q1KFZ2iKAfmjZos3R/w09CJjxU+GwfgycIJ6wsxkq79Wlw7zOgpDgZmLXzCpCmZQ2ZTvTSE+NjUL
zIXF+2f4lARN28OsyBf9l7yzTECyhoeudENdiwnRab02c3P7G9cIujU44BPK1QfhbUSWTE/YyMPD
z/4f047cDUXjOXWw9cwK3pVjfKb5U964r1Zi8uRChgX/4IZEvGt+DFa+HUWFxmqPFsNBj3gwMbIt
oLE5wEGWJKgSZOA8yGJ7MoAVZkWLimqv2SXcvsmji2s7nZzwc5/+RpDDBPE2tseCF7toh7VzFiY4
5hD3rtSvDZwLp50dTRa43CsjW6770kUE/ftfiZyrEcOza6hbvTZIA9q6/D/W6OSbXqsgDYKzwGuH
xIi1VCoBTSp1K3iWLXc8i/Y24LGI0Wlzm7kavRs1RdDgfe+zTxQk/P9paWcIlC8QCMOtUrE+FxZQ
P2NmxPnConO1uYNE9Zk3UVElk2pSBgOf7q22GKcc+/l1dH3dtyNwFjF7Q9kZ5b1I2qG6mzXCRIRE
fF1mmBsLZmLWvvR14k7uOL+iJaahyCtyRUHjMEP3tvlaEeWX1/T8uWSWhSplaMTQs721fv8tt8pZ
sm8CXmO2CAijpsPsI60Z5pdx68rZ/6/BbM6tlhLt6HcaIOcNgX7KfuTXJU84mW8NGK9VGizoqJKp
c2gmbV77D7BXopeDcviQi2HY/iAS1k/2mpTnHXKqxQROlYpYwAaF2R3asM82rsscTi2nZnXxbsIr
TwaoARuujC28dseMuN33GLGulNsbteRaTTD0jqoX1gfIFBJE5KtSwWnuaa28ZQC2jVyJmDj2YLV3
R92NofEVXxxW6HJv8h+9UTggTUdIyjpFrzi9v+dZTT9xw2JAvd9QpWe6PxoA2wVAmzlP0EkKyFkF
g/wXoloXa4H3Z1/1uEI+dNJnr5Fia45r5jjiH1ZJkqP6k4rTBH6SphaE7AovlCcVIRUWT2RpCd+t
bduFdr6ZEvRmBNs4s7FhhtIeVr/TE/nQvs82y0BTAhWEXtM21UzG8tkcEoyKC/IPyOs7SQSminjs
oP/VX+ks0i9HQpPfl/ltGbG1uiT/dwjh4xoLC73S7ijdsPEbXyJ1jI80rqIcHvzffZ7rkwMLv1zi
/MjzFWZKC4VveY4AMKqsJWuHRpEqRv5HpifovgNGwEthr4vqpHvgchSWPT7xgo/GYJUdDntP5JhH
sWd8h+t0kWx6dJe1HW8Nf58Feyu/VeJZJG7fSe5Qk9rc8SfK7buXmSILR896s9B6lqP93H/clCqc
pEGHI6EIB2lmgavFSdc3rTVGV+6sMpsB82M7kiilwl576Deq1p6CnPwmv4gwsLaw83f/ifqJJvqA
UJRM+SYn4fYMOHPsa0MjU8nttgCT8jN0OteIJoSj7ggmz0Vp2IBCjseHufGSz0lTXaHgAhnEUiTY
ipsJTwVfm1i6u47SkktIEA+vlMBeCAuIMnHH5pt7UpqbXL4IxvDU4gdalIPhWTZ3KowFVU5SDGNk
o4jA7UF+ieXOZ7OU7q+U/r0IeDkPle5JNwRL+vJVYMQh3eo2FkcIZcB/eQP82KeEwo2WC1vaSDNf
QV12E+vOZG3A6a1TaW7s/gg/KhX4twMriKKdtp6kmma90+ncb0gKDHhrxmIfA0bzhjvl3/HLV2aD
CFqRi/kmHTxDtjMxseoi49jYNUP4L2OSVgZPaSLYAEr1rC7TR9XsYpvIzCIH3DQJqcy6RJyNcwAz
tzz5sIRX2uFYLGs8KLnxEanwX6sNkYGQPpNhsytSgETJNkAxWLwjgm+iUll3IJGjNv6piqYYVZaj
mBOGAOZ7cpFcT2zvCX+yhhVFRv87DiapKtWcSgBTMmkx7YS3bsetx5JRxbD9r0jip+1e5MqI2YZs
w6RuQu8NbfVKa2/g81Jt5rIP7L4t16ek7eRu6sbgtGjy73QOYjGUfIPyff+fPhUu36mz9w0jkRuM
Fy7uV6p09PjEigH8dZsxNDwPSUuvmFAaG8uomFXdjAVNISOV0SbxYsFjD093LnBKpEJgUC827W8o
gUpVpCQs72WKIAomP+te5PmQUy+Kf5N/QQnZF5Lty+4Ex7X8qTUEal5py/h3FU+QCi423TBWHhUV
7Pnr/oI13u+JEXBIbXhkLkmOR56zHwcWGOiL0Oxt104JK4ZPMUbn+xl1uyUxErHSzOg0HCh0y706
omlqrKbm02is/twyiCltR9NZA0Qjq09rHbQuIIBVlWmqv2hMiYMCvn3UZwAvGsX7K4vNB+LINVbC
uu2SA0B6aagkTLvmCkTW7lRA4QkbR3T3KLW0IUZIW6Sirc8W8W4Che0MhmsQBHP5zSzUbRoNSS1N
iNJDYK7B7r4bWPy3JQkPbrr/s40tV6MGTRJDLDMfu2yaSmXC5pWxrqDE/MnjVFqhEv72XCGID6ew
5YSlI1/MBqXCwcztnzZQN8CKI/j152j6HLYY1ReLcY044TT/Ji+Svjq6C1JVeiYQe/98gxYDEI1/
pizFz2CS9Yl4oRkQwOCvtWRwzyZnLtwHuhBbscqmBJL7LyDv2RxoQ0F/MTNom8oUrEDAOzpQzD6e
6LVoWJElQxq7sdtMYoYIkc2SlgsNJ0k37w9hp8N5lgBckHF/rZOIdzWvede50Ngd2EdboEbXnLUF
OVh4EvjXrBdr9aV5mo2HeKl223BmQUbbAGrUHY7tK+VreM7XDCaK06ve1g8Uq1B1a002bE5gvwVw
XL5ZkO2ePNNrNE55b/fwvfVd0+px+kDVqe6YKw23UYmMJaO64n4gRxJbU0C5dkqbfTYdUcmlMHtY
mbfIvmsB+ut2O8F/G9Ztdbvjh5K0CoPBdy9vLNNHzO/ZizqR0OTXW8HjIVai8N8pS1xpVBihpOrE
TNm665JvoPvcCnRuTGNxa0UnoUZqtoy+Eqejevvo8BwYhO3gj8OhVyNoqwa6FgH21kzTEBSEJrns
QpBYS3d18bOMWXHl6lk3XV4wk05ya53hRv3UP0gqR5jM1lXAk7Yb+LwXo4tfGSBb+6z/4iYbltwI
AdT5k1Y5WfQ3mI8r2jPA9rIap0/BIGyMwsW7HNUgai38J8/5Jedd82kdLmphjprlVzEP5XbJ58LQ
MPXcP2s6nOGrhXrHUBcHy1pJO1eX89g4FcAq4TmAeBleBHyEA1JxaqaS/3FCQ48PjVv5B0QLkA6B
pCMRigganQEQEWz9Woulr/019UzfzovK8dHwfMsCjvU+uzOiUmxMpZ5VXLtCACO01sDjOv3bzyP+
gc8cGMb93uS0J5GBddReV0tebwdISSmDrQb5ZTCttohoh8JBZ8UNH+ggNy+9p76grzkz498slDXS
8HmHryZa6OHcqkRO1ol+uk4RVsrGwpAXcVz0kkIbkX5xoogDyST3TlL6Ivlj9nA+IrPzDPT3Tqpw
N6SAMS7dq4DvJEsYaECoeIX3NDmd49Y0bcDRtTpMyp4ApqhmrGQ5pga1yofGhP5mtUHvmKy95brU
jUlcF/IUEctPPlMXsX53ZRQ1XvU7zmHIUgJ3/AXjtXyt6h9gVfpYHXnkcTwVhvrRq+iElgRA/4mQ
YFm5yfQ5+soHJSBbdmhsTDG1kj3izIqYTAdpmP/7I9W3U2cv329os1h66ohV9njvvw6vSl+xV6vm
FZVAC4lfDWh5AKgwHmsTp+i41PwGNJRIrGQHmMAIJiHoVIUihsux8pY57kcgN81jVbsLhZ8w0DMQ
BbqMJzeok7DCCy5QtgGmfS/AnO5a99guaslJ3SS4Dk4mqyI3g9Xf7wPK5/wnEBdsBNlp5P8UNxdq
SmX2Nx//8MxoqKX/tKR+4rGCnuO5wGzlT2nBxuGuIe4l6hy77H+z3P3vtDs8z6oNhesPXfu0NjcJ
l/5Wipg20D227yIKBZuvE90RWo4JxdufWlnDTIqTRIIZ4xyBVxBgxHygRNsWgDKvIIRRY6ylximp
YT8vOZd4kbtlcsq8aEis8qt/+8CLajJY1VK7G9SMpUp4aYX1/ePkXovwQKiONF7b9pj1OdM+8+ex
w5wGB4a7/bquzsv/qrtRLPp4jkAtlu609+h23ESeMordN7rFkyvfT8plh1zYwBljn+lNDjG4BSqd
wNS1qet4GE7Smg7rFDYXsui/2EAC27wnGLfrAeL1pVVpjHst56B86G9Wc8Nv/BoRsUmmhf2zx156
jbAtOsB87JlMk2lK8NQ4NVJZVyHxpCdOZ6WvG0Bl4CtVhls4ewrowsNkMKJvqBMTUZCSaTbOl3Fb
mQ34V08pTNyeqLeqGLaZc89JRWBknU3JNfYknUDxwRn3gj5M1hvBQHkyZ+Rk2RtbPA/qPYo5KrtG
g8a3t2uJuNDv7RPJZAnESGdagGgtiF3peBehQX41VB4P11FYbh2OoCyB0t0Iqz9DfHIXezXs641c
uqNF7Ng5WKl3UK+qgynglBAi6eTSB84O655VeDr9pp3bdSL3TUo5ekfdqwwEAimG/AjTbJu8YHdK
giUSuF9OXYSYFW6w9O3oY9lfCAgWqjR/BkLYXrkD9hJDKw4CU/izLWbN4UIGok88UK/ftq4X3Rxo
tyk3aPWHMlHaMkpm6lLE+pU1Mf2b1ddElPnjh9U4vT06z4Z0TPqbu1NjncmHKh1JwXr7/vMgmsSu
2P7vwmB6ydMqkFqM68GiTv17mY5J5KxUJC6+6KUMeng+SVbNpUr6emSgVnaQyl1ljfnS7CIKYGV6
rZ5Mdr3MoZTuvkJHQZZhIdtP0WT7t0B1565pAR7myAtDOWCh4lA6Xcrg2y7a7bqK0XIuc4V9rT74
OXJ+U8EW4nl7QpOvEYOwUaoTaUePsAwp5u0oM2Q8iS5m0E/YCRjBdzhWpwdj+EYOeek/bq6ncqIa
BO1iPAB88HnS7uvyMHSba9UW+/2txIWRRubMyawUiY40RhFe5vs23LOMALxDXa6hr29jnvlGp8fu
2nDDYg/ojBRTw3gJ7ndNDjaOpoc5AmUSl0SMkxihygRkVTcr6BvorqrZAjo0NqNTu+5wLuBj8jx+
o+HpJXALnTUZsyuSP1YaSOue39ZA/ntUwaYmooaYJ4nfnY0UGjPdWVNO+KrHUEyBIZTDCjZ8nanv
OhSocQhFRXbWusIPKI4JU6mJJee1M1gNnpZ/bPz4YtCan89o95o2lMA8clr+pDcxwFzXPNXJ4xY5
8XgOqr5ZOTRKcanoYissvQdgJXs8zPBduBSSRK208dDMAW2qmufyBsg3HBqqZci4XGUCGYc4UhDt
/q5Qj4v4PSM+IuHDnxJLhXcXaRt88G/pbeAEbeqhTuz0bdOKlRpoqehYbjbQ8212XONSAaSIQ8Al
tuydvktukc2fCkBlTr/i+rTKLFieCkWGAYwYJBqPLv0J3ScvjMGAQ1jV3AkqZDWe2AeQ1GCdoRiZ
6ZtJbw7an9RgBz2aHAl/tk2yOUvUpWit6aCrOBETlq1IFy37cRpT+72d9JJa6BivobgJn8RLpqGI
d5T1hNo9r/v4V2/mP9pkUNviwo6wCGD3WnG5UipgLKCbtE1sPi3JJJui5YVA1waldKhmamytbxxM
1LSsIbzdfLb5VkdN6+XMCfWzWI/wSESfA96OFkbW9o8XTQ1sIflM3n3t5EsVNXh2GCQFfLNeXvNz
DEQ5nImR5ma4xnm2tU0RHNLaPTXNaDx8NRfdAJkrIKY/9SrhWzQGek7vXm0BE7/998g1XFHqAJ9O
fYgHNKtcHrg4sqG7DvNqtRtFT/PPstaMHH9FoNdk2HsPS+vJQONEb6+gDmAoXuUo3xWKPRaUnhWx
LGSEn1PS3MlkgvuU9Mtu0IkCx7AKBohmj1MAK2YKqy8P3PJsUKJEgJV/yZld4kL6Say9Sef8ZuZ+
k6IbrWr9y+7jtsWPshIMaqG/J63Le8t1m3KvOAxr9PpggtfFhRPVGU3Gnp6/df+9MKlW+3vWubno
bKSKCBB7U/Gj8H0uXj2cAb8W5CFOKPRvNluZ1/CtUZ+HGKAeY2MVeGR0u/WvRqKfrLBoKHXfzXKQ
tfsbiRCZsY0nWkavXw9gcRIpGufcyw043sAMbHEr4wNRpuV8F47RUXVtbIzePfH6ciDTQXWBOSDy
3u0/1V5eYAA41lg9QuDp6/SHib28rYmcuzz2qum+j0NSNC08cQBwJhNOtr6rIb89uI7IA6Q05bfO
4i8PS6g+gJTDiEdigK5kYzKLcmTLpBxYuWI0PSsycFcSi/YT90Mu4a478kUySzF43lYk/HwpaK10
PAroz5Rab0rh22ghLZBU90TEv8qapyj6NF6Xfvjo64VAx9ogTyuzbupS6j3BUgB93vTUisfpkrEV
73oaB6mXYB4E0k+LKBGzCpZbRp9/NQkW+bD3qd/wsp4/d5snF+NifY15ctj3pLbBQ1prFl7L3kwD
n3lPvnV6rdNf6zIDrAvem7/zv5odrf2ZExNDjhvkO4lDm6Fkr2HBpQdrGkP6H5UHVNd612CTvcp8
yKZOMBq/NY8oaE2Iwv7Ox2wpVIj8TIDueJ+Gf4XBStpLLFr6CDGP2bReQeiTSprdr8mpp2p5xSkf
zFJhY0qXNAOc9GT4ciNctmSWtcqi3kson5w/Sqw5keepaD5cL0FD1cWf+H4+Oickuo0BtbEHpNcB
uehcOfJFQM3eaqiNEjSl6BS0LdSBoUvAuPuLsxedF0+hw26BxxKMNWumrlZBkuoVpmmMsmOSZt9a
5il85Ko9PW5naOHi6zGPktotDMh5zA2GWfxze4E5iRo/rDooAUK6ncoJd2+FjNRPCq6Mqq9Y2b51
/SLoFY4E7LruK17GPYuWnWvLwbxhHqfyQYfe++qIYmrdw2vK5Jf91B8XB0dYBzUtNmhNsjUwiUSq
1IbRnFcHeWRR+eD0csplFUIjaLxCh7A2g2Rpo+id0LorGCc25atx3zUnMGBt4GIGrMLZ4EJFj9H7
VeKJ9KZE73oHycRnBjU4hu78f8ECuR69jdQTK+OW5kNvR/cJvRqpxBcbb5Hz8xjoMy61w9RNxmXm
51PrzWraT38u1Pcgpi46BuaYJxv5Io9X6flKZRo86qRkiHTwI9jUkcihyW2e+mhf2zoupAacKJlU
7snw5lyVByaFm7PaBeCtbN8Ao/XEqTVYbnAOIYcL4BGEd6AAKVL+oPezcn7EvLLyMl1qDqulp9x6
9P0YY5Sa4NOQ/HOxrg5i8XfOxcWQdLyl29iPGmGPJjk6oYq1ru0nsZoFZMh2zWmodzueu98y2ise
W4T9JL83CkkkHLz73D1kIuz78cwnRfkchHmdZtjaQegSos3EOwK5rbF4OzYXGiuIIG1u3ya3M5bf
ZhR/gTpLxjNgs9hyhdCqRnUMQqQjWJd+BMM8g1UpU/sc3TwzpF6vDWiuZU9NkB3EE7jZv5ImatxW
zhPDasI85VIE0Z2LB7pWDoXktv2AbkE62OW/ptersSk9fLxQ+ioe0vVklttXbalbqDWt1sy3IbAK
3siz59q2G8MEaxZVzMzqVmwPe2v9Jf94E8Z5xc4pWhrK8B+vwUtLzBjurbxNADXTwBIxWZQesrpb
Upe2ZmVvMEJk7emTMso6BpSYzSg/fx7BXHLUw6hxDwh6BWR6LGgpErLvMujaQtxaXGuhQheSsbuD
nmUIHSrer9P9T0KFTvXz7H0kbPZhsh+d7xXs2MBO1Z8Jr622/mFhGowKiEjP2130T7eKCyoLOuGq
iqscxgdrLER43xQxErEuLAEnZdJkSbPj5K8rJygKm2cnHzjRHT/LNuH8SQzUApd4EVYmgQBlVas9
HU092UCbH52KpFkVKtYGXGtIobTFz4v+bgT12pAuuEQgImq5BVvS13v4JBKhWGL+Zwo6310dARqD
gqKD36D9cYFdmZd6Y3/xgH9zxLcUovjEZikTBljKMsE0XROWfDb6mkhcfIT4m+ixtHHgwwuTWXmt
L5n8iOcWHTT0JGbuohP6TmcbU8ZL4FaXBBEfP0JtyMJhjV3UglPqDzeYfOsbT5390TcZddDaR01U
fqO4ps+PideIQ3D9EP3uQPW6pXcTWx7wZwK0oPqLzT3Bp8TMfHuOcZRAJEvoeOh+j6BFP+f8f3yu
ltTKdUh15dBtMHKnr7YMR/NwU/dED1HmwFe/f5FCr4weSnwnVwDeZLmBl/7LQzrwg5KVT8PNrpV6
lnhqfdJq9gUzlbFuKJldBQa5oHmtsAh4vyojyVl0gn8WfI36HL7r2VAkkWG/rk9Pko4NnSsjej8g
C7ajQJ3sV4H1fsnjLWydHHD64gR+KN00lx/yxUQ+oCQKtrcgUoPF11BgbAR56vtsa9jtXBSHPQJY
oTJMexhFA6AqcWkEb3XW1wSBnsQy2uYSev7R75WVgi4Cy89nAMAX7X4BSlrD3Z+DG6IG4DEGOc88
M8LJvrikfweWJ72Uaee088Zwn2mXah7FU7t76akFBWUYdA1OWCR7TniXQeLdzVm8aCSRP1LLJ0Dj
KpdDIMoeyeIpVTvz2KoicUJuUJm7IccIaauEId8RT0ofnIrTdsMQ1V1HTLiAA9hxBukpvXcE2gzO
Nxz2gbFPX/Y+D5cGF6CMCAjvBZtUTFoeMRy/Ubgi/rfZJf1nSxu5Dmotv1/pZpjDXwwQeJ9ynAkl
jxeduiZn3cCEWe4rfn9CIRV4+9UVt3Okq1g+PtuaVNqIdMqo1mma1r5Bza/2dQqhWoGDqZWANXLs
JkdsJOyKT0WWkwZG/mztKgdbR/cMzPutzOjzH62vv1z3jWDpfEfFQWCmDWe4eA/Yj+UBT7+sQ1iI
rXlAa/J9N2NuR7Wckx/yYkiMbV+GNs6+4/OUVgDb0Xr3h9AGD10rtesfXNsia9PafB6AfDCtyEGP
RwBUPiJmGgZskqkJTlX8d30tR1VQ3s1MDHzpChSmvPbs3wgiz/XuX9W75Ex5lYL5FioltYO3grJq
FqdhtJv4cxq7JTkXGkVFXbRJesZQEER99uSSxOHJ6WwKoFCwVPPIx7oVdPnf6YT4Z9CGRLCdq9jm
J7Etf+++hyvVoKQP/g9yvLNhvP7XBdsh8Whk9iBR/xj9A811Mbu9JiaRJZKWT5wuJ2MeA6QkgHrP
pf/90zFWpl3Qo3xKWT1BD2a6aLUjVWf8bpnHsMJKDWTczU7RNFTC6A1kwkPha92KdeouAgpVrN8D
7Qxv/pxt9Ti4MivUiiKbG/yjt7uZKyFjs/J06P6mL9yQkRwVS45t6ypH+Ec9UkGc/XqUODcd1ezz
uwn4n//4hZ5Xq1bsHpvVzLmJWBU5Bh/ZEGE8HG7VxNXCDtL96zlh7PJfSBL055YfJ0RCXed1DTx8
H+WxbBFYLbEVia7FMUSC4RrKA6VG9fMACxBFguR9+bm5qAZSAkMkJNgpY5UAQwthlQECL2wcmbQl
fIu+Xts+ir8S3ceFwgUwbHSjKWEaPnkTgsS1rMz4k8Y04RU18pgH3aGnicTdSAgYuOM0DOhVrV8S
WHs5Ju/yQF30eY5+DWvykSliABYwbSR6y0zgMeD0O5AYCWOrdWOtFC+qxhDvn/m1XMcBsnJHz5Fo
H3pNhDqBVp7c8bxznJiUJr+kLn3ZrBNqhkcZRgjMpwjZRT7mmHTRqfnNLxd/fx+47DkyEErRhKSj
ZNqk/TfMTmBHCqriiZYMKcFXHFOSwTad5MjD6hCO2qoBuyJc5luqCbtywevarAGGK6pVcHZa9MBU
vrSJ3L7jPtiRN2sTLFTLjUUEPzG495QRKpOv37H3xSXIUU7S0dNA2E7oDU9vqOmYpgGLDHVIc5IW
vM3QmYRNLNC34NzeEEi/DX/3gmC6wpgPtogNjkXMAwufCoPJ4tHLDpOc2lDrWIp4aoC4UTNj48Iz
0mNBjwCw348SnZ39S2bF9xkX0XXnZSvobxT+llygDhgoLIbugBSB7oGp2aOKDQthIdnieFsSAKlo
b4M4gqAM9rkBX6VmWN1rlDaIuRhPEwn4osvKu43GWhM6jThUuEuflx1kRMpjoeByFGvX/8piPD3O
D9EluRdDehIoW9ss15Ie9M74AYtQ8BquQFjnVIIriEoh4+GC3Q1Xnktl8VOn/PirfOCw0n71R3VO
923oeUGbz4KxHWqgMjUfmWJJ0wltwiAh8U3vrYPMIwmkhu1vJVO4wDtU4xFauUot4EBa1qcdEsvD
b04j+qu/q++Q0V1DZHhvIRp5EG+BpHA+bVZr422YyMYlKVPXHDBcPItmK+kFB6GeXHE2zAL3NXJI
hdv1wRKtGPYD4hAcO6VDNwR/3oNBjVGzNNkwjAXz8MaxugKsQeE9E9RYD4YHETCfbUEkVxMf3ZuG
XOujl6VVmJNNQIV8ISjEzkkQaTanxCbqjGtaguU8ri1EttcqYKc1wOdGFR934XyHoz6/6xwbcE7T
Oup0BRBsjF9CBaM4Yn8jZPYXEvfnusK90JjIUF1e2EfraMsNBSp2pmkssHauiSHCGvb5fRurQjAV
XlffZBXI1IN5lwHstUZ28+WL/gvfHHUMC4gEGwQiCORtoh3smLf1zUrSXLhZSFrt1aXRzk4zpn5T
Dh0TEmcLvhxmWTTaDpVfk64/6XtdiYbzIY/BmNyGV7g42X5+HvICI8RC+z9tDRX0NMXo9QmMRZ8L
+MSklhSPgFN3a1sT4mC2P5Lnqr5FRQ3i8bVmv+PD6l9Idd4mO0uc1rFo8UMHja/te8gjZ2KORmfI
8YPWWMRoj/nv3PxNPvJU9WQRve83GqKcvujRVg6QVmHJqcl/V8lxNjKNwpdRz03gt7FKh4SbIf4Y
cCBCS4hjqYKJ+XGAgl6YW/vf6Sg5SrBsh8kQOVs4qkgS0ud87Mn9VtUdPLFncHz36suwYF+6dNWV
/IQIUS3sTcd1aLiNZNAPzfQccYpQS2Q5MQVhb67zWEBV7I3Ea5H9XNstTGgw9Vm/ppvVFKTlYCpl
AFo18ie0WZq1aKRsWdtsbZ3F1h7N8ljDeld+auB3wg4eSUeueFy/x+UabRlF0sHeDbDJu7qQdXJq
/wkhccoYBQiXHvYlS8xTGm5bfs2Lcq+1BuNt3uq7HhRTUPqMraWxpTRIYUnGITs986LlSNXp8qHq
U92OglN5h7rrbKPpSoK4z84KOcjrrNFlOvtk+mxUugsi19CNwuUzQVXq0WNj3BRQ2BsbNZ8b4TVo
Ja6uglBpNsf6EbV3OaA52GFpuxvNzaHQByqYbUjhuRKlDsq0Gv9XNhJ5sDJxhJnla7C19xI2pwvp
UrNzpz3xZc2gbb/l7UO6NQs6xFSt47s0G3b6ZCW1XEPj9ixaeM2Fp6lLAUXPmgSb5F7J8gn4WhQX
x/d4YFJ+Ve8AsO8b3B4SZi3gMSq5532rN2hF+DFuXVBSOIkVwyJ/WgEURuJoC0WrHxUiARRxy6Ca
GgFx+UzBMUZWWtpIc/qOTccaGw2u/DBOXtsJ7xNTnAbzUh3QFTb3g+KusU0tEN/pAD8lnoUUhU3M
yWBdAtIh0K/FYCLcogsIDfXOVxJ+Jx97IbzNDo205TTzXF2O/XuOOFtqZjpJfnO2woug1t2GqcT9
FxrWPyqREiDor5h2+qF7uha+ZfX9YI/7luLcXfi1oJFLjrhBKMoFl6WeK0lb5CmkOBUL5W4bTry0
lZdfKZzPAXGIel4rYR5q0BTujUa39Q5y4+SRoVGcdc7Z72qlpn+ovr2zZrzEJIz/KGrwgtHkhPeN
jY5B52dbtWyFyjofVhfMVKW4jYuG8LSOG3/aBqCazv2THi3rtdGwl9WQc1mymkb5R357/M0dVsPU
05t86qSRpmOB6SO9EDLBsyFg82bglqSsiQm1oiRWtCeBr+QkBYBpc1/4i5u63JbdZkNtdkY3KHW8
or9RArlZlrD6ANPPHJ53p9c63FdclYQpQxbZLC0NB2emtO0iZx6rbDcxTcIqEHkKOH01udf0W5UV
VLp3rlZ0NWeXCrx3hVNlYKbw8L9VkCuduZhQhAC8wSrvut2sEw3TmWuOvK1uomH6R8nbdSmwnrlx
LjqPi+zr9xHPlvJ7P2TO69lrTK1ScBNz8who5dQ6B36FaZznV6OW5Y2xeAxayA3nQR3Vn99ZJAMB
ShnpbK9OfbBCSYQZImeNLwiD/JRx0shHdwCPyeIwv2ArSg4A/YS9ho1JcexJ1/NHyiFMumQHvcPJ
lzaBnnQfUVlJAh5GGAz/vrn9UfkEFl2GHp/fMoGr734PLxz4ucO6PRjjTEmahkTCao5C0HGEA2xH
AVdyRCa6OaUGOoL+1pWljZP4AKSOzNm23Pbw1tQgG5UY1jVEWNib2cKvv5Wy8YJR4mgCGMV+kIDP
pEERmZtPgHUWtOFu7TO2peX1BUnM0fqKLYEYHn31i7myw2ZrJnxjokyt1FYsu17cyvpj2iOvg1tV
3kDbR3rfh3wByhrT1kxwWEpCZ6+VtgktkA3izyuqBMFDfzskgaJAyossYBSYaiGLLzg/tfwXaqVz
8o4Ss+BV8z0ZsrRx+UxD2HaNjfRG51gQwoXyNbcv74OSikY02uEgko8QF4qPrFy/Kdc5z+EIvGXI
XG+Lhb1xyinDBmMSq/MT4uHnRa6wsaCVhx9TTuELXR/uyrf3woP9AixlueiTpUvf8fLxRAtpjcHs
MR0Zf/e30PzJA1Wq4FzAhaAtP+VYriq5u/pFbcLixJjY2BQHZ24Y6+0OPw3NRj9rBxoQYvcT/SXm
+EwtxV7XbsJK08oh2p0rNJcSOcauOuOs8Dl6nH5qPBo4T3+LMZf6LdkFw2OjZwPdoNQ+Uh1KywEL
g2ajF3N2X4HYnx+NAc7R3r45etTB/10kjBzFeF/fkRo2nDTTKYtTmmlhG4zk3mkrHpk5bEuh1ZAf
i294RUmBrOBriywnEO2ubTg+4TPWeUkrrLj2/ybCMDPZLX7GdBg20OTusUZ/okX+Pj0G51eREJTH
U65lJ2pJTlmpECsGNG+v9kpDXMtFMOgIm5VZhKv9YQBmBow67fqqDZgAoQTMSPPk2Sfn4Wd0chBS
FqBW/O3LEPxqEBXb5tCihQxFF8nqDdwi+UOU9QsuEXo6LwiGmdwb8F60IcShf7Xvhoj6eMCJbH1L
ZTXhi9AIJ5ZtLwAF2s48O+kSAwG8zvqXj13+BQGBfD0V9RIEQRhuWYskUjyyDvC9nknkuGQwD2HW
CE0BNK2OwlDThKzZdCluk4G9oqERAXQJDZizcMIkOJyYHRsQ5b3VFzlWLF38Ym1I2PMISJSxXOxz
pvsickfzuQEXJ9EaIj1ocLE6/MW4UmLzzA6u7FnZ4hz4ICu+zkWTG823a9OG+MEbOsbsTe2MyuhH
Y61p0yiNRo7TfIHUw+Ya7/Lr6/V4bGr1C5v8jyrp6KwRYQMDrL9413c781apce+snallbfBxPPfd
hpfU8Z6rqhvhczahqpw3BKtqaflg425nyPrKicomJ+QEinxusP8pdkt4eOC72LJwB0Wj+1YkMssN
71RK1AA1b73yYGb+aqYg2hY6PYuj3KNJQi+cM+zyHWwUs1liWy5PEO1/DHUKBbUuLVtuGXsx79s/
GOj8DHQSM6q4dkhjLQowPFVX9utmCSkz8iDK6lj1JVGphWl7yYCABONv+RNgZww3ewOmpeUuIrUH
w2ZiULn2TJ1P00xZaL2Ldz88nZlSRo7DPnZy7cQDMW2GsiNkK0oQPWX7yiuq2lh1Gn2hEMzR2Jnz
L7kMkQPB3aUasnupBk23Edd1ujNeXGxcwqi8Orxw1O9OAAuI4eUEpW9gCYgPTYDYawYvrnHQwpWX
4oBOfGmx/+eItPWgbywExkVPsHNeA6JEZ4F0HuACiUW7p8eZdAMl0RlUiXuJgCYGUY2eQdDTt1za
1Y+JqgQksycUFRctxXuR1o83cTjIYvc672ODcl3id1QAPer9h6PGBvtOuJMnDLxR7j0covIE5TsZ
hzLjnCQzjqwyrR/ZD088+7/JqIsAuOj2HEsiFWeTfxyDySuv2LGNR/55UNBM7HNZEXOlV9vVUz5a
3rehRttq62yIBBxadgA2/CTG90APYBElbceXPG4ubWESgo+x0Hfl1GSc6weO05MnbEoHCZvyOdG8
BN3h4OTOyxqzPE8MtMk3CJFbJ9sBbhvjIRtsg0YnCNFc9kPOboF8AyRr1u+2KV7hcx6vhIgZkpjl
BljpfiazOcSugZmKcHFQTuokqGiV9At9ljDTkgRDPE/TfnqTz57aRibCFyQbVR5ZYMVEWUOdV8MS
hOLjtMhwcyD3tTamGZWf/zm84xSoORzBcj/TKWDK9K8EaDP2OKOrd6zt1PZpTqj+3vK44GwmWkNc
BC+hgZuLTyIAqN1uq2PsKzWAoMPzEhQ4nFCiO0fpTgbIpQkXR08daOacpucqxRO1ZyTooS3mVW5G
EHNiFcDnTfiE+FdWZR5Z6aGJkhM9YyraFBoK+WxgC9h75Tp3g3YDWkiB9rQ0V24Buw94v5ZFKBJ6
xuQHHJ7owxpiUFye/84zALOVl+OUQib91mOCSfxoMR2OK73Kpc67t9y67sbS/UwVyGr89N0iIXTj
aMZc3oN7jBGuR0TAikGisN6gfYuriQFX8L7W6WmXWZ8Wte5qNifPbe83BPCxEi9Qq2sSPOljwLOf
9Tk1S0lLyo8TBYfz6hl22nVREG8CFd3xdzWxrGacXg0VkW0pbL+fAOaskjOn/vkGkRCLCCZ1UKxU
wX6zgaqqGnz+f1T23tzkOzLFrh6ndVudf1YU7xGv8JxlOdjuzaf1Y8yBoklSf2Jmkwxrgufo/yYu
7iCh9TC70qWy+JG/qSNW26+vFXgeHKrXeIgKCV/t8cDqTov9DnqcOkviWg8eehA3tS4eIm+En8f6
k0K6BXZBhZexiBiOo5isPLG2Fs+1GsRVWWf4KqWu8P6mrzdYktyHXVnlZv7+0px/4eomn730hO2n
Y6v5Lo+nXVz1ttgpC33QmW/J/DJ2pHSNmSObeJrhzcu1s1K3KhlbdfbUcfDYHyYdixx/9tktY8Yp
d1AljFJH3+SPCUTmwGPP6LH1LQY9r1K6OTdv5J+zLHoSImt615RBbznfAxd8E91x40wXD4BnH+Fk
Impr2Vq83/Pa6RL8wPr/bqmuVWro7RB2bFMrijDcu2PhY+6MkVHaunRp8Tjlh0b3WH8wuDBP5Vyb
/wLaxnoCZgwBjR1LPKJuEjCqPYTJjYGx34zEs8IsYYaWk31TfUITYXJQCG/8hdpzIOUpABpI/845
P6AKsSoSHBJvscoooCQvA40oak8QmA3eg9ixHE9YKsefDnXAIotU0p0yskcSiZ6s6beDgTTy/M6L
Wq70q5oMChFOpgxzNw5+WeBlTz3gVKwgifSqK+HWDm66RCwGkQZS4bSGhcpEqYpWGxwP++u2hqxE
QU08wSaBi3hOtWfoRWio3bbQFwV6mO13QcyAYwJGUYU+gM3rb9tQeioDtt4SWS8sqR3+hBOr619G
yJUjuifqO7XfyfAmxuAH93U+2P+oqEUW2vXdx64DPS70wypQuEgvH3YDWaq6UcKzxJNm0lKhnEVp
ygJcTre3SW9lyKoMvVgqVqPFhabSi7WF24fUq93Rh6o0U2Qtj66vOFGWQdVZm4fvXV/J499seLsm
R+1RNHxJUC4uYmH2Xvq5Kv3oLRXp7BotJMkNJ/mQbhHtQjp6Njjp5hdJ3s8S5zuzKTDSyv0zf6mQ
HE+V1uLnr+naUDjthgQSSyYf+de5KHJVvSFlGyoWY+ZKPIyu01dw9/1VAcM1bhfTibAkM9BlEEMa
VYDH3kkqtbpcPYwFme4KQzSZp/dtQv5xpUODEFf68nXz3mH6vnlJxN/KKzQBSuexSprhCES2qspd
o0NUjppsj6tsk3IslHfFt1HcGztfvHfUhRN/Tdl/+/Zx9O7sKWZyXecZ/NaIwEn9yn7/RqbgmYmh
AYWFqLk2wvvNQFCJCVo/cy3QZcGcygSGIoBw6R6Ry1OFwVmMWOqxJVh1OiidRrgSDfOvdfeTmJEH
iqcwUwfPwjn2j/MybvoyoBpenHP/nDltBcaOc2VofsoZp7gHppFdzR5U6rMBwOozhDZUneCHg7vG
aUFTKWNvcrORHmfpG6YkdoZkTwyBOLsKmvR+ou/tHA7MAyNFt6qGuCfP95Uok4K5D9Q/B37HqWo6
WEkHnLP0Ak5wNa34eL/runltmatyOSTggkoWSXyMUq6yHsHghRhFSoH94ogYQbz3tvd3UCERyJ18
d60D3vWY4+XOyBhpEABoFSAwochtfUxhgg2vG/hSRQBDAt6AyEnqP9Nc9rFuKqIxkgtMy5VHT9tK
v8nsvqsbcPbDv2iqlkXt9QtcohE25E6QT2c4kei71kRhFXMyrVBIpqBilPBPWkJloDw1UR9v84e7
JGwwKiJGY2cxxmYhnRwAww2RigubmuBhWCUQW9MlFnMRftg+Qvy+GaqD6xooUQ68PcVN6Ps2L38f
A/VXIpjLzyQEuxZStwLvkUf49V1I4ShksPLe3fdmwyJjvL32pc9384yUvRt9sIktJnh0gFFLhVck
FPGy8JM8ULyw0zvPEhYRy+zzOzhzdqnEsIQKje7KT4G1WMTa64P6j9Ur8sfSY7Jwq0wD8ox6guVo
YMR4Lh49K1dCjpBtx4AvCHwZUAZ504kDiIeEv+vT9Ha8bTxjN+F5opgcNPpbxBI5gNEeQvsqppMx
a5ghNdnA6a7er+GFvHdK+vREZRjbonl7haLIU+Wfz9NdiYpAytt8Ta9vqqsBb3jKQ3qO0XwaZWW6
VfyTcxtuDGJANiJ0UAYD07o8m2oUc3s7LLhBX6yZ8guVXX4xz7l9A7kcCLSEBM4TbIvrVu6WupWa
zVbDlGkyTE5VsIi1/mkq+l7LNXswicCy+iv3cPMiz23BGTtoabWruFLE/IYdtPUgUUxL4WRIN27K
uMSlVCaQfChyio3M8mjp7vNzi6Y8G0oNHK8FsstncMbifrXWCxc1CKBV8cFlaHdOXFenEc4Aup9C
7H6Ljn/dfd923qnPbRSaUxpPX5wKM5lYXUwLHo+vQVoBdzYSK7eQT+qgqTHqIOYByzHRTqBtppoc
isUiw7oeNfI5cHs+6gSNmXckKcXUJXRErskWoMkWL/Ue44dOCEV+u04KM4m8Mo37f+OaXCMg6X0T
/jF+rNAzqWfFylvgLxqFBv8mPuteUm5KUya0R2t0ppByRSys+xPqy3seW6cBvDsXN7Q8yJu9rNAr
KeMDZykKnvLw6FwWtn2hSmYp2g1Fpk2QsPClPHItoBW52ilDAn28ld7BvE2c/Xq78JDz4OW1T6u+
7zBOT+rTs1QP/V1rAt8OSBEXefVdVhpfBcGKSfOxMawE8ReonpwYD58JQOCHRG3H8Fznhj1ORP0V
D4af56rAfgBhemZik2KSXyOK8naSFQXUjqd0ItoEQbka4Z478oAULXLfvfiCrM5DFTrk8wwhT9WO
kisJY9YqhqNdVg5RsUGiU42/6sR1fID9DwtEo4qRZWq7u04BLgnsoZ46wHVlZdxcsq3bpr1kxdDR
+IDq76TglS3wDFDNgm2lQ7yvvwXpGupOJSRbXH8IA0W6OW+0NA6cIm10+a+xAETB0pYvAHyhJ3E0
dZialNtkNlS4iLYwnLHAqXorbJ44QXyyLZICMfeY1+dZTRvS1BcWOMmOTlO9OjIFrjcUbO4qaZJ3
9VWGgloW3Ymlpu9/QYkZDi7RmE0sBtFV8SchDz8C79kdqa/Et37unnSOpN3nyfrROW9QqrUow+9m
7vdQYDI4xUDjy6M8z3Dy7Y7YRzzkw+oBL41pw2q228VjeyauwfppnHXELw+0690Ji+ojsqvjQ4PE
OwyNXc4thV7QDwHv7s5WtjQUgH0G2+YzT2tt+miMLxr1YgQHh1t9dRt/82KNi2iBC7Nz+b0CSBjs
39O/DI3TolyCR96OW4KP2LC/iMCjdY32IBx5NwNC8GOUkYNuWQN0GipW7WX3M5EZgPXQUGqtfzvR
rWdMmmimxrQecV3RotQXfcOdiLAH5H6QtHWKW3xhHIo8Ly/dLEmoEA4QJWzIur1y2hzutsKrbTlz
cExLykhik31tM7Iqybholo7sPqW5bgO//TJHmE5MeTpcJLsq0Ys5zwZx9m8TBRcCEJQa/joP3Ann
ZcH725aF1dp9uQjbtaKO4VWy4YFz61ae4WTrJ7BcS42rS8Oh+QLnb1OiwbY6GcrKeCmKlxRVGZkB
gKxee6h8ky6r+L0qakwZwDhgIr/kmWJpcYL5Z9mC0mlT+O3BdFTdW6MDjbX3na9eyzC6S3XrzPZb
NSDnjkdp+MbCo8c2iB2ow/YEUTm6PLQlSljzNmAZ6FOusD+zCCOdEmhHwFix/tHC+TytLkLGK/nc
F266Wx2nORNw6SHpzexg8rY4JjwTgDm0GfckJCiGFG+Gj+ZIdx8+Tahg+hU9dg2fHX8rt2Et7cAC
OffuvracRJaQafLRs71EL1YLBfiJOBLxW7yAToGkJ/iIgWe86P4v6M+mFX5HW1tiaqkI2sfenBZn
T1LUdqhbzhHv/chE2wp01d00CnBJM/jnnc82m385rjMpOogYrpfWwJbTSc3DXYjtqfSq+t9vbfek
E7wULM9JT9Di8OLHneQdtDZrnwedD9hZJLx3qf3hA9nj8Ba7C0+vbM+TzE1rarirFU4neVojU67f
UhET5CEVMmmS4B23ToN+EEKyAOUgtYGqOldU3HFvT8g/DXT5d9aCizzEyIpOO5PXAdbAMQt+HpLt
DpNwM+kXAW7ng1oYf1nn4D99vVsJrlsRanryZPO+DQ3sGIWTwMoP2mip47Vv07QKn8RcdwyFizkz
X6HR8mMdgP8OhFgcIIwoerVMPOwAW2oBIZtJsxKVyfKwzpVVERzSP0EwmaTvUQIbtLbwD+mIsGKB
t5f3wRfIlbDjQ2RiNkXejMae4vyCJ+Ng7VbYTe75zhZ4Czasc40LmTSeyuBdzD67uk55qa8v3wdS
62IFOVY1h9y4nO3SmaGNkje/b3dCBLHs2c/+wOkrMAvUYuHstyVae70p9z1/LT4FzV3CVrGTWxew
wUuKmbtFxOhYzBls/tyIaC3tNb6l1gWu40Kmo5A6tEfS9rh3XGPR26CXcEL6x/mOzFWYzv2G2dNw
FQ9UgA11nVFpkB61P1l6GxQ3e7rxYrBH6l8BZnDASdCcT2OF4UXknykihU5B8Ct9S77jK5atTvRW
g5nWWjauOaHm2IreWxpHpR6m+jdx4n0V6b+NYFgsfOWlKmw7qrDqY6UxT0alknhUz0ND7wA9yJ8E
QGHjn/0OTk6fqkRpaHJbZxjP6glJMjhngEPsFGu14QeTd3dZcsUN2qTpoyFOHeoE3RPFpaVA3IP3
/nqNk75XaYQ80r+EkHEqTj30xrvXKdCIU+YNpSjsCQwwZdyZcFGZ5yUamsx9GY1c0sE/2BR/1eaB
9MHwE6xeUy1vmpc9bgEfYLZyzpGoD13bR8u87kNSDQ/QVOmPkUPLzLZz3sg+9JByPwd4Oqj+YJfF
bu/4tc6OGb6L69oul/Cy+OQS4BgLGUjGgLHWqVbNXDosGO1gVUMjnMV64ah3EConeEl5oqhq4wX9
YdvMwiOL+mNlCaVN/pGI6L88nRqZO7JEdk/M1E73u/B6LwneAOWCPeuJHavZxIKnRUeWUmOYJ1cU
0YRlaNafkpxldPJFXUJaqzwpun3HJzwl4nmJp3M3WHDW6qxU93wmJq7W0SMGM2ZcP0vHdn06JoBL
4qQCqC93gcQDviGKThG2TJsNVc3ritEIKQFMvG+Jx3VsUJR0zBqdczmOF2HMcgyX5Pz7x97bImC8
GpXbdAzfFpY+dNCWt7oxseBRj+MLqDX3F2ZftPBx2XMtEO3eI1YrpRWXEED0sUFg/4F395ACtl1g
BxVxnNZaK/3qUE9yaoa9yAH6LmXjfgM/nA4cw/azlObZwclf6TKru6ED9aJad9m2WM5LzWUQtyO8
FP7klhcdi0HglcYxv+uJD/9sM76JGUVuSXeGKnbhTyWhltNW5Rgb+BwDyllTaXTNwbk9U75gQ1UU
2SOu+WuKLZkyu/rDj2oIwzbfWydu/X4OMD2eJ3JvaB+D+IiWEf7cBqiTQuvxGuTZRldtnggwp4VY
yDxUx40ya4ChRGe2K9LbYToN0+XuaeEiOnH6JWDp38QZIv+RM/NTp1SXMFSyHMJN+sSO/HnTBK6i
7HNDRdGOVdRKI1schZHvU2UNy3aNSEEAUB7d+h+o2pJVc+zNI2jkEhp0TfkDYULDzeCedvS62POh
MRTP+cjVMmYO01knWmq/yVthgQzTrDYicwX5wTB4Wn2/7ff8gTCjjshcR+BhQeD3A9S56V+sF28K
WSCsGKIT88Exqag+Zd67sPZ02tofPTXOnr/YAXnBckaX0bjoq5eqbTX54ZbWSyZ07+9GlcYdKj+3
oY/PKz+DrAm/xlcUV9h6XlFkPhQb63ktlif4K5212QtVFftssHT7B8zhsJDtrmKbuSXq3nxcusl8
xUU6Mg4L3mDdP9seIrID/BjQs3lhzzlXBG/2L+nTtAohmWKIsKG0lL3IlI6BiVkVv8G9fbcI/dRR
FPyFGAIQ/RNLjtmsJp9flVLfvywrcljABKKSIDJzfcuGSi2b/BclBh54ACZu6kSqIIQ13qBhghtC
zodJQaeGaZAhA9xr587gwtRd0EFNetHRoUxg5pekActWuSYNJRBMWZ/KK2qqGInxIVDVXGIjj84v
OJyt+pxeEZVO95WfDSarUC4Xneq0mjxU7eHytA1q/F4kIO8ZH/Pw7OjyqmIBm0c+JpRGE/oIR/5H
byHab4Wt3mzmk2thIYA2hLSclQF8k0Md3vVlhn3AK5S5RN0OnQVcLLXP+EscPmMZ0Aorvo4NMv3X
GACpwD7YmocH2KeWtYoRf7pQBOQZHeYFc5n/GOjNUZTrFGl0FheFYd2wCFs2y4tcJMMSEGKSlqTu
cM87rOxzKWnlkesMY4mket12HojyzPOc5Jdv8CFwdWbItxTDIfuBx2CLQ94Gldd/OcRrW6vCKRLq
bzAksxrskV0P+sIyt65PTxCb3NLll2C+EhDIlzk2/7iOdydNkEtai+e0Y+pWjvvgMe6Geqj2Ld6o
k3lCFHRjENwd03WPfn8Ou/cnPCSa02acbVDZxU6th1OxlNVtNzezIgmWEQg4dF90TzebasdzJu9Q
5v6zc6u8P5G/gtdeMtuSTG5+uMnow/HpYRE+6NpWQMaSjeOgRU8ExlNAeeBOPRM3Dbp6h5fCyq+l
SpwdPTfEsHg4e4Y6UKN5ikD7nwHLVOrhBooDts+VyB4knvxNDHDOg8+CqoAzFo5VWuirOhWmNGuw
sODwBuSyzTRu9KnSwxJ6Xe3lwV9XBAdBGK5Oo/OYh/VvjTSzxk4yyVnAcx5t8WD4+BRVc73tJOAk
/czT/Ms86zqEEaXOGXsMHbkIlSMyVlBXcppKAKJqozeSGHGffok3F5OxGD5NcFmVP+WN1MPM3KlI
dH2sfdPrb5Y/k0e8DwP8zMYrIWx0COQf5xRpRR52jQWfTgyd0bJHpudMOUkWya+KTqYGf0ZdiW9D
GMssd5Pu/cYF2fCKQe19jFLXgnQhX24KaBcAQfnJAhtJuxIrK4D0C5lajlA0OcU8V0jfJwo8HoaZ
x8EEWZ3s/lUDiQjPsEHCrCETqiqkQi28uauk2HLOcZwVqZfpa9wApn+UIFaS48OqflyJ/ailyW6r
kw0jn3lv188MnZ5E7UYWFIEnobmFLX6MwH8GsJA5KsJ7SCkoEHlpaivmo544FOvJps65GiaOLGqI
p9U1ht3Y87Q2MJVLBbL2haHRJAbBhnPPXslL20+Ii9jyKj3ApIaak8qLx1zG1uIWtf5zN0JR77yE
2ZhkT7N/B27evF2sRwO91FVOSX/asXIK/pfPGS5uEf22DjbgNBypFjLlkDUHidcqwlIj0tYgwza9
uJj0rYtz2CYrLI+H6KfgoWTcLZjZ3iSLs52IGrxUOJDPOsKFJ7yz7d7zi8Dh/5WttRrEIXKVnjTi
92twHzUpa19T9qWUT44BcFFhPZaHSK3ju+r2DKZCzuIs0ovKNKBN28Tg3VpLylz9jV1rc9KUVy2L
IP7TzO8Dtc1LLpsWjIamjIEeAnmZPFo8t2co1jB3xYucEhYHmpGorDgYQRq9YhxmM74oRAwNBiyJ
rf0y0wHnzv63NW8UnvO5QNYfHEXRNl9XwzMBnTCWE76jHbZkpsiI6P+2LTMuGnflvVjdBuA9xKXd
lv8knebiaIKuiFuN9I5AzwebL/iOMHLGPJ3nr02s+8D29x6BlNFgcW4e/pXLH8Ufad+LAzYUiZ6I
ranaXAXZwPNfjEPJeUinEUoOLHIZ0ygZwHanK8eEO6h3CMyGkKIZPy0FyjrTfGOhkDb354wFDwuW
J9Pb6noD1MnIMQrHIWMz4upvKmVEQLvSLzzGW3VM/qCMZr2CE/0tgFgh5aoRTpHhGvlxIa+XC+1R
v7ZLj3kNd1C2kWyGWJ+glGHd/c3wkhiHMuDx9kWpmzBb6pD7KlxEq6k8yuIjYvJ/+MwWOR0az0eA
YZWcBLzGIeMl+E5TvudW9ANLOpgeHb3gDDqq/Z4lSGB6yp1xCvmW85gfoKUYg7vAyYxcUmjbKbHP
Nt/VweEQOhEAyG9s4lR4svV4GRxwO8KHgfPlkgcvyAisEsht6XgHEWtEDQHJr7uK+1yNtfR0afaW
tKDujr8pAyaKm7C0H0mzFunt1Lq0PQldd6ThlveKCL/6NijGC3Jzem0E5H18+VTg+4Np6ApxtfLh
ajTno/aamGVU18g+d2UNYO7//X8DmimYHXZ4wb84gPUjG9M1frYU1lm2UrLtIGuSALPdgo37K6WG
+wVC/+luvpKce9TDnpTLX3Sro5DTXK+dBVO6Ek/6+Nq9NtgS4JEluJP0igmwXMwBpEFbOFXstBKp
ApbZmENIHO3sRNAyMPzpUm4ObWs1XajhIhag3e9OmsmI3njai3HSlInOGia+vcDm5YmEUyt7QFBp
fNRhwcajStKwa/MSjRm2uKXxHxeV/1I6e0koWeziDnC8I0XSElYdxQ5+8QLH/+5pz/ypAjFhtuH0
wWWxL9Cu18nq0tkGcnlniEJml4OQf4a8y/HRcjJEJ4y/SKRTK0RJNfZt6anMGUY4sF+q4zN9xi4e
37HomVxtVjdMnpXJ03vVoYLgs165l2GjVvR35MwONiWhGbVUlPJfnjMMBNBMmvD7xLuXr7nEziSC
+dDGdm/Hy7xd7pfkUBHhmp6HtnI33SvnGfKdpzJZWni7CCI118v59d/+sKOcgovOQKlvIea6xiZi
Bb5MhgaTu6n3mluNPTkSdUiCkaw0GoKPAVk+ujPNcuuj4sfpPC8VZuXwHAKB0guRKdwLx+q30u8R
UzyADugHyE1Xw4h5rv4Fx4hHEKOdcwX7ipyxsOiy32GQH9omx7vVz7wMuNhCGG92fBoItX1qsEcg
kUNcLuwyelJ01RSZAqIAG4sZkuiSj6BtsVWZf7HG8ihmuEuI/8F8ay2HuR1FfkL4xwXkfGAoG2HZ
x28ELw3qBKEziSEEMf3mgrpFfk1TcwKydm69lLbIqE0atVjK492Azg7wBqyU3Qs8/SHsYYDgMpmV
2nFOTt2+KQE7sg4aFoppZ0WwHXa06JjrNrc2pRQkDXqi059TU39OAfNPbaBOGgL8q5KDRFSbxk5O
V/Li0Wpq8DLsUWJG00h525Fx783sqctl1BN0nSgPEXCJywvvRlbHrkPwuqekYONtiW3B5HQU8SlO
FnCYJOjOpQqTWShVkTLZ0V8uKaI7LvSPc1mODp347fRBYMxIewVcy7y9Co7OGLhADQuKw5cqaXFN
K4VkkPGpCpusxnjU/5PeSXnzDvXb7zGUV3K/9AbhL8Kh+dMAizR71bmJpXr41V/eF/bebWEeAIew
o6na+y3tR19HyFELNRJ14bM5AOhY3BN9T8kZbrFPryYGMn8KOA7PTZF/XUX45Eb73oVGmiAB3k1Z
1ZRhRUkoHqbOcOrnsCpJIsqkDCGaIFnLlfR99JrCS2G6+nENss6dyseb1KY1HlGjuvhpKbN59YtL
a4uMoXv46+jPMIvr/YwJfRkeNDrc39KUR8zTLHPF4T6oP6cEPuhkAVqdNEA4xrErXLhgYfEqR0Mn
McB5HISFmyalzS5ej+/6RgM/ff2cillHiOjULLIO4wYz9bE5BVht66OQZkL7SXuwxp8NXBVaU0KP
/Ytans5N3r33qK/oCaqBijybz+0LK1RvIoECf072RsEX3ZsFcDeUe0ZHwxBmrBPh9A405E+7MCjT
10eSsz+CrKajR6jUXmlSyXMx0crIbh8NYARrT5JbJsfrnx0LKDiAi/OwMMNiluXpi3ig1qjICYE6
8IVNVCFnsq9jjkp3Aax1gx9+I6HP8taQ7SBxtkEIln++G268/r6EXR+pbm2DkgQfwfOOxR0639do
itfv4D47cOXpcrJR9iB4TM9QjZMHIgJWol8LZc0CxKCigadtB53eLqvHQQCCWsJcP25JGgmxsRII
N6PE5LBjt6osdWDFVc2sR8aSVbhEfbRT6keJKqDIL5dNdZMHGOvVT1l23/a9RUhsS0BJ6LO4sn3a
2KZ7m81aOWxSXUoxV1pVogVLWu0eo2et0WBpahxQEHdMPAQt34eGfixKhTFfoj9XB/u+CWfcl1G6
LF1/PjxTI3SrbsQ6ZTArUhj4o43Ofow1GuJpFoC4fWscsRBB8b2SQb1Ck1w33+MjEg1UUi9NDh/x
noFD2pfeRam2L4ViYfjx4011AFbTHlFLv0PkATZI7aWUCySGNA9Zg/3+kB2gYxGcCdetlus5RFvE
szS97T/3XSQuh6/rDddOnkiVaJlFWe2IZpFx59rRpASVXoAUwLC4nEJ0BS/EraKXur47hfxNJHk7
kFvkOltoNA+k3CIDiwi8Nsg6Rq1/oKJ6g4Qdq0OUxI4JSikCCS/1T/pM5kI0DWLYL1JbHKBfYR1Q
nD0t9AUUYhEUXNwzNEyaze2ripaBs25WvC6V7JoVGFq/TN0CKUliJfCWLhmMlPpq9iie+MEXDTRx
3Pef3aXcC+ZDaE5Y2klt+ramey25wO9KgjOiREEgYNkY2aZQhgX1yEUNKDDfVKzPyEmLk7y6G9bp
fBRJJKfVsuyPDUh6a+Sz6mI/kZKCzoczebW23NkXJLiSCni1TckkWDkTPXl3G91XWDE6ANruA5bD
HbthP8QYYWe9wHAo5M9x1L98goRt6IAq821zCCav788gcfQWAphIY+ZUSs367bFckl+qmwOTqpPx
3sROPm/bdTcYHpUW92u/mtBZgeOVaFiIEhQDrjmEggAz4IKqCfVfAf/PgEPyz+yldSAF18xgRIBg
wbhH8gJjGfvxaKon5VvaKc7p8NaLzMmYmuZWCbasWR7dNbjXhl9xBX1S39r2zYzd1UvFHaAl9fH3
oOB7/jqr2myAH0FryIjx1+4V3ywOob01UyLxhEsLmPVF3iUQ4KTUW/UdjvhKpKvbXjXVcnU52mOG
0VrOYLJDUFBRzajLckyfQ6NoQTO4FksP1leCsv9f7woFYW9rFmRdDr4RE2yvI9Qo9/tcS6gs6G39
UNq7W2DXJUc5DusIFPuwh5IF/of4c1dEVClAk0FOuJXEtNa4vgllY9q8+QuW9QL/7qkzTf+4kZOa
qLfsGgcsk9kDOszVe5tJJ70BP6TLL34nU+aG6J92RqugbFo1MllZGsEBFX3REVquMjxRQy/Ryxls
fN8llBZR1Q5PPceo8N7bL7SjUu2/IsJzoExW/oxsqNLud/U3kZCqPSHOseC9Bpe07I7OxANLW5LU
jYAbRdyxOFbOkCNXaFA9SUwYkQoHRjL1Jzy8oo1+G45zTt+/Ze4uUC+W8BGqUMIhfxvAALe1ftFb
TRy/4oM9NCHyAlVv2ymUJzUEAGlZG5Bay7vCuWd1xjYUEP8ENUI312IoHLwNqzsWZ36xVTAi0rgs
tk5ueQ4hvcaXnd1FO5tGlDfNzAS4dFOvKDQrD7gbAMKhz2G9uAHAgPOLrVcSjvo+p1iTR9Mt22OB
mApyc0SxHajG2m+nJZjnsUNq9aux7V0bp+QHzHM+Z0ED/60HRGqPSN2h+e705xelZJ1H4a2CtMar
6Iu88Et4VlPXFy6qNF1Iyfg/Qd4y4krCGVw1LarR6P3AoGk2ODp5EuwOg2IR9J+bK61fqBo18Oj/
QOpvHl9r+jhurxpe6G8t4GPLeyOx7Uhk2eW/vCAyBbCuLltAtjmO0+o999dF4m0ClYJMmCujoKXO
RJMO47SS47nT6AZjvI7MvmAgl2mlXXfcCJLgIpk0UzDYuryoDYETd+YSePdnFZ+/RVhnbP2v/bt1
sM1I41vgXD9oIgpZseBaJR1ozAy6EWB/rNld2+CDnOGZQzs/lp0XzRkH+rmdI6vozfksByed9Qzy
zpFyh8CUTSl2p6lQKcIS9uK/nfSFTY2ljz3mjxM0yiIig1D9h8MSuyjwuhwyv95y617ONsgWLHhr
j8V3OKrCFjdGZqi1/n4Mka6koNCwdM4z2jRTDBm2bS1kqBMleTMpvzwcy4bEaZrdiJDVTvlWSNZK
EOWoWAcWqoncpwWEPWl0xkqIrjGeMptIZEQktj037+0RfKQ1FTpsetUYs6dxsnHFIgRM6lK1Bmgx
/poEgxmzCb4JOvuSxaSouqHIfLZb6I2r++xi4yLQf9sLzr7stTe2Bmv5LeC8HNvK6/SrJ5+n2Tvh
U/W8bMKgD3LXAUfwaAw9Jx++yVE6a/HUnwjODhTS/4AQi2QKYjtAiil++C9QRrmvgeSj694kYdL0
O0X1zzY3dpOVtvzc817zIhiyHQ+H7HpfIcF731gJid0XyGoD3Va47AdxOiuuAqDMUu2gGrYM2vIW
LXJn3xHQ7VilOQWXoOIQ9NGxH8xDlbwP2M2q6Ou6b0mij1+W9edh28MvplmT1hkkvEFpb9ZYrTUM
y5glDjb3Q1xb8cI4JLSGnTc52fs93T2NerqZnzhy7Ru4ym7L1K8dAjhyESxtzM2Buhkx2hWtR6C1
E4bV6JUv01eu4St6uoZ2Nsd4338Dj6/a0oxPBN12P2S7JyTO/gS+Sn8xHOw1jeTEw9CGHzf3RaER
8oIMpUMAbpOA93Q60hs9wld+WaxnVcaOXKAIQewpDJ2tQqLzJ3RkpTHVCXH9bcuZcgomNH10FoLG
OIyMKtRky/kAs1evkG42n/hwU8cLQSGwX39trbnalX3AYU83PMXimyBOAfd8VolJoj061JJQ+0v5
VmZsZUYsMqlDw4p1eCnCF43NKQqqQAXz/7H9bzbDuKWAFPwhdGQZydN/6HBbVaOX7JyLrY6JsWpZ
g9BTEl37VnHvfhJl7NYrqtF1/m6DpFassQf1QdNwhFf1mqIR82+CUmQdIeKQ6CzB+Xdr7b2v8PVo
2FoGTNPSCnVsm9ZUdiYR5Z/abaY2yB6r2xWkdCnfpL7eg4C4trh1cmroagqT+r/yxW3k5n8kkevX
lTANL5T3rIjhIt+ieKaZBsMkr2X7a4DAx5WbgW1qdeP4Q5bL+cDEOqdkOK3SWCndoqB2uSYSkOZW
g2KfY2MxPs70mB1KfOYKG6p56iPoqHktj92bKHNbA4r8jlhvAyaHk3bbzZP2qAvLb5/3+PHx6qI6
cIqFw8xu1syK7X2LXMoIRgmPdgQhYX76a4xdu0fypWWHvJypD3GCS1W30UgJS89zAqwHHT/iSm/q
R8OcPC3LV7x5kW6wtS+zHhD6bVNMPkeGOlY5Q4K42SjIhBHBwO+O96aBtGFBDRJgPz6Nal5duNbs
jzbenmvyQ80iDLghrfTcWxT3L6i97F1EIKd/0Aj/riKJTeaszyTRRcftxxr2th6NDyfp6liGRJM9
+tt8fuT92/qknojW6wyfYQyuPqCkEsbTe44ZaeAQU2snMeXm2UzVr39oZsFeS/8EjfLIqw8Gg+ON
AS805Pnm1/6HaXvtPI7NAZBQv+g6z8jLTXlhKVK+WWuan06Fs0P1qCT2iPp963rjfC7VEuU49XIc
F8JIluEKFW7YaPwzxF41Gg3EzwYaaCAFqhc8hmk6B5fh0zlrXW+fucojmVVvJQm8iaFFKpnj0eyp
GjZZMRnmyu40kqVBjtVZ9PpyqyzlvtM8pUoXbvNVtB0QWnhMGDqo9+jCsIbkeC5E5FlyJxVgFM4y
aBx8xAIKdLDwBJjUVrANPErV3F4EzyyfkmSoTys3ji06THZp9mV4WvJNy52j5QSShkXl5HfsBWzT
QGtGYfh/UZPcGgNo//l+4GtI6Tj6QTPzb26A5VpE2oTszzei4bSsAfW2juaafMZEYiwY2zC63SZ6
uqzVpZXxpLekl8MUEosuYgn6hkVxAdOxDI1Wkk/Zs5zfZRdXYNXDw+pe7FrKOkziF7Zjv1z4WzMf
ymD1UhLi4/JOGlpYhesKZdNanQF5XcGAjgv/SY5pF6zb4QSU9xqsAoFGdlVRE6nbNUQ473PlrlFH
nl1BSECBebqGbUmwueh5MAzg0TiXVDcSWuqujcp/vG7bM66qHSJwMQc0RCmA+An4GHkNfI/Bl3UB
RrcC+Ge/3wZargb10ZddEWsCH1PQQylxlHGz4je39A9losfobmHQfYg2RP0jP/bYuH2zM2XeDv8G
DJKJ7QvbcmITVoU7aLmogoeNsg5jUbLP76K62kv12pHUI6U0/Y1HGzeR581oGqvNDLpWz+DztBsQ
N24VufNnVykGGWkDrXHAYp7iWdqOwLscSPmdNYoMnkgQAYrYTyW1dawH4JOfl5rJqzVSKjwtAsku
DKLoc/KK405TQFxAmQUbu5ZtfGf/ja2DSaPwfrUmpE/hV90Srwd4LYRxjzMUURdQAA5V/tUOmzem
Psqt2nuxZs3mOxGuPdXu7KgKE1bFSs63gBrOXTBoDeCMCREsqzq8sFQcDkHmo7FSubM4tg12dCmZ
z4RcV7HyLR86d4rlE0TyxDBIDuiMC2XgGnu6s7CiinV3H9HYxkBLZRC16Altob0Z5RxNvg3AJN+x
zxlVbjdGAEqGPjqPNmQZGYd/8iK1sKCiQPRoV2eQQ9AvnBbC3GvBBlpih2rDfIJzunSx4BfMNaLk
r77tsOeErgIPlQovz26Li9fTn6D7MDg9eS6TR16xGdccXB7BTPr4bkXWFoC1Ev9x0+uBpZjY1qec
8UXLxnqegIK7/+TBGFbSWgSDTPio9AdW4KSHK41+RPMBxjJGvf6QpV2gPmhBIZ/oj7OiQChANPxO
42BbMZyljGQL2hkJyKCl2V8G1opbxOV+YLaGTVEXG1uRXrfuKLn7FLlOAuLhkcK4tipEPmzvqkYm
UD1GfqHBIxKRs7t8yG9C+LCJ/jKqR3YpliCav8AmDFYCdEeYTmpLO81RCqVpUobTGn/diViBpaat
NGethc7/yS8gan6baWkdpXVjm/asK767XZM4f2ITnmUJMDhpRUjel0DGpNgTtHX4jMDQdXXmL2zE
Q4D5zAVHlwz84x7ZGXFDsoig8yc0fWmlB3oGJH4/HfZvRn2lV1fCEQSYGEpAlzQARu39Qdd4wTIz
8vbMqAMg0VQKIR6NRVB5gN1HGgcEzs6bnYA6r/xbeq6lHWCYT3VR3TL9TBCUvTwQHOT3W0PTE6mM
Y1uGoB3uNFgwDub9NwJHdWXme8x8EbN26Vsg1YtNFCwaop+OCOh4gHum00r7WPwS0+ltMxSimfxH
VYKYabYEpQr8JdXBWhjAok0Y2ZJHBP8qDW4wmciGLiYd+ZcvH7GhTqafpMLA/LFME8j056VTn/TK
fd4WS+3NfghqdVUa/cyYLxQRXVnO+unE+dWHnAhI7TiMgGBnA319dV7aEP2h77ua9nJetbJMeRMg
EL4w+t54LjrWo+HTezQgucUDboFTcNmmJ3fdXgkHVdXqHhw1p3ZGIdS9PI36EllS5d+zqlfg5i8l
po+WuWDHV8BjwT99OHqyr1/CGhaCv0qCQQORxcn5sNXSfuZhqdBa3FgFFydg5WlKmc9eDWlkthTR
o9NfzJ56b2IxzhJFOCgIogIaV4mpoapM2oZ5ftGdUMmzWcerWb6DN37qb6Yx42YWVJKwrF8T2xoT
4L6sBJQ+6oIcbS8U+m6S9NspR7lV/LBQHussmNRyrAO1uyCTZids0VxFqZ3b/fK5A2yDYluRyjqu
iS9ycO+C8Y8W7hLlA4XBRXCCua/2Khclc0KIppIGoJiAIbNvFSZvFAlslnBb/6ZGsV6dxzG3nX8i
Q6RCY6aagjiP4fMCd1SYaryHy6VKwtQqWty/JIcOMZ0wIpdrCY78qV/6+r9/K7YhC0y3Y3ivGq6b
L6rRFeyoqSb3fw0bivlO5ABBr6KLAZdu1UbPB0ROz5/ANXwmgojh9B22QixyTlb/pfLouv7QmBTY
ISg+xkqeHRtw3EJyhwBeSgZ91PESe92nla2ECY5sJ5p6zUnWT3bP/l0FCS1xe4E41m0Wksc7gGG+
EH+ptRXnSZsmwCp879ABxnZIPFr7WYJhX+JK5BqPXpM0UEAPrhhi5/zVtTmjgHmXUL5r5x0zloiE
wcR+V4Wh/6+U+n2DMqRdtmxspOr3/xIEZ0/nk797dV5A6ty/PZT5WiUIRnQdcogqedBbZe5fhZT/
DfDuyNcZNQFH+AvpwZaFYO6RI2riSbgZUQNRKLuDu3MBJ84rxK7AIpnkA+FNs3BssgHxvUBmXMde
4aTp61n2QK+dVkYSQb1YsOV3kDPIjJh7F+h1+/jP72uigQZQPS/jdtVNsAeM+JjZCBbyGHij8y0t
Mv0BJToZUb9U9MO3AqDn3IRBVlmtqGXyIaunp4nOEkB5K7OwFf/4pgKuarAhMGo7E25R7xwxtwOy
goif8hF2dhAED7hH8BDktHRGGqLS4m3iG97xZEG9aQez2/PdQ7vnKfJrK4zAUrMOrOE2NZbSGvf7
fVhFL7lisabkKaRKcROKFLlFs65/3Eyad8MVtZo7cOf0VdnmeRoznpxhwKEkOT8d8r9zEmC6CF0w
JPlL7IQcnRpifCwnt1I5zuDqbtlGvtWl46ROQVYv0Oo3OHI6M0WnVhCqFAJmgWzz1PvelX7+jvEP
hCCN9ehv04szRcrtuUOBx2iFpYRQrveYjUuFNbO22mQ1leuU2FMt2zrar9ZA5hbZDdlmm6UKAJcU
MGv6Tv1X22gY4xCge03zQp657rdPggCu+sCDyTjnkqkUoTrUEEgypRLpMqs9xTUosY3Mz27+3pMf
KxZjfILUpUMS3H0i4WDXsVArms/xKvlWzLy45qSbCCqe1ANJlkMio65paXlv9SHMye+seo+3tw83
0oyDRsrV4Qd7ra/qO2fqsKOzMYk19Zf+D3LK17+EldjDjVwKj9fCnxE9dJOXNyivU+XSO3ZAxwdb
cj+/M609VqbU4hIMGbPH2wjJ7jf1EPbc+IaQujqOSWfpiO9/dtA/cOJrycjC7VZFyhnpnU+lyNc5
oRYBb6tDI1i0Du73OQFaiKJfRj2I7nDA/5w85oDE/x0ReC3fXruX+9WZKdAvrNan62i0LU1k3j0h
tlg+Nfj+HEgyzXSI5PNcpnU8acEl9+xvTNXLmOQJDdeo4SYL6HDwyYWyokRAOIDJJFHkmxcr8rs2
5EXBw76mNxYMbstMd/N9Nef+z/GWLCeUNYSo2dMxrOpztl2MxqZ4dxqEfOjLNkIyREoqyNmGn0xR
CDm269OXo6MmMd/cduJ5FDiAO0Y6BVZy8v94+Tc46a9/uBBhOJ3YGlkDiTd518uLVN6dQ2l2A3gT
bb7y2DF1PObzKzNZQd1VAmb+hUfQoeVdTMyeUx3nq913OoKPu16fljeu5BpbziYJG7vqXEHQ661M
oTnGzSJ0rVR85CmLBZ7QRvC3Gj1aHvQdwdsdrEUhrNrhMW7fJdICR0drq6vaXXMY8Rl3NfrUCHNa
xD3jN/53N7aTGrbf9er6XKgyc82uIWeroQA4OXSnSRV3cu4DNk13eMJj211Rlmk7tLxeFkHPeTsC
rV3PzHxEysegorQ5fXItupNAkDpR68FrKFhMkhSqd0+eY7ZqV/NrZ/CRclKBzV7evdHIqJcSSsMl
XY89DyQRnDGUmPvXqsWGxndYEaE65oh9GTnt8C4l03itzCJni2+0u4395IFyej8hchxZbxPfFppM
bPek4+RiqXE1dtN+ZDaDpLLnLIHOfzhb57f13KAVSUKDAy59p6ITVSLWrqiEmNcaxbTUsex4Sw01
Kaui7HAAEoWeCY4V0joAecKKTYjBIsOOTEBkisBm37r2/KZ8qhTwR2eJKqSYGBO/2WuNLppwypLx
ZRUL266EHxhmHYmjzLFV/7DaE9ZvOdhr0Zj52Th8n2i8yVMD3LeViu2DnuZTEkieEibqS7Txks3+
lQODGTDyUMS2Cr/+7qQNNmNeuSi8hxQPD/E14daO4qNNgzMxgHjBsATtHY5H2E6iAnPiWH2oaHBO
bJPxQE7ApfkxxRXFVj+L2JU3S8MBg9zBDrcBA2UpUY83VwEAyp3cpLk7PPQKToijvfZQOZNMW+VG
sPIeZagj20TMOTfD2tDYenjwuHwH3Twu1lhVFVwFjXyuf6A2tG/ItcCOrAQT+CFIAHG6pRWhIe53
lRIT89SKTFdHzePPdFcvfO5G2h5oHXH/UuYu3Y6V5LnxRONdBeGBq/EFTPj/+UKaNsmDvjq6363y
PYZPmaWvXLRYDvP1yFLxSNcR8UC9Aa9Gv9rmksfg+t770oXQ0jI/HGf+5HY1ADF6RaYXVHhaTNb5
9cxyJNiWkLa2Ml8t7nJwuOLrWZbgxFO/gE5ZNIctztV33E5WfHzxsGC7px9ABDlKa0tTSboCamFl
1k3HFIDzMup8wwPGtc9w5xg79TKVqhXOzlejJTr+z6ZakgR5aW3dQ/Krw3td1BzJ3mhylQqOiGH0
Jpnat6OzMMTrPNxR7p5RIsHvzJjlZqMuFFQyr++aciRwpzOH6JfVO6e+HvbxOq3D/eFYgf5CpQ2M
YyHscOn0UrjeZuInbc8RAmRZKML3kKnNdYZ7JclSe579vEEwFs4DcIu8GSLrHbNxgyXnrxKTN8v+
WeiK+UdGNAdSd2MJEWF9n67Lw9giKNMMO+1CTVloJ5i55L4+slpd+lNGnkxXObQuECwhAJxFbilY
BzJZwu4M4QmbaJM/yURMMWru0iCEjEAZ8LIIcz5/wzEiFou+5RuKWeuFNfZS2RxwqXMY8jnHmPgK
AEuRx9YDU93CiAGYis34ify25yLtT7LraNh2X31vyyCC/VLcfGKIcqAcCPKueJSEZITaQJSFtCxh
rAGNEslV1Wmjzrys7U2JU/ExWn11T/XOttDZ7IpCsbrG3Od/8ebNUfNTSsR9y5zr8laejL47Ctre
5WkDHsEOyXWS8VGzusBSVXKr4BiybZMNVL947SYJWJ9D6F6CasmwBjZGkvWtZ2nM+Cf0eZ5/cmgB
iDZDpXQTbH6Sn8dOfRuwYJ1j7GEHy2dyO4eLRmEATjXR4fkIR68DOwZU2VyeJnYK5IeLtNw+ELiZ
CFN+QcENu9+4X658p3E1EuGsKcTPbyUghl4rPWMMh/1N0ENR5Fw6dLss5Nbcw1/oEi6BoagfvhO+
eBJWtRfR9VTmZuxsVXDI+KaEvWrQwfTPLnR5h+7DOQqtNTJhs/N9rHe3qIQFjRxO/PwYSnD/vmsG
Un7nxVIkFRYQbKNLr8+6dL7t+8psNMdsCm7Vhxbnu75hBu8clrKpST1HzStRUJ1sr6LfCih9PTBN
o+7tQWrxPpupAZNwiwQZScV4CZK6t6LqBvcUaRyTA/uzGdD6mtHmNNeo3PHNqiilb6vLBgqz/Rsd
Qscpyu6ENjbHXWHz+X94vfiU7JlUAqJQtjBC10GHd2DbxbQQPNglO07QJ2VMPO6Lqu3F+dOsXJYj
pAYf9yg9xgMrhhiUFsRjHk6hpd0A0O+8Y9uoHL72HpGTWfsmn6NI1mEcIjDTLs98Y0cg1ir/3Uax
cM1xbZb5HQTBb8Xyz0fPA3SOI0mdHllR+2i3nD2ll6Jo2YYpgOksHqh3vxetDiZnMOimNRirDstX
1zP6hohSdvA8UYGU4On31GSlFMIrLh6dTmOZ82WpnDRW5dINu8sPaCDcAgRlKMHsENZvZiSA+X3W
5MIf+ZzyZ/g8l64+Udcr1Z55v0Ve72D6bD0QiONr464NaTBFBQKhh+laj+NLtz5dRibBXgK8aEOQ
AyE8Cyf4kBqSWStzMrFbSW3mmaRNQvtEtqAbtFxEkJbc/OonijTexJFnD/4QuXbtB1f+Av1zj3ae
9GYDwgjWtkDR1MIoIYvjLm2JxrRRU2uVyLAbDFUhzBTJ0R0v34mVI6EeOUF8GGEFSK3dJkNOD0xr
/c/hn85izfyX3ULhUn5K52kAxAHfla+oXEmb+mgKRlH88CHY+ano4e/royl/7fPUNNUA6vd5AeWe
RiFnuVel25HUpQEFLv5PWRAmj5VoqTV4ePPbG4kfhSxS/hPah5seNqe0MlPL+lCPPCMh2PIQVwcZ
J3mQUsAUn46qnTdWzi75kZRQOQnYMGtQRr1gtRpvvOLclWlyZ79A+v7yit69VotidrJt+eNpzwac
jJDs2jPr8dJgOGtWK6DzdjM+xC9H/uMnexHrUL+mKXLh9sch/L3hMb3ku7sGR9bSOIk7qvrD2M3M
g6/XnBb7OlBWumqBn7c1MpOJWGpvM7DbRCAzTXQ8CLry/iMJvmuwXwuD6WTOqqeSp31cFVLcr3PS
w/Rzuj5F5OjJOmc+khPnt3Bv/R+T6cmnmJZ1TDqHhbQlhXPFjc9ZRGmKODfpx1NAYFpDspXHmixh
tJ95jcKNTdxJ/T0+Fyz4BlMERtIWy6+sSFjhe+RWJ2W+sSp+dqbxTu95y2OMQG9GH7q2JFxTBuKU
J57buHiqWUrzT4b4rL+GqohO0wQo945p3B7+dw08V6Zox+hY1QYopoE6N/kxIaATpElLD7o5Em9w
jjtu+ksILgnFjQXAQ+zabCMNAVQ3uRf5udpnuKk5QaK3E3m8uaMUNWjn6A47fwxxhanzT2Pgzdtq
mFk54rD+Q4Po9JQbSlYMum0q1HfkrK2ZBwVLj75ZZ7jBZ+NIwiUb4rGNKjRcY50UGTuRAdmkBwwc
DM9SGfGyRUvlUjcy7rHCJGinwVj99hTPTP21o8zx5idzVy6A+rT9I2Iy0J6H6R5FmWOCDuzkvDG3
i0DtgEgeowY9no5BD5tAk7iEEtgidKo1lR0/sbX57CjWLKqIbcje4FrwVq0VeMU5NWe7MWpyAsCm
jnYTvCHn2pQHtjOz1TP7SW8IkPR+t/bpX7tVLYbsPMhYvu/90ATmYRJJuFX5eMaVV21c6zcfeglJ
NmLlUMhgH/ZRYJA6xT9YFs6DsA/233mcEjzD46ENh1z91t5VWA7AxkememdETzWzp+G3INwnAoWv
0w58ilEn0pAd4UAROF4DW5ZFSwRXwOBu4v7Pu4yAV6+cUVxXu41zqNLP9NI0s6lXXeVBIKcoFlKP
PMKSWgyWUM12JER1A/uFJw5CAwQyrEm4gRZdchl05vqCqQC0EXbXTXmf34LkMm6tC3ykZ3fIWA0M
CZysQ5daUy0v1fluaLHKJ/4Rk5bzq5HLT/0PN74IKxS/FyPVIlbBY1viVLzkFeRfIKnJNzL2XZ2C
tAi0bHsDFNKSkjitErHpb7yGalzNlJ5ewIqnfhKt4gHLwoqKMfl3rklVlbqsqWnquIKzsEmytVxm
MKQdZXAkQsNVWsANwZQfjln83Q+Agbfbt9WsHfB1kyNkFxhYLrE1cDzmOlxcFFiXP6OhpGn7VSns
CNCH/AzA0/EniRXzOkiMKLNEZov9hTxQEphoXev2RZnhIyhuGSajJOxaYzdvuK25Jh0zqsfgULrv
nIiQIi7mUXMXRfq3gyPIOEvXL4/xFnN4T86ROo8L780s7sDo3G7Nu6KsmlTUfO+WUuNEM89o1P13
QrChTDFqDLYe6k+620la7F+lM6PGC+CBIM0V/2Sw50D/SW2HdR5P+1U0f6DPmyITHjlz3CZ7xH2p
QxzG8aVO+FEfSQzl/4QIIYmzanKjKSul0+Gi2PAs3M6lG4zGaqO8t1NueNodVOV2riAadJWrM5r+
CV3GQy2lJ+3wMrGc8n4X6OQMWykecbUbEmR6KjZiTlBhtvlZ9Ax+iPwBAFhdpwAA+r88XHFzoxZf
M9c8DzhGH/IHIKpQOhsm0piknvBAiZ39ZIlwD25kpvwHa/HqjF1kUfgBG6qRFo0+rQYUxXXhTlYK
Y98wacH1aM31W7++tmI+nGRR9Fx32Y+/xhXGUHV1eI6L9ByQp96tCYnIQ9WS7KQvInzE/W3KHYZj
Q+ZWF6F/7fc6n3zWBK5pF/ms8LzSBTWrCpSuFooGlFnANEHHGuGAvmNFaNiY+JI8ZRiOSGuHhwGG
tQodEjFsxERwMWFpemGsWusunVmtCpb4S5ZClIBGrdxGuGgQCfi/nIG4ysbT93WWFg0pmjRo7nmd
pQp4sFtN9cMDO4lrk2vFHc+u0K43x5Ib+QL4X6AwhQK6oHOgaAH78Ab/r2eh5m3hmlyEl1iajuef
tLuKEzyyblKhjMcd1ijKWqW66cMc2hWqmbIwZuwohrgvrW5ei+jywwAjWiSH6uJcQ/ThSNXz0T00
JeaduG139bPE/opv0pLyYdibgR6XZFEdMEBpVw+P4cCDuVH+peUJ3YfvDRBmc8HPuh0zI4J2nq4J
oYI5ffBLI9Wbf49RxyTF6UvhOEOytmidwmLp96L4d7fCyc+vKxCdEkYBGcVn3EobXN7rl7/bG6v3
5S/Iqv01E4/e0Xg5GL0w1qdKEiF/z3L3xDqzhNUPMGxtsXId+lbzVKPLAr0vTcX7ike1KOcOD5Pd
pXr1e8mCwZbWz6oF8GrNXdzg5AyE4E++uHi93qmcd/0T9E1/JxsvcdHuHi6wGthhONoxcCZxVzBg
xemOcA0Q0PhoNKyU68ahqx8CYhvlz3h3eHuXp0tZPd0j+Ll77zqV8d+5u+Kz+LsI9QIM52VH0qvc
7YGEbIcfF1Pao2iRoa7NWkOcp2MeF0fJ4joQC+Fp9FDDH9tLsY/AM8mw94injT3E9jS1kxlPuH8u
O4WZBhEnEH6NNoAR6iDclQ4wr9SksUO8JEVRIujydZVpZeu7RfXfDU74wywaw4IZEv121HCjIS78
+9EIHJfUn7s4mFgDaSGFkOOTkYFfEWkyFVvHZUIvLCFmousiGB1SeHsoBQtXH/ydQfr3uwSYFCaC
xzVZKFr2NVpUYObggFKBXiWp4goVRerzolROhG+Mxij3ZGHLiN6z+cfjJCkihG3OfjGgu917ZL9B
E0OOPY2c1d+8Zh3leFGMqcQk0jWNtkGPMMrIoXPWlj1dsBmPXC/CHx08dzqskFrIMX1dFVjWVY3u
vXk/6QGrP/rcs3QRdphcBaFQ+lWwTu4xxYVxqyqg54PAl6NzcE3L+qbPiXsTLTL3WQizzNMmMg5A
10Y0sR+6GLYTEnugJXJ7t23KKKJs/nRQNEXxBMpGzMoxvnlL9eR6v/E623ElUfveFqIhENAnl30t
LSyF2IxSKi89xlmzR/L7eLpghf2BX21b5qwhjwQp5zVP+Xpzt2IYdiY2s4hN2kAGHwIFtdtDrmaF
pVMQCwjOizyt586Jy0kEUEJm1dB7PBF6VnBMPgWEO3SXH2qhO7fxOrx+yXGzqswYxEORSnxnQVGo
m8x8POKVzXBGABuDruTkWmV2YFAfZ7M7BuEtg8ZR4bd0PskWkEJK+i6NL/OKBhAos48AuMdyXsP+
Jp44VxKjVGhaylvJNr/xIRta5Sbmt9/EV9f+9xfujETcgwbRf1TnWqzRcUNxkd8MmX2pBi7JdwCT
w0cjJgXcIhnoey+Ve5D6eVlbdFaeVfZGXIda4YLWDpcB3+S5iiVcc+X4cQES93yEdM96mZcyN0q0
Jglh96igv8GaANQ665tp3JSY6dey1SF/BPbMwJJImi7YILs6szloDKS4M3PdDTnEfbtPxLiOMUJU
znIYY9HYUNsYC2e39CGrhemthiNyqRK6gcESidrMK2Fr6N9fqEV7v7AMp7U2fZBFEgVktyidSTo8
jkvYbN96Cet1lQOKj0M1/WzFicJJ/HurJ2mXD7jZCx8g79TFCb3qiXd3LLUYWiNLRSyGOS+/F8G3
lDZ0SSO/xP9StjEWrS+B/eRMM+kAeRKlTnjNwpEzlvXD/sWRYR588t6GTwa/nWg8J/4Fj/70VtFj
raFQu9WMiE5uVy/YNeYWww83FkcOl8Q4L2rN/b23zHDz2BfXqQAWY6cZpXa9hmlCZUcuOLTI6lAW
kUlqiCqvBL20t0ghvPFdR1SsbYoPn3FN/ZdGfLmbGeBu6DMzT6UvNfj3B9he2xsC2ECwdIe/9hSd
FEKM4OdLA+CnFQtjmPMSoWTbEnzgGQvXYgCLkqVTBtcER+kRtwRNv60L0Nf0SWw4eU0QA4u+kiZ6
+M54TyR6FsHqKXLOvJXfLlYFpxWZpqeW2vnfDSImgejoWYSgKv4SNzJWfRDE8WEyYp+HP95h0JDE
0uqv7zF7ilcpi90H9adn5YN2njAUsoEilXkqd5Uk7E3Ic2wVEcIFH5uf71EcqCEXUYsMr0Jxjl2E
4itq/FTyDnlGSmUAGuZbGjb7D7M4jUTcubYjLllqkc8zNvL1R+jucqZoFEz7e9p0xK7eOW5YEcOl
s+XDtPYfiSxIuM+HnrQUxvseEkKnPfsKvz3AVS3tNBFNi24VRoAVtRub3LK69Ur1ed6ZfYakPAKE
wKDzpDHnVLJsgoIEDOxGwazo/K55OfdAG1+XaS71Po38oPLq7/Q4PknrLHl6tWvQzTzwgg64fdcM
cMdrVy888eYCoTLn9Ymp8nsOvDsOZ2k7X1Bg62y6DQZ+YjGaUtDwLFfn8Rx3dBoTxFeriD9fER+3
i2zzaQpXGxa4tCVw7TBAhLeIWU0FYozTmIKkUccoEZrn7tJDgJ4IBKpXXA1BWHRVQZgYvvWfabeo
UWMxigUmoz1n56IIC8V537q+aFJ3jYH9HeY9DlmhpyR3OWB7zS7M052P/v2HzIdTUak6Fs9OrW4s
t7xI8SFFMoxrRiRMAS1p3wEfR2MMuKG1uClqYzEcTYs0Vzx0VTzpSK/Y+qsObXiyheOswMgqcgBN
xRG3KzzN6jg9HWN4MTpJakNADpHclxptqyjY9pPW9O3yzElmxDYGnsnUmqyK7kUVSBEyp6gi/0+b
35UhQJBokvBGyReO+3rw4EXecZibzk+ElVE3g8BosVJffz3WgSMLDD58s4s20fn3A2Wx5Eu60vPc
xZs8OR2oXY0rRqVRYpj968+EGea9xbe4iGOSF2PCZqbg6VxE1Wm+Qx7mUpKrtcVVDczBiNmIlUg/
ZZsc/pYuA2crNaIyUXzioX4UlJF3gp3J/WN/3Xt6VNdHsnWY3jb2eDtDF0LQ9Ikt+oU7NUlKgndP
Uc/xMrmh6vj2GhIGOcN135AHoK01QlZReA3qtkZZPnQja4ZhgnEwjK58G77ePHFWJT28v+3rjI2b
c7dONRrIFxqSKniNYnztiDFydy+rlpzU6XdLfDz7mt7a1DUzI0yIUEy9oPDKVMnwDlauI01Da/VJ
DkozwQoQtAOnkwvJ0Gw5csYqqjnHPtpicMqfx3CuSeBWSh476uSQw9gZnxxEye2s2jfLymiyjc2A
H59gwF7A9xEKRUa2lZ0t9uYHtiQ3ARkpcDF9wEY+yM/NThamVorL9IlxUKlPLXUZk5Nkyr+BzRAp
sKC53dey5UUTptOVTXzrBnjDtlL5Gd44oWccPURowWD+0y3Yvuc6D30h46+dlv0XJ65wTbLFLCDR
Zu1fQrSE6FWzZjuiODY+jPf2JsPWAhhpPljreLmezONxWrc3xbeDsYFMLoj9zu6W4Gm+/eTGumqB
Skphw/PSO5CwByHyQCgWPznUXSiVJDxgswdqM4q3aO+eM4RRiQcKm9zFO2DtfPqkU338vI1uqCqU
7BLp2cYbiwmooF5Mpg/wRSnl9NMI2rZw7gt8qXZGlI9X3C21AqrtfWpclozf4S1avkpfnHFdze0/
m49P7YxRIYxeB6vpYg4Z3XaFRM571+4dWuPccK5V7ixvgpNYSwPl3b+WEUr8+5D9Im5OVI0/Ud53
op1rRzawRexTqbJWFHbsVdcCiGI/kht3oRFe0NpcBG2Met+GHh700azFkiD8sVUCHQIhNby/1jn1
GyC7E5W8wZuKIzNsLRzrY1lCPp1DiDj9tCLgkOHe6saqkis57c2LMEFh4mEUkOWYNeRcx8GYN6oQ
WJ8/9/LIwqqmBwdHQp7fFp3QM6Iz1abCHND++2EUXj9d0cXidGkLD4veSP8ccIgrc09xPFXykVOM
B/v2BUcIFIu+vxBXemm6nmLZON6h8gbQLbrHf/UK3yT0pSQMmIN/wsFmupS7yLIscIitBIu/SL3p
l1H6at85KES7Ppp0An+M7gxttm0qMd+EbhP1pqo3Pom5uPAJ7Ua8PeyDmjIU6RMGoWdPC9fddmX9
/AY828rIh2X0D+qj3dLqIc7g9h4fbFhhOVkNxWjk6JOe5RlYkf9clgvpYq66EPT2HgFR5DZyeefi
x5URwZYsQso4w5bTXtOBLr4nYXw+QdTrOaJkQ0+uzTptN4bexF3Q/5HOUASk3eaFtmIP0XOuW9qk
LXcJVLzX9pYEQg3f2q5R8EWBRINuysOugs20IKy2flTDpLCwoFCIKclLv14z9EPks6JPu2wc0LKY
mGfvuRQlCS4zybdEsSQYjpXscb5dvQ4RCbparT7Av6TPY466k4Nt0EHsA7NA2ck1udxVDtV6B85G
17obfODJh7GPwnM8LsvIZfAJIAEARXZ1btikF7fJq9NNfAqkcOlK7ormKu8IeyWw+HNpNJVNxerF
Amy6uFkF69lGh/vPyrtrhefI5BGLbOP9j6eLUtAEafOP69GWFK7zdrlFFVQBoo684HmOHziq50QT
JLq5S5/HrN/+rD+h87kLf5c+tVjf7KD3M/2GVFMYmYe1n0B1YIEjM/3A/wh333ex2hESMI5vf6+R
94TZFJiC2uPwinyZInMSSwU8r9ZgLw9DlN8WEjuJOEGiDKvbxsaFu+d1ALCGojNUtupT323ojS16
+yqtio1Rnt/nURuuLhizB6QcRg/Ij2ll4Jm1uR4ezZ+lkAe0HPQ0l3WtARrv2Gfz+UX2hH2xNYJa
eqtBiBkLrPnQ/snE1j04kieO0v9a0Hft9u7FhZVnT2LefsQ7jHRw7Foz0XwDvtrzbA2vaHJ7dupt
kjjn4LKedjEXlKzI3ugV0hTEt2ghqoVNQx+PpqQMdgLHR5C0+x0x//4SrmvyOtztkeOeBjbW8jIP
jkiRES77QqD+SQObc9LTZZkopDc+lh1FDilKOLcjYm65xgIPWN8NB2fO/2vka/1tDhVfruHBGIuy
zQ4FrOpqTszyfQfUylZXLN1n6jzfE3G1pMWDoZqSuG4azg6sDVBacKycU8YScOOXJgLV9aDIWpZq
eR5Ls0Sq4TKWSdL5TyjlrZCo0DpbbMPSdNlYbGawd4DUoeHtEp9QS2IGYy/NcTjc6iOvWXL5wzsS
RwbBbMC7DzpuGJl8h/PhykgM7ZlFLTSqtU10pgyUpdsi+YzVCv5pVIz4+4hiVjQfE2hMBhNtTmEp
RIxhj7KiYz1XZKCRsYE5JZoKWg86RDoHJzg9wzDt0lQPkmfFfgGJYJMPgDVmhgI4MeODh0N8FC8a
ETaUqyGeAH3CQSGV37j8Qm2kGFdkBXiBVFADGYxYD2d15F1XhuNEmRBEk5misH4EpEf721UZ/EP1
Vooe0FwThbByQNCOWwYHgaXwePEqxEN45iDTxRU0BJpHM0PSxyes3IthuBPbsiATvdxn5upxKLxq
aWdZFhgKzfe/Q+IzWc7iWz9/FoJwZzikD6NBy1Dq/5I4w/BchfRzUg7cpezsH9w5D7Sbn8SVuh6h
KXgwBIn8+bASFuQq62gAkcSMlg0rySh95esIBC1n4OMBBDHIr2q92cQEWFeu1iGU5lCO8ErILXz9
aA/RV8qNkf3gUWG5VjG9ytOzwrMKPM9kHaoMKXAwYD3IRGOVjlWF7zq6tMZG62kmMB8XUddQh3fM
Yucd99b1AURwqLf+4Kgphpx3JMk2510kpHCgHbjEpZq7G51heuZsBvtkuwVsk9Ta7ivkclppE6HH
nrzW/SCubtQeRmbojJjJnj9dBX/UHHJZFDt9NKRN+O/3sIo5keIxVTkbLrWBjb+XM06NahX7vngE
SNVFP2Dt5Rek0iHSEZ6OR+3eSQo51mDwkTNLvIIlPAI6+R6gYSD+EPvJ0yFZ1b+azRlExxvStpOO
20EXOb0Fu/7l6vP8CAR9LfWTMvXw46ABvWh8v1Yx8W/1+6Oy4xT6zuQ0a6vtl8T6oB1LSFtGjGbM
z5MV1gaYuqE1mrii/9ScVVn0mtjHB95OhDYcfEQImy1KZ0Xe3e++KT7DipEybCz9kJn10s6Eg/IT
cA7xiVXh7jwcn6AgUBJBeetA8awGvMIAWz4hcnOscbo6EiPdFSCQZaIWeRvdLFT6EB5w+c89xaNO
bXVB82IGpKL6rO+Gldt0G/vhIKdXW0HmL5nyjZbv1/BrU8Mvm5eDLmqj1ALr+UT6NrF/ouKPn9+l
o8/dXQGi9BLq5o4YKrmwmaLDiDA7Bd4s+QfNh0JmoZVeU0IzpV6fos169u7rP9Fp9YjhxuakhN6/
pulLQ1/MO6DFD7Ldn3m9jm7mKrcArS3xghTtw394Q6ha1o60FovIoY7zlsWP47ypzqkruxXcI8mO
UBJCBIwCJfo9DiI91zS+3ntgDUxod5WU/1TCIHMO+xiq1at8hCoP5zwXEs5NF/3sgtSdu6BT+ZlM
nquNy4oYT4I1v/NnyI/X0q2JKErIF5v44G2y7U/nyTfZarDlaeEZ5Xv3ynDqh58xwGHfD0uYCCEs
jgCKos4k9LxDRekZOCyGdHb023uYsC4EnlSxLKvGy2CyvrjJISFs3+VJdENkiJTE1WmxigXPAy21
y9tQS0z53wGCxvmo5GzSpXKJh2t0E3WRuvgCs6CLwarSZuCvJBu8+g8pBTc8RRsTo+Ka0y7lb+9G
4Pw67m5MZ4bXiLy2aJbhVGVk/tuKTGMnLYofEHIfK3IIqpwoSl0JvHFfBl7Tk/i++Ywp61oxe08I
KMSF7BxtqyYqWlEYBnA9Gdj3ssarVYg+4bXpvtDT5u6LEnlwZoE3Uu6d4pP/04pLPdCI4oqluSYJ
9di7CvczR/aXhhaX0e0YhuEF6KZ8RrAP7GdiTNk5kKKcEQqIrF0t0E6OthWmeUTteNWn2r9Hy7n2
GyTBCxKsufWCwdc2JtdQ/6Qb2I3ZAFbmsaWVSoTbcPKePds7pDAJcSLAAxbmjhAmt282WVskhD0S
QpNqpwrGsedq6ZCIq78i+vbuuFN9QeC5ctwpLIBDkjcc9lMtRHT04ilP3Kuzfq7SaHoTrVDyrkdC
UNRTwGsNOQnIXhfeCjvDTeX0gSBV+TiTHMLoc+Ax1et+gSPXswEVPMkSS8NW0YRRtTTz+r7YuzFn
o3rt/opHjTxhfj+uuYgHOehdsW1FSlepDWvVfN5q0zjPsSPOPLE10EM7WdzxHle5HT4KU3psb+F1
tTrDtovTz6JHC7p2E1CwRbIx6IlR5UWPEQcuHvltYHtpRnj6PpVvuitgrSdSHg0bvO8bDxaCKU54
r5mq6g5KrQbBViZJgbc420qukMxxjhxGRdHsLt8NjabAXCsumh0A135HLjhlDFyDAmS3dlkDx8Mg
O7q0xm5/C4HCCIZJ0B5LW4asrBNg+H1VGviqhZQRXJwk1i/dvToF60NBHzYEkZ6RR9pNY1+6pdQt
V9m4NXVIReicZUqZ2VFWNX7ZyXKnNSZ06FIZ1mADxZyXfMbpQ4+Bj3CyUytQPm49lJtY/VAwF9Rq
+PSFA3bSeVjmf28tV5giirIx6fcROH+3K42TpUA+AEarxcP6F7qonAPxH7Sc1TOUBWV67ITdrLB9
nLgI4XbtzhImg7JorhitKoEMNZHxBa6cUtCS/2JWSlBITUmPKLdtqjfxXMT6RYgqdXWK6OvsIJ24
WHLqyAq4SlfM3BnzrKjhiZIZSl6rdCJYQkJVtjUDEDu4/DMwlaSXwo+w1zMF4nvQCkHxqwZIangH
cf+Qx0FsD2KM/X9mftmElaoKZbiVEyB+mwBpjxuVTanbBF9FDQdybpY5dQB0bq/Zr4e6WZ2lQe/N
7Y+IIf0cZm4hQHNrrGh1rp018h39XfnMUCpty3Ns5PWymFNaNK3YHc1tLOpkOpiEW09l56NX50w8
kvzWcEyOPG1QHmU0Z4vyI3KeAiBSdhcsP0JzGjNT2yVoZjDGBF8eDMEEEk2kXeqgrlXHvpYpygcQ
uOcbqZ1ObFwd+/x1GWVLQComFVYUzTdtC5qqM9TWJuFG6I4I0BeCtlbPjcpMAYHRQ+5P8X52wM7m
nawwDmCZ8SAB0woqLBCXSIPxBG1M0XOsVxm/KsAMKBVRHvzfBUVg8H046ouIHk9DCLyl0NbPcGfi
Xrxo8KYh+dNGE727wmgnG90rvBAJtqImEQSEl93RYNDt7VmCmKAYFidC4JPtaY2ljft3UKiCFuaI
jSeCHSG6SfYeLOueRckP2I44+mQ7KegR0M0UkRLqVT6Wgi71Thjo/q4LeeeH68tPd8RxhyL+Pr74
jK+j61boMcSbN/QyDKr0wU5/rEud2OXXXaKC3jGOW+jOcqUXwdaUUzRI7yxA8vb/yrDhYV/M96yV
iTOj0zJu7OxJD4u9e4V1YaJ3QsSOTJsxbtwz7QYikyiw0It+ZTfIzMzMRlJAUgOk9B7/A6Sk3B+g
bPyk3nlu/CK2lQZ7nQTqJtRAnY0zrCJFI35SseYXgkAP1VRZvcHrakgugwdz9eZEbtyfvQptRBBA
qQ4hoG38awwcMlnMMltU7fCimmIKYY84IZY5hc18cbTuNMBV0vK/0mpWEJ+XpvNQQt0Su7bD9gBI
9If+d5AJUHKPknouensTJcc/LT3YZFPsgqcqiveK7k8rwLi5PulaD1yFPZm5ylcs9wI3fgG//stF
mJM53TXzd+3tEF1TdP1qseGv8cXxyItWZ/KLgDNa9vBvD18MxZnqvJM6LM21Av9SEgtyWMeh1T9x
NHSUORGg6TaH7NjYQR3e/IcDQUa327cH+WbEyDaWyO8+6vJcYqZxhyVii87i2Cth4kXuAlm8EQ1Y
31xCCMqMNkhG7t9F1vcDMvEWrvfDCS7VblukXE8uko3170GeEvbddaQUGE/0g2Cduldx0n2WegYf
GTe1w5PbCyS+X12gnvBc/KVrcz4qPCE7eylSLsGsDdHfBfw8G0Q1TNOHHewpcoXXJ3W0A+nG0fam
7eG/qSyIZ5GwEHj2P6fPwWbyM8a6fsDHPXJiZsnMVpy1QbfR88Tablm8ieBY8EB76FfRClkcrpM+
To6NSD1hfgHvRRi5mvNCxYjoaMD2PcbmxjLDLTHtz9kM8daQ0x6FiRuKweT6NvcZ/XOlyFuVPIXt
GGERV5CpDHVT8FoxfNVYZfH5UGVx9fQ3RNcAinuJAQNKIz29OxZijzOIasBHv6QJFQzAWyJYupgi
U22iSjD0/IkWUeoAFF/NRewccjskiWVv9tJXSzuK/tjwzXNXfO7bRqJlHTMC4sEZAm724sHpS2EQ
+/Jyr9XALCm8Q4/2rdZl0NKMO+tapIhyfWnV+NHEqnRml0lEirLCND9DUElP6/GqxAMJbmtkLzql
xNb5aNRy27K9uLY9HbcjWQArPMN6ks5avfHtd/1M2rwPllNnTAeFZw5aZwOmwsaIp+PpTqulP3Bn
K7mrF8x8vf2WbFkMinxMnRSJvc3jUDsUrUzL/4zKa38xSRgfqrdvpqTZLs7P9Wy0qceTreQbFqup
xAwnyPuXqATNq8w+Z8hy55js/xjao9jlksdpKk/ks5+QJYw8ekroGFLdBf/6KT9hT08cRuSw2gmb
a+W9z6K5Cm9lhWrrPvKK4SegEusIrdmVnEjycZkP9leHRCGEuGN4hOPJB78WBTFCGTtu7mdjVYsg
wgM/riC9v0apBzi+TJoAAG6jf6Xr+446pj1u34mnreskYnHdpiVpKbpH4EyUN1Ai0oFxrrvc41ql
TsVfm5eYotGow3RJ7Dj8U1AgrweStIM4V6z7tsns32VzaiWMAOSHX0fj1XXIy8DiHGYN3t9WileO
j+0WCcUqGwyN7JC9f7u649istLPP7ax0DzDbuPnTUxdJeyrlZDnHrDOpAuq8KU2SzCmdc+bP0WO6
cqQrUYhELqkKipkkVFdjzwAeSukILBoSFEi6VaxqZkCS95agk/wWBMXd8w3gWnLb84jJ169bcFF7
xJuIhExeeTXyweejH4hkwPddYd2gVJpd2/2tfBbqaPaixnkRDFOXm7ZOHYkY29slWT4KGAOJAtco
waLsG6e2kGuTHVQNXgco4OzPUiL8pYxLjYVst6o8CWou2IQIBAqQqHY+CVc4eUtZZDLNA736rwCO
+ukag+v+Yu9eRPxLZr0t/tp+1q5K0HxubYt3lMAohiyuaRKlJ8URhLtsM0BqqsMYDtGGgyxBD32E
dSpOpCRkx7M5m3dcRD3NEVhgWpL1a314mhWnYQZ+neNInw20iD2jBxDH7bPuDH7wyRve6XpkTE9n
qw2zu8QrFJ93gGTGSEMG5FcaS/VJXjZrPkX+/N6ohzkmvDm3RTa/Cefy4SCdJdk3hp/UG5Wr65OO
mHhUyFEt9Tb3I+u8k/CYm4voAmcs21zbiIs3istIRyNptRaA6Kf9Uj1KSJnJj3YffoxZHVFsxRwe
fxw+vugufB1C/2ew4K4ttrfcRNWInRyJf3Hoo3nuaRGZ2NIO1xRT4/QmT8RGjQDPkbCcdtx6Syvr
Wgg5CJEpWMt0mrLBdr6X/+I/0ytHRu+jYAKI8hmvblY8ZvL7/cNLj25qThgTzbkvD5AzjLeWBsOy
Me4h3hDen/dNSdfcuCXyakZw34AjtowcoYkhAE471KGtS3gwN/LXV0f453+hhUpInsD+9S8d9I66
TuvBEczPXasxD3n2ku76p6igbzjeXGVWwdY5e+SjahaKqfqrpEMo4CMcMscbxhfoQO1RnIYG4LiI
1Mj4pJ30lFYF3OrDV04hAoXltAlYc2Rk0BGtY8ZN1WNqYKo1Fd0DB2KhJHoHrAYRdjE5DQdvRNGL
su8G7VTMfSJPukT26MaQl6LeHLnY7Y0AVrxruxMmuJUYGlBLXwOI5rnuaPsWsNc1eJ3WV/oFOjnw
wM/Lf1xkIgAYHZ6DJwQ4TVUdGKNLL8AOjkGk+Wck1zhD0XL862NoNERZghRQZv+WXV+r3iTVwq82
XsnFn+4rcbTQWZlGjrt3DZwfrYa3Th/Gc1CtRu0MqOY6kCujCfR+DulB80RanOMxFkgqHYpvCIHn
hHOtjZUBwcGHE9Wt7yRTCI+9cAwsbP7uSlJUILl0t641pqIY1QkZx3TqBuaA6BnVcKCJw33d5Ebp
S8x+xwtZiProPLGgAKSScuoHrS/C4A8fjqiOFwSGCwGJp7YEAiD1w+bEe92sHcjHO6gwNuWoDw2u
c9+2PTIGjhPOERpa7eLxnkNLjAjbhmKvyc6RnuW0Nj08vcw8dsJXDqrk0tiQIMM+j9IXQ6IJ46iu
nZdLqJVWBLLJB2oIkvNI/xXdvHZx7bj39qtzsxfG4CyKAuX1d4jGp1mXzlY7np9Bc23zCKEhd0t7
zvkiSlLS9qzVmXjUy6li7XTHVvakWiDvAJiZRrNIfx3oemQpsi8U6wW/YVjGvkqwAA5YrLZVSPDh
bV65QZwSFV4Hn1diDMefTFmZnfQqYwHV5yr6iOyeruUawMPhq5dQklYzNQbPTexaA3tgo2V0LLSD
/hBmZ2olMTVdVPpogDma0EdYdUUvEnnTaRcKhmHKZjoHBQ8s9UrJoLVj9f5zZc+TOttklDblY1pe
NQvgQoQsIvn04JAZFqihVQOLI+Wlxqyz2cuug3ck31a9Z7Ujbl26L9ttGUUrR1OLaQNitFv1qbTl
hWSIyx6emp3nKC+x8DtNEzNDfs44q2/BntlgtcPNuUt3DFx0Mcf/T9YsGoz2PKWnAliQKtZqBCc3
D+jaMXcpgXdOCfRG0Ni4mvvamI5FxYigYZwUAhjVtXq8ZW8XTmR9fTe2AREJ4sAyeOGQJy+Leos4
Icm/qUiovQq4JRnvRyo58hB0v/2u9rRp8xT9aEqkEuIBjymQwJ6uhcWAbhpgtavMQRgOY+K9dWdl
8MmElOvppPbVQNzD/0+hHEUsV9QmsQE7vU8kEJIEgy3U1cD+sIKREhERJWI/4xmGBTbi06K7aYsG
7kzyQfFeUm4RR5Ub7YmsNJ1Va6+INV+xCAX3HZBh4Ct8GVPfee5CsqT1yvuufiaC/QtQuKM+M+Pc
EGLexRWm6QIVG7LVdFsxinWCj89EW3DxdUtWTx09liuGLb0Rj5BUJjMU6T8Elu2tQy9LB9OlSFA1
Ma4FIpQSrAoWU29RX/iu+yKacdTmMaN9WZtmdO3Jt7IZ9qrvGPhbo8e2mjw6vsdFnHGR8qhncUW3
KfxZhRk8MWdizo273mM3gW2QW9IGDh6VC90XIpkKEwARNUO5p1gc8F+FJKmv9Zw/dyEGa4gdWIBn
D/LhGLH8NoF0XQkYjDL6JOApmduksDkA45cxSwIQ8eb2dABbda4ISg4/qAttc15P8ij0u9nq9DXB
sJ7ZdttQYX+BL1zp1iAYQ1CApcS7tyo9LRUKoKUM3l4DycVnoXJz7SQmS1epzsbfpT+bq3XXNVUc
88v26CUJC8wur39mSWgAJb3gs7RPz/SdVyuje1WvcIKo1tNZqbhOQNvNIwby049DzDIcy6ZiT0cN
I3DcQHJVHXTOeRjIb7dNX+0CearEstlHxlR8TchRzQ/6JBE5wjDwVXTMLLo+QlW+YcAZZYR8hj39
GepR3vgqnW6IjIPsYeHmJMHRa9m7QAyxJ5eOV0OyhJbPIhO2llnVEP397u92dVL8VRUeoObAGDIf
iEWhnfLfVk/dEs2Wpq72mIWMPyWm8+QuT6B+OF3Qwz3yNTjokVfqUxsoKarHWwTIgbGf/fz2fl1/
mP2V37OQNJktlKUu1Bv5kEo83NgSM5+N3170REj+3S/C1Yq7NqPf8RHTRoGpzT/Msq+f655Uy7v7
AXJZWkLiVgHGZuL2hPHXPHKavT8U1LneEqdPAUgkIEOa9HeywK1AKiPr0A6EhGr8QxFVZxDYx9zO
IaK/+DjVNFMbVNbMuCi+ge9Qaye7+XpQ0KoqpKizIjVgIiv3/dv6vkto4nyZjiGFnx3yzaorcvul
g11gQirPgguhY+nVWXKi3/nlE4/gXLRoe2YoLlT9vJ8c1G7G3KNeEr7UJj9gOuFar/UwWytw1hnx
+LCZ0qg+C3aXcwbULuduN0QhY66GZfCiYza5OwYqITDk3+4vl+5pFjXtGwjHt1pSTwNHxHdMU2MI
57pYJAossFtR8linQUjYcbi9c4YTEi8WMiCYWvH3ACut5V2uDwn1iXfFWpRhUZ+w0hoF5UVdBTj+
dPH4R1Yd+HjCEfrdDNRzQGgkXv/RieyzFb25T0/pQ9RKNy7hDHVnYfWpm+cVGWwnUF+5KiUXw7DB
AI+se+hLMgc2r9p4o9Gt32RaL52d9yizd3k1iwGNAAYlTWXmqjQfGmDpPm831Eae2Y38bvfLIY0N
xw35Zf2t1NcTBaXf3cokFblUnGQ25+JKne6BsfuRDI55lreEo6HZem7Pddy30Mrhss+ep0L4j5rf
Evdt5thQzAigRIiuMI+/2OWd9WNwe+qD3Dl0LK4+rBtSThfMklEIVyE4IkU4y+eV1eT/Ive0LAEd
Jz+QoFdgEdKOHLEmbvHj/O6jZT63lL3Fu1lni25tJkK/EZv0UDPwZ+RAGLUDTv3u70BKLEUddzpZ
1H698QaDkmcd6UPxbadfaM5e/vAODaFG9ArpTbkI4BIzeodqAEPm4weqQ0umZKxwvJkcvAPgMYZD
zcSDco0fd+niMd1IJoEj3XhLqY9q+LttSi1l8V01r9RAnSpGUM2cyUn7dtGmuaXCtssWOj3gqavf
ZwmW4B/J63XkqNc0TSdfRzS4aTYNKJc86dIHTrE+VW+wTZtcnXg6E03oiAXo35S+mkUv4au9IG+d
9Eyw8NBZlJLh3hUrnIyFucRoHza+5mNDPR0tHlUdNDnKTHjNOU/LkQ+5gQrSv5nGwPG+ZfIvCm6Q
tafd7joAzKBR9ICy+flBYAjI0+irPCdZB45iyG+Y8QGM2lGBAocfZjG5WEhid88rYPl77N2ycdQT
IpQxqISwEecOQhGj5FjyvcynMttxkFGy2yC2EnsUHKTlvL9UgIo9W3yhnfchcXw8yJff1wvVHfU6
LS98g2OpZdFei0cAPLBfuWsnjuSDBsSPv6w/Ti1+Qi4pd2aPA/KwBaibjU7gOOUJ91NZCMc164y6
w31CR9h5D5cPDHDSOq3cQ439NN6X3kjcqyMVnWqn3rgXdla0i34qy1bcO0qE0+AHmhCnlIrl5AgE
Vk0zgRzNiG3SBvGwa/9LTwVvYfIuWccqSLm91JtjDuPGTItcaZe6qONw9eaaGDBTvsM924sQthr8
937zQt5otX4CzI1emvNFqPieo83esMI8uNXRKtqx7oEdW7/zZEC8rbjzaYSIy4Hleg6mr88UBviB
rcTervVxDkCbd5eY3JnYOlmy3YzjFyZl0uvlE1vAj5XaGvAJCQuqMK8dO5fdfsXliIYivsXcX9w/
5RNwhhaq6LeXn8QUV9XCe9BQvOGplNMlH6gkNQ/S/N3PMG/I0koW5MbBXcojw3em5unosu/wMTG6
qqrbF2EbZmR6cefic7aL1VYHECU6CtykPHPNczmqnPaSjzIeaU4z5T3EfimKzgkb6/3Yj6qr9D8Q
J4Zx3nl65zqePTiDuM0TSHQlmk77NCoocGmzojdejdGcCOyBBTcqsBLm2Fuhyyx7xbdYC48BzNJf
qukXr+v6FHrMKwDZQaF8wZmxk6VyjODh2cQJwLq19Ilymz3fRPO8mf/KJqHjGR5TJmZ9fa9Qdlh1
Mg6Ax87FGwmlsugQKULsmZ0+FPavUwVGpP0+dw0xSrM9w7s1t6nK/71J1ngV8LlLT+RuuzXw0at5
WN+Ya2ZEkN3EYxi7ThtD6wvgIYaYL4GQ6+LxQtQOGFjoiOIuv9LmKwtmC8o3djNrYYQhs7cTs7tO
IQ3DjCLgfVDtViLx9+1hlg09ku+sXMVIwI+0yt+epf+mT1tAqEYd88lCdk/3d9CJjm3TbxG2w9MF
M4YmpxdsaMETazRSvH7VC0hxO+0+PGYYUPHwnUpJ7CfuTULJW4kDPKrB1cbjCYDcptZRd1RR+CdR
Bg41hAzM6BW+eq2w6J8bBDDjkW44RfuikqF6yzsc/AdisWM2SCTu7/gVHvSLNu79HDGGqM6SA/nh
rOrMNIcs7XBOCJLrFvAhPxt7F/3l4209fZH/uNy3jE0j/e01VNFKKG62F8bbqaqbVFOUc/C4TosK
BHieM6cd17Rt4wTWG02CneWHOvswUWHTjq9P1V+GfI6r57GbAzOO59FEwMi2a6pVexKSZWRQk0hA
jPww3Sr90ElFa9DsVghZrtKmWE0m+T0vd2YvTsEMK95w1LWn9DV8QSdMHQJjxQbv//8EFDCopLOB
X/dOetNTzKjDd7bO2v7AMgU62od674mp4d10bzKP1wrbL3mm23o1+3G4sxPAduP09B4JFE+rFdhe
gAySW0TkqB0rQzTEaSQFNRlImNd7gvph/Kq3HS9z1at20KUv2AXpRq448dOXnI56SFVr7C8YVk7b
3J+tc8Ldb9x0Nva/YybUDwXX0RmLt7WTb8fT+kaheGtiXI4BzAYjxFP8skXlZBGkT69UUn/gTwSh
HaDwYjs6R3Jb6o+KrdyPxxTKSYdLIhCFunjogWiBBgcqwf3bqbSNwruO8xnTA6WbBaFinzSnmXlT
dWdlwXipJW6DpG16AbNwwRbW6Sdg5rAREM/sph8NUvj7MnpizA/vjeKBilC2E2Mkdn5UZ1diuBW1
TYJbTBASWiXFecOB8bEkD/vV+m3tFEwpfucuKAOt/VGK6UrTr67ymVnf4kcPBEtCnbAVUlXyd4a7
qVImVJW8k3KwYESlRUVreCsl0nJP/se7lmFlyDi4O/VAJ8mpvsmRe1nJOlyMRWCc11+ecYH5goW4
RbTQUQU093bi2AS6HTcdPA7ZVFQvWBQ8Av4zka2jePfUKnMHcYN8xuZVl0lysQZR/uTUDMjVLHQR
3SZWPFGSHYHzuhQ+vDZdXmeiRT8BNc4WXKQYLLYKDctbDauKioWX19HRPNkD4G6K9TLBEZRnDIvv
pNOEIYpAokqnt0llD9YWNu4wyVLbMtxAbZh35Fxm++JC9K9y19tds2GZ0ISoxX/lrTTBpVM+yxaj
2T+j1VC1pggQi/2WDK23qkzr7u43+D5CRszHyRvj2zzRn4YJySsf7n5WVZoHd9xX6ST7m38aosM1
B67Z4LXPs44vF2TDfEPqYMIpLe3CDAjj0qoXOwlWKlPCxeyfPRK+5vNkfYx2zWpz7B+KiBr0oW/T
u0jLKcYwmK67HmgKUatGHHT54CjpovSn3Dfls329mabWWU0FvikbX6hZuZfYsW6Q3qAixkWxgwAG
yeT9IfsEXpt7wQZ7/7e0U30rE5SChhOwjj/489LXnSU24VT8vbQa+x80c22FOQ4vCphn4hcdfK+U
NyFt7wazpUCZB0Awwl48o7LqDRX8jLuDgZivz6L7r8mwdzapUObiTQgOXuWYTmOkPAtKuN4yuMFo
kf0RttT6NCldhm6E65hM6l8pDN3jJdT0sCbQGpidojCTz6YZRJKX0wEVsZLN7hTEAeTtId442iDl
hO8g++ioX7vX+THLF5r7+zVnodXElz9rvmxNR/G2m8jzq/maA7m00Zz9SQmfEzFtopR73E8RE+pr
hYTCX1zflhfBtJArFpuE0UDsmtm2AsIFLtSh/21X7EVR6XvmHIEMh1YmlNjMa5wKIWMCK2nREiQa
8sgPhm+EWUtI0/wHhMVMkDe4Pe51F6qmdqMwxeC4CHa8xa8Pq6Z3Wsb72wbtEuvu4jAtiIxebOY3
lBNTGDOTqScUOmaqGUtSEwd3+PquDa7OKtojpZUiMzvrcXrFO2snTHQmS5HhzOQd3qa7tNm5CPRk
qlXYbagRlbszD+GlZyqt2GQyPsUolxFazugGEuA3RE4LmMTfy1/TT1z1x7fYdqZ3+Dloq2cgsW1n
9o2iBIsZ1oiyT8HudOtxwm/925qOGG/iGIfpRu1AwENzXC5+SxAVSM6XFSZg2aixJqShh1q3AAbS
W2zW8x9VGgxhUtmtPGIVMNn+ZwlaLGY9vACiO3rSZugGMilFhZDZsSUBbs7PSR41hol0Gg6C7BxT
EClerxHHehTi510iNOGhyTWavagojMmrqQ6j2dnDuMxikzvKUwvM+88FuOJZoSAP7SwfsfHetSg7
gYtYpxS0Tkh4qqmobD4nnrt5Ih6eW4ynpmFeDB+ykoncBXNyqWaieMrARP8TRN4/Djvj4rxdp4fm
wLK5FwLcGzq7Z0P/vsD1it7l99Sj6bP/ZIOcwcf3CdC5VPBJ6KnD3F9LJDnUXLcsJYKdHu+rZMQh
zp16odZyHHD3o4hq8D6e4UrHJVb34Y3qO+v5SzDHHrIJZlk9yIYsM1O8hoFJ6GHfFkts80LSds8E
OWNlABxz1YvQHBwSz98E7C7tvxLyauUXMKsy4jWov7KQ+UXvTeIk90lpBUJf/uuJyBpFwwQ4JhjX
CBzMOavE1bszN4sRMJi34WS7jayfUHQwkr2FmTE0lv4dWdjOphlTWdXT3Kgqs8tT+Qwv4cOzu9E2
y3D0PVJPxz+hd1smW+xw4MEfvNWzG0jJmtAs0yBGN58/z64ERGDBhb4mnGCRVj1UFfMr/sdOhkP7
PSCGsegSs5/5dLBe5KZfFKaE/jyC6ZeJP18ehN6hnR3j1jdKEsnsFB8Y7BJ1pWwMp9muMj0GRSbi
g/XkcFZ4KadupdxLoW/JwzmToVfrAU/Yl2pqlyPVmeucRIzbzLzpfbyHgcKMhuwf6o4BANYth5no
YB3uOMZef9Vdf3YF8FNKgu5Yq8ZzQV4py+Aepiq4yrYPGaeP4iPKich1I16GaPifS8m117gi61u3
SfisbEZmTz5c2IbdF2oILv1hn3cPorebZ1CGUWOgIrtzPveQfN3MZXm1z8JRHv67l6ZZ1LQzBtgd
H5fDpB6L+xMbhoyIhJmKPYNjM1G8XalEA2XiPfg714WjgpAQ2KO8AYmBAd6UUUOHIDqk88UpljC8
rjimDq2asEQkgkdiQcTFSCgFTfHiChQpWp+5igGFJ1RcVMk+leNAdtcr/MuvxPltaFvNXnhcAJBY
GSganaE+CWQBhFaw6tpngjxt4aruIbrZ1zhXj3smI4A4lBcnmp7xRGB81rRasWlHyzQFrcoGndIq
/bUCeCYzj4uhEMi8K00pRDVz0zS04oR2YF7YJJqfjzBBfehtbgME3U0uBHIp+QXrQD5WqxcVYOr6
P2xziU96GUYR1yITuwm9NPN2KQS9Jfutm8oucbVvb833PVuky6VNcnj6aYLv2e8bFltVMQ03AifF
iEx8eqXLD4wwMOX64FcUh78S3SB0qVEZjFNXvwdbt+Cu1WsT+8Tym2w3BFgmTadKQRRXR9WdU0f1
G9HEdTf6b3Mprfs2yC4BmDirl5GTm/tnRJ4hXHiNsZ+EuVPSCNM2DKkh6IQE3xbakJFI5ZTSDd3I
LqAQDguJdXX2Hw4u0Iiq3vwIaR+vwErohjoQgSp/Gi7Oy+yZH4JcHsZwag64N8+WZe8bxN98np1g
PF5tAkBKz1dRq7nXIJQUFM7iVsUuJC3AkfAnogbiJ5WsvGL9RBtlT7n9euitvqux0d6k0khnIf5L
SSu+oqQM5rz2jmT8/FR0HbC6UeVnK6I2JJJTMA3Zi51/fW4VA2kOFXVQZu7mdrAds4Sr/Myjxd5J
nOc/uilPB8EloQRZ86tW9Z3coYWc74U/UhsHod8Nt8Pz3NtXhANXkeyVtXwmk8CE2iXK+nGbWQXX
5/GJMxUuvTCqW07j+pRLkz50KW2wYsuKtEPkvtdEkVKh0nUZ7tcgPLX6YEGZI8xr3f63RQUriGmx
00tKOalOVAkkhtarUvZmLHPyVdMqJAAqJ6vI9plg0iU1GI1LcQDAGfS0jIUQdMu12GVbsWsfse30
vKCIHM1KJR+sF8zWR+4RcywXisz1hKaBXnrwbd/snxVuVQiWxhfIrpkwKZb1JZAPtf54fv87EbGc
Hl3zE2ZWh/Yddxo9pSyeHuIYFPwgwHIJ/D7OISoyd5ZE/D4SDdkzs/mQSn9masqCCdcJPb9ndNcG
1Y+ZfIiZWsV2E7vtwswEp4X6uA2AdsxKaWFrJ+Jm7wbjUw4c8o8CPdrhLRzOcecgPKfp54rkxh+Z
Ro0+U8Bw56uGi4FLSOiyvgKLav962HsZeU5WC3YdQ69IblPHl1v03TSg24DbzfFmtB9KuSxKq4nk
PaYtafUIqv8E0tpR83bbzA0v9dcu7RW+EHHcbffQQbbpKlNFjFxi6QAogkcRdKGg1e9RlhD5GmF5
yJk6Xl5BeVIKn5CY7lgeFgxGb9Pgx09u46aNErWKOW7ISejpAtyHGH7f9Ot4XBrJ6duDtYrU83Ni
tuLx+x4bgUQ4qpT2aBiN70QjFrB2RirSDCNio6Po07ce/oX5hNbchv3XIlG8e/r7q1cjTT1qMXDL
+cPURD8C+RgNVMtorY1l1ozPg0mWgpXOBvQFtDg3noM0YkPbPciOiwVS4YFklouu6sX1s2mV/zoP
FK6FF5NPVGc1Er6q9IhnEb7t5mFuOkPKIHKTz+glX9I1cGjI4BEdWSP73EopyzJiYmQqVFuyP5IP
7hIFTbBSZUBQe2RZig1qtdEEkyJTbaS0GoOlHzTeH0XlEfhM2901Q+qappSmgZptKr5/iq+9OvIz
1x7Y7KHEM2BmwSH3hRJKKbBRyXOmC7LIlDsFRyM03BSXCZqImbAdITgF4rF2htnhgu70v0WDQ1Y6
OcjG82Fe9vfCvcq7FjTneRHxufnDxL3JYv75CkhuKVcK041G5vYGTSkVWWjb0wHGFomLf6uhOvAD
hOLXVwSx0oytn4RBa0vOIGxmZ4q1BrhwXJj3fRZBnJc5LiFDKE980mQ0zwaFKthKpvfNMAAGSORb
HB1IwA2PRszgztIx6DwTUAp+YRS7MXRZCcmChSq/kJW6TD4uWzgp1pUefRM5f2ZaJu7bQRX9wqq4
H6bNDHTpju/Lkub3XYb3G8VbBM0QDrZt7BLW3/qr6DzuymgJ9cZZqh91E9hzi79Mym0CvoVEdgRX
RZ142zVYaSnCWP3PXrBEYgWMpmsU2yKqswL65v5FzZhyZXwCMhM3WE6/GKOhfTCFWxVt+ZJ1dQG2
HY3HPPmGOSN+p8vaCMbTHgKRK/IWJ8KoAT1IjumqYVbSoY0vAcm7iFusmKdpLUWauAymv2gXzNvt
2KJu4F9UJTdxl/9VLe0bdOkEkfFSoe+pSSmKFebezCo2/rQi8QNv6gAGP2MmP/iiBXfxI1KkmfpS
C5MjZ3/Wqdx0HPw2t32rdhL3k6vAnOBWOxWgZlM7KUyUAW53xI62GFW1DBjgBN8MtbymvR0WTA4y
3YMtus87SMEwGfPLJvCAAwL/AmqAdYmF0w5oBzyFz90AZVn8eNewKbfDd440nNa0Ef/qsjkbq4rp
H8+Du+7R7pZGYC6QpYrHZzRTrIkaMCxx2lErWTTMcoP9ryFokYnTE6khe2cZ2NYz5uiz6a7mbtqa
rad3vhfR43WFIYjTwDcVr9gC31QVtFCQt4Mw5iEofDmILQTgqzzGyZekxYM+LBYVy2yrQ4+0Lcw0
R7W2pZcp4Naak/VyMFodFlkLa6uJTNWfXhsH0rRZbYkIgbZpHANv2R77QAP5wHucpHMjrlzgOZMS
QpTMG1wvO/8cnJjqWH15Wcqaaxt78HlLzykN2UasW314oydIIGikqoL5bAeqKbMozJFYKAe3JAGv
sEWQF7sXADcCynwFu8bZ+1sCJaJb7Bw1gXhyIdoKUVzmiAr/eykOloSPnp9wtvmt4pj1saXfb182
HoS9gnP3ha4smlvlTcntBAKwns22OUZ2eVbNYo0fxr4mN5GmQ+LeBRFUMPCMyr3dlzv3MqeaAonc
ux2Zd9PtaSG9KvsPVkiWXdaMmqi2UzCq304Cjcz0u1aK4d6BGgnpyY+xLaDZeqMsOoFstarOEUT5
8YlzZFqZ7hAeQjPXsMeuDGPc4EeXPGYvwZEZ3FehwgdvqI3GbkXUycOqvclxfQ/9uWRJM67UJ5+D
A6VRFOuH4DD7PgJGbBDt1m/qNdTwTM961mYTfH65lTNc/50uUBsIWLYNrzOLRo85QiGP9l3bUxYS
3kIU4ujD3XvCj5ppy6PygLzwe9oU+1HMq12ORkckQwevCJN+n9HSH699iqvNX1n1CtrUkWhto+bK
5bnTlOelB9LJMRsI6/jX/Ao3Ae73B6/WveBpDty7AfFhBSluaApOrFzptfub+wkXcgZL8bDU1PTG
/63tFbeHSktDfKkVdvcTNOPtQwIEYmaLlONTBxOoRwEFnsZ2yfl+hHDfdvUOGHkweKkAOTiT2LHO
nbFuTrf3ROiij6I/E0bFW0pJ1MU5wIOWG5O2CjZ312qDwuKYkdp8qpQhHz66bKfW9nbHm8G91Dlv
83ibiK6UGTYC1h4k8QTWe6F5TNyHxictGeZZiRFi12cuUaCpyIN/pJ5TCWGy+TrMeVoR9/Bm8794
NNhLC/hgbf+aEvgoWvxnbzM38zsXHX5N8DNzGrByII0SgYsIXuAoYbosj1kO9g7aBesQnvSnAXS1
ZVE8vt09LhEKlYjKVQsYp6SV27UbMCGEocry5yqPLuchbXhXsk0u3DOzBVlHwJ6bWtplFvoLvQ7G
gYMoOMpBOFN24dDvT1tSjBtS7W62dw9eet8jy7qWqtBzqKWwZ7H9vtpoiQuuaN+LxcOAvgGY2/EC
nf12xHqRsVLcU9uuhGKMnaaiwopPHrwP8FAxMOlPEoE5Xclk1Qius2RcMSsncLDJKPp77XA1XEj/
qbNHsXoSvwOfTWWpiqqtdaKACF4jvU1dzffB876ZHJ3eMycD/LF+fovNHXlyJaOhjiRNM79sZ2uw
NJyVFdg9JLsh/uOTGHBd0HVisn0rQ/8OLl+ABMYJR2xRjOUgN82HCyhQKq4MqNkqE7jdpBGvROo+
U3ZbMrAI0L5y73yj8WM/u97wZB747s0YUtjnXDixwgzgviZEBtXfu4GeI1GUktb6y7ixqq+eftzP
SWGsSg64TilJ3MxYnZEl2okBm61+RPZgdUj3xFd6Lzh3rgx24CyuGRGxTf4cKOtDf8chW1JXvvU6
1YAnhKE10E/wmqc0IGBb4D+WcG+S4ikJGjFpzLYRrSebpNKb8eDzJublyyryHdj5VPnToKdjJqfq
KbAgVkodVZzmwg0gJpUsolMIZFlbcsGtWsEbbUg5c5oI8p4GBFCl13OY5S2L+AYWcpv6AXPq14Qt
9hy+joQukOCTc/rz83iBz+yh7m6pTEPv1/khURvpwpIVQ3m21hOHkIrk70gFPs6VVB/7drqeC7VJ
F8xZKllIr8N/zF6GyZKacQ5H+yCSmRR24S16s/uNEhquDhiiGQ1dXTVFQrhZsCKdvTgFKrDrXV0A
EAJ1N2vH2GNdWhhCq2sKLbfDA0EQBWL2ouZh3X8GLNgnD+GlRrSCpbP1eFaLh5FZU6DPiOVaRlxY
n7njgolaGDGGanu3AWZAMe1sz64ZbcDfw/5PfVLndhx/LAwWbGL9phLPWQUVrAjkYC/1+klpo1xU
+u39p9HSm8i3iJzVCCPiGYA9G72cgYBeCHmsQbbcNbg9vaPikPAvMt/Kv45YRru1R3mN8+SmaeMZ
sS/2mvO0iaXhCWvBqK+MmBURwWjJy4UOjErlMH2jBH2jQp/E8DGtyxxUI2ZXuNbR4Vm3pcDXkHfV
Y6tcKhToDF2llCLx3r/OC5WqLQiFNqCfYbQ2oGz9je1af8lpXfqC78dKlV3RmCmdv6xYfk8/VFM/
b8X9w/pEhPFk9o6M7KxbYaxYarqNNvdZp/A5+uL191JnxZZSJv4g0G6WVO6TqyNmYY31lzY/KfMI
z0WgI/gMjANKJOSk3zV9toFQrUNed97ei3VhfZtOaursU2zXEaGP3MJ+OlhKMdECn+KLxkt0zfwV
/918zkdgtjymFOlabxkILgbZJZvoyed9IwYyYkjgU5Hdi5MyTCUXist6uQbUlNtQAwHAinz1vLpp
5xWk37Kj9ihYp47QE3HY6rRlSKfRj9+vp470eoMfZjN17DC4+U8M8RHaMFHDYOwORZe/uUBKjvWE
UqmZH3pbemqewNPGY8toVelOGzsnKkPgvCJwdfR/ecINF5xqbG6Z7pTaHAuYuRrVIRrYxfoOhMWO
MLrDwb6RbxnWAsphP2JSFTYw++HGheSVNunock2HKRjubqbKmxJUCtFdMtx9zD9ASgH+D4HnGEna
MhN2nS7dfIgMu33JLKaowDNTRQohoNqY4/MT1fz5xB1kKSF6atAehgvTwul1Q5y2Cfah0wQFba0J
pdX9zVBWEJZpyUNuesHWEuuPcWtLzu8cifRhHHZ2TU71rhu3KyzBIbai/fNbfIMi1NkPA2ZScwkh
0QntRBne8wsUMrztRi3ev1B64zt/B05XPbtSUhMZqFS9bpOiTCrzgKyvda5QVmM6HC7OlOrKoL5B
JWGuqx7osWdPhvpCRE25t1ZOALbhd7o0vrxSp4YuMcTa7Th+ZH518fdVhIc9/gXAQuJSwLsj0Z1f
caeMH1OBLhsvQIsimKjJmDuyW1PMbMzo8bj3np+rQIjPHRJGaznWYgIgJ90WZ7MbnCr/9seduz8b
GleKgVezVpMsis1R3ioGg+qFpIU5GMgRwe3h8GP7wfuwW2Nq8oraUsWyQPOHpf4Tjka86o3MQfnQ
/4DNnBHmLmTtMTeM7NlMTzxIMK9dKPiIHWgm1/ZwUNjnkvRZVtYJIeo0HC8Tc0w0pPuIEmvBRFLM
osfjaYCgg5ZOvS/NiHwoKXbeBGb6HjvRGbdV5fxaVS+vBbxTEAcSD68kUV6H2s3cbOg318iWZGfI
+o3DX4lYTgHJ5Y9gDHTv78Tln6qdZszxYd3GV6ToHHdFD/2bTdirCYX+8qqvK1rsSeRipDoeML4F
f5nuerZ7JZfXjls0G+78LapCwLxOwFeDBtpHf+HAU2RGaKRGikyjBoX7dx33WmKlxuVQowpfQFWh
IzYY2OpAQHqnxssICexby9qvHm9uykCxh1Hm9pdZkBzbSOP8kMYshZGIGgsjsf4q0oYCcssdDt9V
XE8Uhopqx7ANN0w1LKhf1nBNXJs88AnByBTCcTAa77OETwdaSdveK7KvuBOT0bm4ZRDthw8ImY1W
aZzk9VLDPeRB1zvZdYuBhgi+/lc6gs/2ikaXaRxfDWFl59rHc3xSxIovVU8JDO19Cc4ztlMGhT68
cbMgahSCAGF0lSMWhs9dVsGMZAUNPT/w3dV64VyusY1r3xZqv/9bdHI4AuFL06K2VZI1Nb9k/g/A
nx/shlmEmzur51M3sRhPs54t8LZWrvl9P3ZV3flnbuJ0Z7N9QJaFl+xMAiR1OT4ntUYzy2JMEZME
MDSqnM78pouNsAiW05tHcw9Ebdiu2zG5iuWLrrXT6qFW7jdDBwJDH8vJed9H7XvDFBewTeCOng+k
cncNXGIIdP1anhPBO8a9MJ/RQ/C5fGJ81IAt9EmIInPbJvDZIg6qDEfgi6qX+wSgGS4enismxSTP
dUzLDxAjfsgi5At6Mbw0LUvbaH9MoI5KnMwFi0AiwCBE3pULnawgTWlCd2Jq5IwR+I9gQrEpWPmp
nYMC8a33c1u7DfA339ZjYR+K3S1rBzkiEHW33CvDdBJv5W0XdcYsGb07qgtJ9B7asIroiRQHGSIs
qg1p7Pia6zMzwoqmcPfo64PuHYkGj42AgBNi1AmCqSuMYRUr7RvWJrbRKYINZa0BBtDhWBSh4Vgk
gUghBIW8yAw4kqCLh67Me9jMck3iVbKTyc2eBkb7L2eiXuqg+Y/AKkoEOiwz6PPxxUuy3OQ72b49
NiLijmDjIFNc9Do5xv3ba+PNrwESn9VzzsO5av8PuwgiZDZIOUaJHxLl6HnLPeUidwET/QdSVd2+
AWeuoX8+OzxSPsdYYNZtX7+7KdinsrmjdEO/fdQZ2lAy3mJjD5d36bqyymNqp0+ZRjNHtWK65E23
GNTdEMLQOM0r1IDEM6BjMpYmfXb5H0r9AA7AH0yfbAElWfQ2fAgmuDUpZGI2VLYmHLacCnwhWNUk
eJ1wMOf74Z63bk2vNz4WcIPxBzUEsbnAYbGLo1gJHLc9bVDlSFsy28szuqkiM0cgIlFq/TEkZa3N
JftgshfoNqy0Bw94zHeIj9CdpDudMyN+1wRK27HqY/NptgfQlwaYFxH+l06fYxuXH1rgG8y7jRHo
fwNYmcwBSBQJQu5FjlleY72JpseRt6SWe3txqSdR6/lKB45wMZI7BxFkDohpK9WRE/09HQg9u7JO
ROcb1a7WikqEXVPfMhNAbHZLfENuNY1e6EfDqmgT+iKQI5wFMy6mgI79IGcAWgFLxq6s8OXNkD5O
YqiZVL7XoI1N1ySDhen7CT17BpflbGzmntSrSPbbzh/GfpvxGV+tVIixTny3fUlNLvJvJuIIgYUm
m+XLPtiXLqQnbNKE5AAEVDw7GKps93WHumEGHjTo+H/Kk0fcuTuyD8v7eTj89ZkQVMWgIg3ASR6v
mzxoyBnHUXS3BUm8PGjbM/Z2F+WxkMVRa9OI8ANkubbeWJVf0mf4hdGDflYminwGR56Bfgb/IxlA
4hf7QvMEJgXXfkjkPDohl29ClbQIOE2ze8McURF2B81RudIwGHndFbCwRyFiFSWLGJnqsA+Nwhz1
2WaUSmlTU+xeyIdQs2lH1SApsjzdQ+q/qce+5WvyMmW1yDG8WcRp2gGE7EJ7Ku9xUwhcoPkdOrkh
FylxXhcKLLN5rxiG5Lt3HU5zaRbmYCmcylPhX5tuTTyy/x7KZ/4+czyfqS6kmrF/ZiEbuJG0/uA0
jpNRwOoaHjJawczg1kwiRx9bZS9sed2HdnlwmxXcQ0fNCf+nnD1Lul0Efcnah4Z06MXRdtUfK0x5
SxL4sA6csYY9q3ziYX405Ger48OW8Cv/Zg+vYETKN6TnXrsZHCkt+vbz/+fkvBxbOLnpZ1fbK93z
tDqh7KW4eOxTSr1blm5iFiQtDK6JPntTilfjNKI97Z/2TEiDkkJEzVg7qKwFh3rA/T1OyeqaPjZO
6JEEKb1/cyfMrzifNwfJDPjSlxz50LwnVHHldSfLLBcqp7tCSw3BKGY5Ep4uEF3z603LGmG2Wyaa
WzlP38fcHHsaCAu/9HU93ZTSAajDBWlEsC9UlyIkXS57cu2DaSg0NXyRTW3wLc+vIk4qjKouYQbB
3fVb1W3wjMVIm67dAeUhv1RyXoi3L8olC2GP8p72ZCHN+6x1wawuKNdKk+GlkMK1GcctN+HmbjVY
6Hht3eidloOgUJRMtiy2zXNnuvwrEctrGDtlnC2PcfyC40ix8wIbnzzr7OtwCjqvkJ+15qFYYobR
RHL6YOp5ckJJFQN0svQzTXsfPPZRh49X3DUVxvCZ7Z6zmmlAcgqngMG+fP+r9ZJR3veNUh7B0hT/
gRIHpnVMBcC/Rx37DQ0BUNcfmjtRKEto8e1fGRTYmMbQHsD1K/To99hg7NafRZsJu16aS5fwbB/L
4qwzzRHjEUdE8Gsh6lB2wTWCOAl4pZ1qroIdFBDBRLqXancdaveaD4ut7tuaqvWeYu+gZD+TiE7o
O8x51KWW8+OtWTf2PDTMKRZ7GQuAPMnkpUcmnLJq9tAK703sLzf2DPKzJx8AwKLhJ6+fpze7lLLJ
0y47UH3yCIJaYLvcsuqiuXnYNHi501YB0yCqKcrn25pbm+izngdhoUPLJNf0bxL46clYNLq5zujg
nOQLGGLAuh8FQOrczbfpm5klXnvWxvyRWrX1SIBQNS+OgcXXAcCwdPmNuttr8cpLJVuooRo6Igci
2ozq6gU/xbdJXhBAzyoRWL+2WiDCnDTBX2IjAYt+E1thAmoOe7aBxQaCGtZUaYRBTpL6z+D2VPMB
nPkufqILUInznogdFHRjnFH6LLoKnAKSYwS01FX9LRijfATArQpR0bcXAxcy6mbJpSrfT8tkVs/R
XA+HYzwg81HqZTv9vqIrzO+X3Zdt/mwVj2VcVP6+qzsKxnYzoYCxwtWph8J/Pgg9G7S+PjlSB+PH
Fp22CTc+AdHdBL9Z6MHtLeSkvIaywoDY5yszEaUVn5qmZBa0WN3dOnDlojJxUGZ1PAYDeSKZf/uk
KLJ0vmDk1eBY27akG8+XR0PMFXZ5TCEggKOCRqFmMvqV1CWBRl2ShJLBDcYSDUILdlzd+B5msy0Y
wIgx/zi5YlaNyRItS6VldImeXy+MBQkpmdQX4v33Z2KBK8lja728eDBQmX7o2E8e+lzkYEeIJ+YQ
yXsE8BSZoiV32rCD7+4SPS+5++ZHDPXuDO7RujOa16VHqehzrupQ7PWQ2aWBn2VHElX/pMKbGRnb
kVTK3qKqmx2Rg5EqQzscoVDjHvU7rOyBhSU8SReEtfl3G5ZH7WA61m6n/fQsZhmDs7+MlIBtk5Ml
xgr4f04ykqiyWJXj+kC1CXh6RiHUjoFLtRMQepeUNw7LESB0Iyl6+1PPsET+/avNNYCTJoLtp0iE
ywaD4KCHugxZ+HyCMrALxLVg22MRW3IFe7D1bKzDPYWz9/qMf+CsA3Wjs0b8pqyL+zRaHwKM1vMd
FPxsLXAV6+iTpTdyrZ1lEVxlHRhqsv3qwDFoddEZT0x/+aX276fde1RMClbZzi7af7FVQh32IZbI
ZAB78vgT+lImna1azlMdupoCD9rbpiipnfDGXuPnQ+vGvz4xPTZjrvn52EYq/kEQKd8gWGlvCWy6
iPbTLVcJ87UNC3w+EdZG4H5LwNLQQHKOZabw8vFZqSDaGMkY1Lm+oxEyLF9tre++T6UcHMY9vdBm
X7kpBbmzCFMwePj1hQYlROAqqdbiIwAryPQwPOn5rU+1yaVLv4PEn7PmsFuj1hNj/e0ZutmJ8n1a
UH2ID6VQYqzHnlbotlnXjOm07u8WJlnHvytHGj7pti1mjpSQHTY+zClkfrkAfyXNIdaIt/NFNMdq
+F/IYLoljVhTn4QTaKWv8Vhefg5M4j4tL019pSfiJlaLi3p93NDtA55xEm87x7h1ZGQ/OgfRuK4f
+2vfmsAhnuDhBTRODEvjvHs792Q/rdrVrRDNMTSuO2LjkNPHN+XyQAPQWuMOAPR+4LfShOtLXTlO
awnRzJeXra+/4JMMSL0j6DsTv4LwYwLsJVf3ZCdFlxTxdSvCGdepeK3eXs/hZ2PFZ4vclvjnZrte
0cG9REUR9rwMFyMIayUDQmm1Y1OOmB+c8nfvmXDdl8hPQMozlNxU9nu+Uah5H7GXmQot/QGeCiiW
EdzDSYbLMVWXKogbPbNLWvYqL+d9cj2pRg4nWYNV7xFLEsmqQIlEL8+7hP7okUmLtVMwoOUfCWYs
Ard6dhPC5Gm0HkP+1GSlGEuHjp0u3gPUmgQhsMGCIbGKjSPxwP1g1/hnN7bpCuJBd9nt2H07hjNn
XnCDq2yb0HMhJ7h8UYoeAgvKDR6S9xleDDURST6F4jHLwvpyXpP+YKcdar7zO6S1N6jN5wnPglBl
HCAkvW2maAck5/UWL0rNxZpNocaF/q6GOdTMtSw3WCuO6jae/+68VcZu8B5BRozqnajcddVgeaL4
Km+DA+VT8ySasTPjqyXIwTBw+yuQFuO/g4orAJQssS1/1JLdlM8GjQLIOH00nQuUrmYv30+sjAx+
s06oF81JkSLS1XM+JVeYuNhbEC2c5SIVmitNJTbTRRoMCmdHjs1nfUkwp4rI8Kc3qi9LYe3rTyvV
tnLvkgeqNEENnf3zmFEuTZvsqMN2UCmnaBF/qXb5HwbT74lkK3WV6IOLwjeWo7NBe9SboyIIkVBu
x8n6wBsZ6TUCjKihgaRYgxGsb2s5NnVlqD6PxfqjP5uu0QqfDrkMJXQi/gCwnwA3WE0TaG46DChG
QlfiSv4+xHrk/qWJsKfRmm1RhQZgu69pkO/2Sr+YblKKAQPMTgOpkRa4YQqCyy6Aa012ILmGTlDY
wgwmbADRwq38Ni7C55uSq6tXtc7v2CkAJoda/+PqdoXcFviU1BA3imAl+Iif5VCU5TomWGGM5NeO
2Bl9fQYDGd96jyEgT3jWbalYQU3LlmsUrahOtjnSV1wjrf++QaB71dlC5v56rBABnAXA7smrkG7G
YHAJZH3n6ZYtZBtR8QW7UIIV1QxBb0nGl08nMJuiyF99Jeo7A33kVCKdOj2q7Iouxsy601zGM0pK
wJmo5SubFKVINFLvqpmN/GEm5pZAhD9htFI2tUZJ8M/OHs36UmRBiC1KASVxpe6ZIwCMSRfGwO12
7KOiQ6UXtMAh6FV0TLYPfNKA7HSfQoiPRwIia923pH2ZmLbCrbFYca+EWU3oOjeS3H0jMKYQjD7r
RUigpyPmfQfxYqCwUJCQvXNX9Hu7joWPGLg8GwtCpHnBtYbXtHDTApFgfEK9HZOpY8MMXRqoWVxk
wwcqlV0ytJNHX6dItkyevZH4pL/6g/3yGH9CDjLgstq1T6lFUJYJGMYKDY9/fdBBFyEym7KNTMGQ
XwKbRcawdoRQSQc4xy8KDk2NyuXX5R/fQdUcd4/+f5eLj8ItCtCEBul4/oTtbGwbCH1Zull0HVkZ
tViEuvf74HceSNkIow9cB+7v1jWnQT/rVUKR30s3dyV2Axr7r0ufp39unFgWiAJru/mPHhSnRDrU
ALKbJgKqxGegW2OQ/z59wrvZqnGyumJfpqPJGaAuS3uOU4yCKpJT2+mAv6eO/vFdON6NgvrIxD85
iHYMmibiPROjmhCiv7+IA51LdXczTcp9TYlDq4RtlsGLvESN2CfgV4bp+XCTNPpr6EKGarMOIdA0
1DnfZgDDN3KTpn5AHBj6kvhBf+pRAhmlTXhXerpFso2H8+KQeqTujSTPWMMrSDrtLOI5w3aea+6Y
t4S9GRGf+K/A6DxV+OrxqjdBFXVker6hzUBtFJIKGzmFPneEUdN8qeYE+O8jH4ZnIKbyJMWl2djb
erGrw5g9dKu5Yw4eZ/LX5vqD7+Lfpolx3TLJIho6FpmBnTydSdemu+rjzcibOKwqL55bAM1Xs6fU
YNQHR3Z4FQS5pGbqs7Mz6tor5PG5RfJ11K0P2OwuYbKAoWeVgfh9C+5yv1UG0uGYUv98GSGXlNdS
tFw+YjBA2e7d+9fNKM6HeLn3jwQsLF3yWDLCGrOJ8slGLvBbV1dBwLi98/zC9UtLiEG9zthTTZKB
FEWuIRh002RORfKQCB6zK5vt8//y8nQI5OD1nwmUSGm51j0k9Ra4iAPUoT0rEmcfyLcuHX3MdXSC
A441d4nL44KXABVi8Spl/F151YF8TaRn8spRm8EmgF3AIfyfNsLycrUWBmlwPJ8c/rmAoSEe295o
wiYnx/I8sima3zf1YnbZwbS9uXH55/JN1kuy5+SeTaOw5cyphDRfdQzpKM4Yw7owlv2MTa+P2CeF
HCJBhW3MmfUXV6T+SNkPPCJbVhKA1r9xLXhVAFRC52RKgxHQdUYjHd8TrlZM0BBJ1XoTle8UxwPR
wBUXTxceiv4ZKLbXPWYPlHeon0/HsydEPDbpObf4BNtfXm0QCNi6TuwzJC5Urf04TjQQDr1OQjei
aVBz4fe1TYUGAgzuN+T2ji5yh0MP1ZQlpNKSA/aDYP5W5D3KndU8hJfHQ1663uy1akKY6a/hi7pf
PNTCUILktiZHcL6C+5efdrxgIYx+PJJo60Fi2dW1Lb6kkCuX5pcKHiBzaX9puAdoMjU2LWgH8gap
hWzOAqGIsd8TbXW8W8IqNZhWgp+S7Se0xI+9PJTbncdaN8GgjUQtgPIDg+9BmIz55ykilHrOmG5d
CzMNisJtXChzdvnuf0zLPCIBxroPuNVObRXVfoRBOls0kONx1BxDof9yHaNWmAyHBE4hBtM1yM52
aRjEDZWcn6HNmHsLEsoAK5/baRPp324dqMXD/oIhJ/F6mjUWCf3Z4PFyLQVxB5jKLcpgjUiPcuxt
qOWr59RUQa0JmZBnv7o6k2s1WxAwyjZC7DJgJg/XQwlhPPgtJOD3TVdixpmKoys/7x8og9YRsLJp
TX/dC1ovmY+hlvnxBFCMiHF9uN9ebhk712C0g8x6n5hafyNf1NsJvAI4YHChxwCxV57nn3gFvNH3
VxRT+1+ymzUQkNz4nrYucvVG8VoGHMYl1z88j5YU8lIH4ZzVlV95XXddsX1UIbqC8P2QylLBdUyF
uC4ZKwEL5Vff7OjCEFLo4aYTFjM3RfPrjjuqhzofNnvT4v9m626TW0jc+HErLZTBq3spze3R19Vs
Qde+v5CjnstDeVlYTTOKyv+6FT3NvflRvEAAncN5KGRDIwCkKpc1nKr8pWPzASo6Oex7+UDz1SEK
A8gu7fJsnZV2oEz/0Q8sBITpdlckMjysdFEJVPoxSaRylTkIAuvAtrxgKtYqkccemIwcqvT3QBOO
IdI7ueIHCRspl+1Ps+GFqMwhi3ENFfqWy0x3EJPJEoeixeL5HQrP5/sMJUETSeJ35+UoXWusUAjr
iiYTNEnV+5BDyackhezcLx3G2T2r5j1/VeZ4M2DEbYrvrxCD6OlHRJsw5SvxWNwsJC+Y03u3wKnB
UC59RY+68O2T6x7+DUDF+LdYDb7b9uTy3kZQoAajrcLE6k1dnLL/FXa4jEtqPMSETuNHWcUwyMOt
KHHAjQVMVt5PV4AjoXrWP30RQBZ6BvJxXECe35jVopLlH9e8IVUutvAnMeOmgKWXeZZA45R4QK4Y
ZM6yCBwwntBeitT3vJzJ9SNu9Er6gmqs+6i6AMRndjv+Ibnn/6mMeq/sp9p40pP0C3GcET6UPy6X
/X3YwQzENyq0eiDWcmEyhAYgMadzpYoffY4V38C4XfNRpGMSqU8VT7foU49auoUNSuFAcWWeJpsn
brygzWEetzaid96cpq1g6iq1ZMYddWbOj0NuRP/kXkYxHiHqUkjM6y2+AmFIOWoYuAWgYijmLHiy
A4LubzVuD/6v2FDlv3b3uwQWQMU3En3Z96MjSAQ4ddcRfHYLmO8KB0hYra0mgrUb9sxcBM2tSTKZ
x8wwUnIJKcOovLQ9DD/8q5/MmInh6MbWj9FG7zPkAzJDhD8Mw/R0U1a1r6oXL6nmtxfP9bHC7PTq
5sGxBnIFocJeIKXJTYWmezavZcGRtpNN4pJZdAC0Wk4/rRDtm2DsTTSVgrTHPGqZjFk1oizZZs/w
FG/2eB05w3CrkOoMO1Btsv0dFf8yuCwAnIq0+6cwrQqYQ1/ugv7BJSRWV4yNl5Exg+3i1DN62Np4
yIfjaA1LXHJpq5AfgI8pguwWD7w3QYV9JeXRP4FpOP+RduKr998+zvWWtzDs3MQ1TpSh8PThUU2D
xoNx2huDti3VYEHzgWBa0V6+1iyiP192T77QVUXfrPRL1DtKoJ0+YR01qNmtuhaTXKpMEta51xvF
DJQiUyTnwLwQ9K1IkGgS4hEp/+ceDTC4Akjh/ExYO30fgOrJ3Lw1Kje4SISQICScOyVYpMy8zGMj
LB0/cXWoMnPvcQdLfPC2BeZW0J7zo8/T0/9EHeN8zaokdmQEdwlXf2iczVir92lVqhAlgOjIDq0K
BADUDrUYd+lJ+ffuXwvY4CsEt84ZFHqKhYsh/nH0LOo7vuFPMRrf3M7IIHvzFk5Gg3CYi0hjHwl9
hipy0BYBRJR/GU+9OPLq3oDLp58v4hSbhJbId79onO7mtfinHqutBLRjcfgw5JQ8geyQ3CByUhK9
KBT9TpL45APdXzQ086SSzmqOFBn5qAc6KfPjKezqdAlIxteVfcVWcFSZgj6o5uI9AraRyvoO1jlO
+FeZtsr63Zr/1AJO9EXYdy/YqCPgFe/3yElyxEDnUWJR8emMTJQ4MxgSuo4xYmaH25Oi20oi5wNj
mOjZZVgVn4YI0NssK0IxAel31zz9I9NdrVd6nH5TMmXCgCgp3vBEZfUqCffoXX7oQ26ZXAnW9Glk
q20QV/QLVkZEaMNql7wL9i1AyCM7uFGvcV0HpjA0uNmIXXbA1LW00jUqaA/vUGdSQauLHu2RKHUu
rW3xj9qbTKfbqZ8Nh8IEh6p6RtObkjqYDsj7nDlmnpC+hx82DG/4QAbxYRTC3pE6CfJTHW77Yisk
DTB+51zQUh8Pr7+cp2f4zknRvudEJq+6s+JdFloHYpRXJAda7O8EEzy3Nzq4mrECmGqejVEPg1QI
/jmpV7NtGqy8qL05vXPRZtnitgdDYmrELgDFfAz8AJ2WKxiUadxHwV4528NednRs5T76YV8UvlQR
mcPoDf4QF4V8Y1E7YJU2JUnzUs3t/LzSsp8iwm98t0oQnfANYNUb7UIa+v7Z1z2eMX6GhT4dHxKa
iLJBgIGw+YkUSm13SX9Q98Zid3RoNbjDOJQTKsSzvKhI+0KqEeL7SbVc3x2PJoEBoXUfSVOXM6Rq
UUGLteCNXWmUZ3vy5p4qq/ons2EtM12CuGvyr+u67V5Vz8wyG48P8qp/QYHqHmxEapCd72qcgggi
/JHLMvPPWp714XG+1PvsHhWAZoVt+/1kyxNbahCROu5dzeFVclIZuhAGJJadVGoxveuoTERy6U2k
TfZcdih0l8mDLESSHj+S/he2zJ/s79K4dom9SDR3sSH1mPzD+UiyXq62Wt8FEIUyoqwe/41byfhF
qDhnEY79mrTEPw9fG+HT4F7RVgVwiKySXw2tjlgZZfuIEV+oa3s9o/hxaT62zXBruDMXEozYLO3E
Z46qcEVJosJJDwdMpkDzp7b6+7Q4UqTcpL0BQo842X6Zwcw7ATwPagJ3jEIbmCosLo7sVWqk7By+
tJUyS6DUYvpXQ+6X/4VIlw+kGDsLE5aVyn1kOkFy1i3Ya0HWxWMTrY9M5cyl0tcGM/dyXNwPIl4J
0/hm0Ho+WPPJMF1M00REUuuWflQFD4VQYifYIhvw1YLdDjyRsCWWpsCkqQIq9C8XhU0LTEtk9XKh
PUEua3XCsMbb2A9iiL8ieQkH+HhdDYU9v5nxyE0xuZXbkjj5ZlAOvJP+dvWPPgYJJ4Q6a20qeFG/
i5M9xVqr9F0V+tlU9fMxGZsIjf2vyqkdS0z13whZH06Zi5KtdgAMrSoxP41EiPwUk2Fwx7+DLYtT
8EehQ8MQivL3G/dd7ieWcA8lrlUFjB9xsCIvKW9GZMM3Lq00e2yGWeP10GvmGRskvmSdCFXa5HsR
LCQBhwVUA9cZQ4gb6NzWE6pQV6fuNlGLpe4gO0PP+YULdMopk+d47qjwH1MrktQHpVLIxpDpsZwC
jEG4wMi+gW71WChvB7lzdkZombrHALZyJujHBO9pWaoLVVA1BQY0FlH0HCmzq7+qF5bVmlhVJ9Z2
nwNocDvOVF1mi9x9jgpUOsIHX4p/VNyOXEsSX9ZaH9N29Fy+u3hptSQEu8nleRrrdUeMoZhvV6k2
zf8M87WHJDwKGhGOobDO+NgY1UoyZxhAXU22rU5JR+YZFaq9sinLi80grasIjR5BzJdD0R7Xr8Xu
mYUp2hGGqhZHOxFJpsp8Jx7kkCVHH3NALqgEch4OPY8jBe29NxnJZg9qLDuI3gm+e1Xmq6sP/l9h
sTjDv/yXBMz+EBX49zRjBiy2W00yJueTXPBodbtqwVETjrr63/pv2ecV8n9WsOTApi+erTNSmOX/
RvdE/IR24vZdn3tYlczq9g4BGqcHSfcAry5bPmMJvSrxhDsuN9a2wAmTyqe36DhlRIhcyQ7oUHpI
QpHMqGuAHLyszAy3vQ1P3llz/1tbYt5fD5idOzbx//tMXFoC3rHtnfpP4HXp7z7rvDY5auglQaBJ
IdEzuMLFyYrU16m8bdl/j0kgfF9mA8hASDKsKth8fwlpXZ7OKKcSwAwjO2C9YpGMDC4/vW2igfM2
J6zbJS3DpwYzOBcytaSFmuLSmAvlmsHrsQpm6mmvhQQUhXOZcZKHr78fGgTbYNdkHPKlT2HVzOtK
5ZpQhWzYvlCeW5CU2I6RmJaxcZNINBlMpmJyVHXYXLp88TBb9TdTLFnAiwoVacg1UZT4kzpZV6G8
BsddosirNx3zn9Z30/kHkd6YuJd9gqutJWLYu9wU9xvBWvQdmHa9/rSEQVVy2IpqL0ziItRXzAGM
BWdQuwGDP5pAI1XehcRdA68FGC7pUQ6mYfkF563qIo+ekpYD/Spil8icjP/SvGfh0spbXWHqAC/s
2PbyLCYXpP405NNfB2nho5NXtkIjbcWgm202slLsRLU2G7DJaxn4yi8meeZPzVKIpqB/1LhtY+vz
m0g5xN/LF7Z6VD0mQMfl9r7tFtrhupj8SIpTJC7lLjodFre+iX+ux8drQCCxIw3SQI0Ta72oMsRO
rfCgy7t0v5fVEFYDFYR7OGj4PwSgiePpcKqrOvrtdoDyfP2lKOIyBbtk6CuyuT0uh5NO9+L1A2Aj
BlTML/okfKcR31Mn4XXKCUwT0LgS7LUgXnhtaCnRmfmtZHK859j1gfCAYMkqgx9O7GVrqVQwPjOW
2iDKypMJHlvstH5wNYwvx9mdQiWxcGsHtn92j1wCkqEEFDb2ccbszgXZt3D0Q7GXJEitSufSDVgg
fEmCUO4s2FNzRNvvAdKC3aFf1UX1EkBQHqp1NGuNlYos4NEBgjih+A7aPGb0m0xfX4uAaN+LMDRD
l3YDGaCCudZzNsw6SgNcarAM1/bzTogx0v9l5vLQosrEdW1ciEYLTMC/qUXe82RsEwNnZsdURi3D
YVD8wIChuZk1bsuGlbceafEiXTNZD8vfHWAQK1KtLM0qa3VGXn3J6wGeSyITSXKWGt83Y3xqU7tx
O+n5i/5mmYPSerOST9RZsKj88fU/iB73QOMVA1mgGEwjcAO0jiJYIp6jdhfMipjByb3uBjfwcIpG
myC3HXnhkO3FCIltccC9GGf+K4ghOcelatSdO7ic+pBYOjeGLYp8lKPPtDV7yQGmv3ecc+b0WeNk
3qcUu1LYRboMyejd5oRJV9oztCCjWQYSxvpxcmOcnREK3H91/OO+2ZbBLARo3mJoNa/MRuuDEdsK
mfZhHpet1lJdrgf6SMLWOxCakrN6cb9n0e86AwqKQtccW1rFAuOsgyFE5u+W4m3nqp+VAY6TehZc
20iYyQqWRgcWxtyxI0Owi5RNLXjnxxPXTohvq03gTZc72KjoHB2jcLQh4vzYzx4VhHju2rvWRjEd
sYR2xEZZecPjZRZNzeGvtnfoShIGS6ro5CopQeBdLhSLm9YDQiCja+A++bjCZP32Gb7tgvQvx1V7
VidKc3qUJ5Cr6ejN67qXpq+JwHW3tiSv3Pn2GeicKKOXnwF9iEVVHwsIDE1/O1OJY7CZnpVy1uTe
vfGt32xvQ6m//EvOn+xpPAZwgtGqxuJKKJxX9FseiZI6x2d1KwPFdaZ8jzswPVVzGdoOHir9r+2n
8e1OsrKF0dFFJAI+kiKFefArI4uai3GbQf4d2GT0Sultwwa6/XTxkSorT+zQNdtBwVqCzoqh05Hi
Y9ARwkqP6bDYX+rCCEuvCG6tKMpk7Wg4NYrZWSsyWVCughcJzP7+4UT3OGMIiaqYKCNP+xcVAh3X
zNpWjPHK619c1OOe4+3xmxdp1tIPHMlTttTXFJwA45OclCEdJy96/hSeguEtoMstxuaIG60jWisz
XJkGmv6h2yJGyt3FwmspT8Aux+EdKLAPbWplwyGlocAlIXZvTamVbX2K9jVqr0wmVGdxkQc8fPL2
NxlTGgI5tNuy0GOXavbMg1jnhkO6/vCkr42pITI//nO+cu1q9iCOD9KW1lhSW29WIFtLnoP4HyEg
SH0dxvt/NC+NynIXH1We2xNtrYe3InIRh/nXHrH5sN8ayt4SW1BrvfI1tSvuAueKiVaUcI2w50Et
m+X6Z2aofxZ468GXyKlU/MVN4QkGMrrqKpLO7vpJ3grgyzinYavrgxkUt+agB0cIuwzurQttqDle
+lIOtEXQ9U4S0upsiaGxZaYrIEYCdDPROwrsVUY4nCDNthOmkk09K52dqCr8clFb8K4PXdeB+2tT
9Wlxe9vowT2chtOLEqMZN9vfFJoggLvyR710DlN0szyrccrdE+T+2VekJoGyD2A/zVkxOGBfX6na
SvkuVEIjjzea0nv5CkQ1pJDa9zLyvyyJB7BVeGDWYquJBTu92CXOPWHCum8iRM9aOpvaAFKVVaba
x5FUZJXn/yMhSlxvPtREo4A8MXwoAJbzQhVatNQYH/5jRHQtc94yGdyxePJmq51OttsWQ+DOhzKt
0nuMXgQtxcl83o+wrcYNIclIBygqekVjcizducOm9m7+FaywiEasei0KpltUucVTTDDoSD3QdLvL
c1wZ14RCUDacNB5YPllMT2iaI41gRqeoYkO4keooJ43AxZ16zE12Co+QbYZOeyx6jCrJNF5SIjBr
SH8dW52i229hNuYSzRFV0AvhG/c8WYGLJiIwe4T5CSxn828J6J6Ws03fkOF62GhVGnA+IykxvXyE
vTi19+ULezhO4YiQAkAYLp3SEKbOLSV80J2+c0ze6lj98jfNVhwNdWVYaUlrlaG9paXWxJJg9PY/
JMuuiw9i7IU9MWqk7uiwJ874bE1EbfmoXNPHQDgb/Ni6pXBHIBxOiKhQMsx3AOPWEO3vRQPdNfkr
a5/G5fSp8we2++1pYwO3Ls5118NAxwVQbBLPnvxYxgdGP73QZ3BUqOrWml9lWqARkcr4vpVRJ/oq
PgXOWiwsVeiU7g18NaAE08tKoAH5ZpP/Q4b0YeelLyw0dDLuE0rDS5bfm6NUhgcXziQ/hJt0dSOO
VdKLL11CI6dLMFjSfpBBtRZ3ngfiHFHPHoApFm1/IsxL/6koq+MekZNc/VT5yWbqwoygC4uvQYI9
PXpsByVbItDKL0U479yyLpe0CJOdtO7lGe6g9KCwfitz4dXMZxilVhGfFBKZ4lgC04Yxx3QvZpUi
xBiTeN5nXb6YESQjbqY6RAGRrfuMH0kcp4pkYW2tVnHFMeSSR7D7SQzTVkfRghNglNTx4evtQsyM
q2XstqwYZvXsXq+hEpqHxOCGT5Cc0KALjaEG+wiUquO4lS8HvFCjC+ZAgMdgQA2lag43e91z2dCl
B9fpj57mi503Sm0u0pROBMCYz+9xrJyEfuu2ZGl/YdDsUJgUxAkCMB/nDjnYH/YIbrug0H9Il8wx
ACHJPJ5bqETPzO3YN771Xb9jAHeguT780xl8yYwNDg7ZT1atBXj/iHrSOziIJCNhZTo3VbIhhqqs
qIzfpqUOrIQgWG6RwuT4eVxtn+lwlCJyKRYFrM+SdZEisQDBGt/qCJdAnauUZGIXFaKHG2Uh7Uzi
sefKFSTSL7+VKKuO7SFn8z5HvEfzUE44WbsbuZxwEkazyySIq6KbP/3vu2ve6/TWPPE6z0Mge4c8
9u2fPaYbDJuG9IgqAmadpEYgvn9Xd0+mFJxcGHFji3KTBIVg/BL8URfW2u15wbCepRaKJt1CwrXR
UcPqcxHTpWYqmUBsXXPnqLIOeMBkkv/l3/BHoS4R4/KS9+vcraX3Z25I3VdLqT6S0Ik5q+Uj2plz
vWAsN8F3bA8In9b0iJFwfYYHER/PN9y3ipK94ZLSdIeXqas4Uk1KKTdiEyj1bs5tHz1ZbHG/xqxM
2m3V4KknKFFcjez1KPZONbAyEhocxLLSLsxuO8wnUmDb1xcnIqNykr/pvGIH6OxMO8/Wgh6B+XT3
6aPreumkwmkz+o407QR1r7SWmKQCeXhAUxd9/xk8BThuLpMogub6ab5u6XtoQRwoOZCnsOi7Krxi
oSI2sckGBLUtSc1AvIhX++PWyLZPiert3J7wzng4V3m+oHI5pyUIZO4f0EwKwoAdoG/hFQyqCaRm
m9NyYJceejrwIOwg1eJf79+4Gr3PhYYWRrz3acSZOW8teqphIHE+qx+q79AunKN0DrLWJc7AejRd
L2iCi8dnrVnHspKAj/cxfPnUHMqx4Nj08Pn8Tm8o3Y8vvoSsXNadZqGRliKEnrtmwdxK+etk1zdL
DG/mifISw8w+F02FwkZ5DWev60z2s0hSOtIJfTV+HXV9nVIhXNXN7gh0gNmJbtCsUZFyXHljIgbe
X72L6g8EnSad0sLGb9VVUNsx0t6/LvCUbkPzatjpPrVNyeH3Sp147CJOGrZQTkTsLyGIfEvMtCdh
ge9YQFBfW8cjzAt8Mzw6G8x7hScFNWbCXN4nX0Cyp/NhlweWALaHWo5swLqXX40C454eZA+xbIEA
1fpdQRqt2+Mb0VcfudDihaw9ieelmrt9iV0O5MwyKrdkUJ/iMT4BeZQHuIZRupolJWb9n6H2EzA1
brYMUcMuhiX4w9wuccNfhm42sqDmsdTxkH8xQ4ozoVuEoaqsG08POKMx97Q5CGKtkgm3og3cZdZD
Udga2HoJB1tJI/fQUi8Sr2mg1ZYjGHH2IVBhkK3dkAZUW0kpqIlpKfS1DzHZlB7lcaJ+ADMR6Ikf
tQSkUlD1E2+BM622WNDW7NzQcU+m0GAC6r79yuLI9VHZ8R37p5zdacCjfVW8L6fVExVqeo2alcz5
bVcyLOxgaIRbUVDzbxFTIrnjxTtcf9mTGGzJw5yGAkEf1EtJTa6ypA8/vUtC3OjfW8D/0fv9C5vG
9ElfRD0SUGLRv7dCOKbXdR1uEnIzOV79VIY8ceCDvkiaFJwj7BGsDr7MP04hSW7fL9f9aKC7eBaf
DK9FG1vlxSTTkt1F7fgMqrm1Zre1HeOCznnIhM3oVyIgClTiU1Nr+Fh9/powrDHtuH4IpnZ+azX8
oQ3cdSWBpuY0yKR/T+Z6Q6mJG7bPG4GG9uS1ZSumIBZEltlLOYwew3Zqxc1FoI9vBJsbqzdofDkw
cXqRE9egaMz6PvdRZBxN9QYPFBGHhjzwTmtYw60ygEJEBVdfYOew55szL2rpmzzP5jD4kcbLyknS
PaYvEtqJN3b8qZ/uAAX9LEFjD5BLHXFSNk0cx9aZbuhLIDuZo6MxhwZyV4ovxOFnZFcEZrzZFvcM
TyhH76RnKMbE4WkNi5Jb6wNGkYkTQR0se3uJ5w1+3Tp63XSA0C3EyHhV5/JZBbfjXmUp5vlNMHgG
ZYIW+ah6yJ/1djEzdRACb31I+MbZVkb80ZdFYiSPw9L2YP9c8hCQLX5l5SNVF0Y9YKuKAiDGV9sJ
prKO1dml1B847ak4838f0vcmdInQIsQgmgLDmq6bkd+HHI5QrXzClgumNFQdvCdhTfQnW6cWxK4c
XgguMl8zOLGWImcixaek8cDkMHcT5L70EDGeT9aUcyWgx0LxY57BUbHV47i3yChb55By46gv227G
1Vk5zk9cE/+RYQxYrkMmkZZl4zz0Dtn+WWW20608JxapCYEBrncPgsKf7ZSPIhH1HL9UDeszlPU+
q8SxGuOrOO0m0X+clRPmPJU0HA1w0cgtDdufv7yM1CyNmjXBkFmFbkfcpYbk1mTcq6O1/7Lm6UTv
z2L5YqH0k3I9SLu2dIN3CMbTGbcGaxO8e5jKTykbbjs7ZG2oG8yls1PubX/912g75hUbq1nyuuzg
ctoRSdQomoRbiaGnmwIOZVREbwSwAIS8EbfY4YlGYMm1iYjBwepGgnTEFgc9DFzFCGnltBTtqovl
9jHKazgShOLDVxb/5Qa17COrhWpkzIumQzjw/+4KwrWG+xvmxEJR5KmrAVhpkxMBG7nVEq7t1G3l
mZtWONUx1GL2RHs5PN8jR8wH3vs2xzzxwUAwYuE6U8Dewm+GI9H/aVH4OB/u1oiviK0dKBwwjBw9
qB5DJZkyTLJXkv7uT6gBLao1nqvt6cTdSoImO2GzqpfTgYFu+aIwv7fL0JHI/oZqOTeYvQiQZLqG
4toLwiNhn0bw6+RiKCupo8sD2YqPGHZhDk2TuUJuPMwWrtTxiXYYx/+HZQP2tixGfANvGH0+aMdb
9b5+bwhF8u5cR2LsiqZvrEFoOK6WFc8MLrhOijOipLDgOKd3XDW1gkFxfZKt5rg4kchdTiHaCl45
zubnXtYWNyhx9WgVCVpfr6Ybc9MZtytOotBlTOf3i0P97dLo+iYByyF/8ikFQTfs4UEKZ6/QPAMi
Pm9hiUm2/IK+g95YtDZkPWKogD7vVnAmkpXhiv0SDjWNanWeNQeEBDcDw87MhfouTDIt96TQ2Qb+
LQdvc3oF3Yde2eTyx6LX51HIVQ4p+IzsI7ndlNgPlz8U9ocjMTISQ9YCbTiN4bgxjbGxBV0zY4AL
K9C62WKXy48ZXHAddudS99FL1uxSadm0tEBDtMWbL5aoygBaqRElP9Qz92pLRCeD7hyHv347ULDk
hr9TpY7VS8nzqh2vIHmIzfhx1NE3+SCL8fK3w06pFICGj3E6s57ZwYr9ldwGxwVXMmnTdm4QfMAT
nCOSRwPZzRUMfpXru/wmEAQ8cAOoN6pjGuJimlrwj5xEhnSeffI0uwxeEnzkeIWjTdh6gF5oy32k
4vPEMNQwRblhFfM+HxMeu+CPE5Iy9McDTxCUdfyBLC8qy5LNvYi6oSMCYfeGUDFbmY4KQHECJ08M
L5vz3stlIwwb075y3kgmqsNQ37dEplMtODo0UUIvNXiLReKLp3amsnmtKDe0UB/yg7Obvd4yjKLl
tYwvW0qnda2DpbDa0fB2AGcLiEfBGT1P5tLCc2rTuJlAkMWd1ewke6Y6olFLa7ejfyKvhi2lPHCO
s7OVWBn1z0Y/ThOv76hy4ArlfAY8qqOsc0aAVgThhIBCCnCv3Vso+qkRmPAWvI0Srivj5nW1eRlJ
CdaZrB39f6Tqy5guMOY2mrGCGRIr41NVdnTHUm0zJlLPFynXFIl4qeZoAu1CeJG6UWK+my7a8ZrW
foSeWvlSsDWfT+AypXFtUNBUPaUH7CthCyx89GX+vTmQLAvK8JNifaKvoz0fPC3fUJ5xMvV5mR18
Ibij0ibanCQ/4o5vaHPgEBXwlvEOkPgSqoUK8haKxY3DwPfEZEm8l6Gjlqp521un14m5Np6iCave
d2jalK4XtIqk9TPkK2SQQbcyvfzSB1TOkFM2tRMztSzyluiGf5aS9Fe323cl9SwxzaD7Z0v66yTH
qseLC80uqgiZrFaB+jWZaGpOvyL2rwlWLmhGrQALgWabtpsM+es3pZwg1GAmLBhnaZR19D90xJON
cepV9Be0tH0dMDsWwSdfh+Ib+WwPQ8CKDdBMZeLk4QU/p+H7z+LkgQdBGKByT3wd3EBZpF3Xpjpd
8OSlphCbqIjw+iEgvaSWuy4tkqljs0l8yvkk3WdgXFfLYU2nXHzwpyXHrvd15EFqnZYm7y59VTv2
QeyZwFcSzVKkJyouZ5X5De9kCBzbSgfw/73MiGly4YqJG0/pTVndK0fARQbLGWPLWqsUIfVG5EYJ
kgM9RVUUscIictRUsd1YHPE32hiEflba0yWmXKtPhKALcbeSKaVvkIiyyg98deeOrT2Adpr8OOYE
888oZZcjA6BUSbpjCtopmoddHOL3KC2kipyt/tkyg7LXR0fEvNaYd8+dz00hpBx221APFRRD0U18
Yw6x6dZfxItkG1Z++/EcNHaGmKLddus3bgq4D4WyrDOOJv/5T3PC08gzCodBP4m5iNRiOFO6qvsd
YYz1H5wcYtQfjc6lBxF77ALQUJUW8p96fMOtv2Cc22y3wFrMkIuEk13oSQVROCX3lvnE74c7kKMm
EAIwOR2EHD36NhN8ExvuVDfOkKFYNLHJMTTOZvhVWezpE0VuqQ5ozo5gQ11ryYAbCbdZhmZyR2sR
3JQ76JJMIypTBnC8VJh5VkufM73hNwo8R366rOy0h4/GYzT4T9l2mVFhoRhBzz6UKXh9Z/W6ymRY
gVR5KxMHxeZu+BunP3A6oblqmR4583JLcO7LSIR36h/nSgf4BJ6W2JngYcvHBXb3kmBxsNX5v0Tr
GaRCoi2xv7TOBFfMPjG6lguvN4pY1iQFrSyYI9BlwqFmVmiUBOEGTDTzPjkUwbEmGdSL9tFtbCGz
QQmRYZLXRNeB6J3JrWz8TSda6kwxc1OanosGaGgqvFe3kSzOvwb2Xmrbt6RKYIFvG+Bb5aTwp9GY
/1dq1B31mynWqX/WY1k9weOTgrSy1jkGjKmaNZjsIJfb1AU8Rtc3mxhCaSZXuhJLC40Zrbf1Pj0r
OjxvyUyjEyorKzEYqdoSxPxTqXzoT4AW1c29Rxc+f/fumu2+TElHhSM/QJ7kso6dI1ZubY15OI7W
9rkgLeSp2kGgG/uAqe1Th3X4VxMHA2SOEibEsjPRhEiYj/la67qdV1k0R+oGalLoAsewnmT0a7F7
tXUXkfCLXgK5NXAYlURkNXOYsWb1ZJxLaZTm8gLA8mKY7uGWvKY95ogxsVW695hcGb+aA3RdOkV0
3DSisdFwFlqdBOE8pRoirncB0TPPwtUJQlRa5q4/wyDHy58zhal1cCmI/4oSs2l11p3bTZeJqeIV
Oa+vWFa93+PpuHtXMGcX6Ewt8nvFcv0wFyy+cm+qQMUjPwM61JPgsJN0OsQ3Tga7IVjREqxb6KIk
WM1k62dDa+1RTjEmQB3blafpGaZWBMrxdspE2D1Psa60dZfqK7XB9PvzWV4K1wix5DFrsGDQY7Ak
AhxQXN1+dBJFv9Ra+PjTGY4tBDlM7t/VOtJ4XyjaupYcmgdZ1cQT+q6dgyMqPIfy8rGpR7CC9WPb
wGSVEwjiB/lxzTWcXOWjHPV5ZL3IJVW7h3ZyMRwbkibLuTps20zdHGkihuv569rUSb9wUAce/9JG
IWxztlD0j54xBKTjYbdhU9MVDbDZkFaxaHWjTTJK1Qn5TW3zJYwNfwtP4TDLSCgr+riRzLLy5dLX
TNfRj9anozyFHfmXpO4p/bOeLlH15rvhuLmtSoW1AuVq1xHzxDAV0KP4Qtuoq6jJjZY5rRWiuXUS
5/oTc/8kabQ9mf15QYnC0KEaoXBOnyZ0Qy1RITAi3yLBIRyyH8kfAdQqu57aSHk+xEcpdyfXsqMy
gGHdxSm4zRE67WBUBYyrQXByx7L88Fb/FO3nBy+eY37po4AP8Fwit5f28BdntMxTceoC7GVgFq06
wl35IQgOF0ufxiVWi1WF/mF0raTqQOc8/jLfKfgzcua36nobHHslnkHCRpamB18sd2T37jRgOH7G
KKFKgdALHuALgu9UyO/w+Dari/U/pe7JTJIWpWBNjIFUjqFJhVLSPG8GFtL2FTtraNAz7jcKZa41
IewNfqTNNNoki9zhS4+pJuiR0iMqPBuUVrrbovhQkB+c1ppEc7bkCASI9dgJAsz4vC6gTDiGkF2I
7pC22/Hzj7TjwIrO+B8V1IHm77zV9MP8WUYJN2rLlNYDkHwHMBsWaHu1pE/MSMSykKt+kTdm9DvL
ZD60pobnLc2fhVEcp2+3LQTEGwJL+OG2SgehRDgiBb3HwTFLJNOhy8VYXrskVdg4/d/3qU0rQ5ao
erLpxTS8PZTV0QrIavb8iSsqz4GuUC537IspMK5mwjzLPaw5fzv1HKzqkTamNDWLvAFzN4ik/GXl
f3yWUXWiWOmvKpRvhZiTcGgX59VAsOtL4Ye4V7QKxiKcTtkYjGdGANowzpfsqTBEzc0gov145RP1
XuquD+g3/S1fUcwRqQIQulTIBmDIxA9mL5hisOJ+6A0BuFGVZRJYf1+XP5HX3fPRdlJ3eknhAlT4
YE+erEjiTlndaevwGoNCf5SVIJNKnE5CsRprc2yLSHkAQfEBfBKBFr9DWJ6roMTWMTibZm7PC37M
IU1nx8EPEM1750VmcTVLhe9wUUdqatPk/bMYW3affU7CGJM8TGUc8NGtT6buT9gMdH6g2/bmHL59
TyouKttEJS6IYb8cVh+pmgxfgH5TyIwk0uXVtIYn+ZpH/wi0dCim1uV/az39QwjTrvTJ0ZtnB6Hv
clgi9yI9Z/O6Jd4Gm/R4uAX9I0bpglFDMJyi2s3kdJNlQZksTf0vlqmnlort0W5yN8tlvx4KpRif
TLJlkybBBDUAo1IZoHbAsHUqYYVu2gGKtexWnwDBPiQso/tnOllbrq+IT9Fb9LKyjfspxTMp1jLO
65MUAFTU6/ImYTD8zHJj6nSxksxpt/264JLZPEhql0IRiB3RE8fkzsEztytPifC5fAp+0AZyXbr9
MjSaCKMIZ8ZNBYi8j8REGqtDt+rgFFA8e6opWcUdJzLQqtjkTwTRgofhLwyCtNLLecgcC+6hFte6
LjSr+jj2cbQXWbO+vg6zTSPbXAr01saA1ZrbHSl2itGTT37SlJBtRnMaeIdv47vjPVsgdapWV2Xu
+v4Q8f/Jm2VhQpJL+OLRGTQFCagqraRbZvDnbIDgJWZCMh43Eo7LSC2oSd4C87Vcn7UGtooJ7rgA
eqLBFXy8M8fUINqRk/g3G3J77gf6igv0qA+tCe/LNlnks5FIZEMEIQZvp2KSGxsiQcxGEvE8gyKO
hdiNge8YH/MQlswRXLOGLOGH/lQ1HN5PEndWYwQ7QmnfOJzWIYptXOW24rAy/1PkMjKR+jnc+jXs
Ov+npT9ije6gatpqYgXDT5yRx9kvlxNB/4eDkZnOgwZqKYPLzv/jVmk2cO0Hi6dYCMZklXZAXeEm
8A80Ka4lN0+HnlNj6NYJE/n8Niw/jJ1c38dCWBGECSXLIrnNM/8y3VCFTMR09HIZ5/r5EFayzKsD
/8rQ0hsRN+R6O4rc4sfx8SYxQN5uw6K4iuux3SW5mxdWns9YVNw/No7RFjfc1QK28zZrLrP759fs
BOyH9ORmn2bbz2x66zPcxdX/bv2t6uNaxlipa6F3uLK8rifabh5IszMUm7XP0FXusWszyqIBew/P
rsu1iFe40mospnj8JQ6bKve2WooHecLy8GSpsn4Kd0OYhxCUmXUSmxHScbQU/ZMMBu5l//Ur452M
QpLijFOUz9nIQ2aZ0Wute/IiwM2LMr661y8C10/GH+oUIa4OO02mu+MPI7m+AlAAZqSK8MDrFWPS
VXpsmnmUmrvci95qgqHfczTSD7ND2Tkw1vR68AqOj941UwRqMwwnGOdoIbXbQqtxk7hwNY2qJ6ez
gkqGYBu3FtcwOO1GbXzPHuov4t3eV642eQqWjtds5/bkJvMCjm8JeqgkOAjDA8iY6wOrh/FRye6q
12851HE/0SP3ctO4qcaMS9n5dia8DpsWmOIrwD6eUnzfmeb7U5FT72KsKxexT7sKZ7FKg7GlbIfa
9OoHSY2pGncxokOdHl0df7N7veBnd9aPD80fA7D/d+COzShFYrkAaaMXFpBVCBtWZwChGDSUlaEv
AXCtmT3MBP5BkAfyjpxW7ATzFQpNkcCTwVr6/9+cSTquvqGJbPTb9DUHp5IxTON667TK0HQjKCH/
UHjtesTPQXQarAHidCBb7uhBz9PXSdbN0183VlGh5zA3KbD7C/tSdOi55Tt2fbgQdbl7Qm/50OHO
1Bv6TcQndpWbuHl04MakjJyB/SbDamtJoV//JFz8R+VRbJHSsdYFcaYfBDvi81ZbZLx+geeQ4IGo
7JDmFroS92pzjbzoe0oxYoSzKCOKgJBRe1/qNhflWIURzQrM7uP+e02g7Z/ZzTYg2TZpPdNyI3ZJ
TH6KaUNxZ3vNTBCHHVXTa6nanwdhQp9vrtBcDtOL+LFvg9TzNVPaGL//Yy8+ytlBRWJBIMY0h6h1
FRhKhlkll/7goY9UUBnLoiK4xxPnzQrC3/9JFdZ7Fb3+Jr5l6S+IxOn7SgKloaZlAaokjk3f8mDo
MqfCfmI9Wq1HRwgE6Cz+uqDiWEC/1q8BtRSnQ2rAq3siR9uE4yhNz25qKHvqKWYP5xrCn1EbyYhe
Cc8i0u1SYn9lzwc1SbRO1bcg5DcTrynljIfKrmOP7S8Fu8JY6R0zCRaGEImbByi9t84WTnRtb4f1
pXPqogi7/xX8hHS5K0W1KVq7cTn/tKr5Qm1OUN/qEgHXL474VsBo8Zxez5+aTw+epoufgr20N/nd
dVatq+pc240ikpaPPZQzXFYqR4F9tCqbzC5vzl9Dis1Gr1T8UjEn/LZc0/wZkWtnO4VomfVtl5sO
E5uFzSJGLpMdwL/cKVuQLio4/4w7wtCtyWMLxPVpHRS/E4dydl9OLrev9TgDE7fYorwBrrK6+tJx
O4dfwJueX08eLYx3orw9Qcj66ktjd5AO5y1uiaIPLasxfnYaYI62kKj+DO+b+Y8IUFcc+4vd/ME6
dwJsxVG48B3854rg9RPIamSSE+BL2XZseYA91Wqg2jSOHsFohaXQ7SV5tkoIH7eiNePFWC94oOKc
FxREUq3WXvHiVwcBQnnSmVWfa7FcBquNSoH8GWrY6/rbbsz+Z9haHAZVjc86da2CGMoZ8qmzCThY
qsI4wxDbTpBAwd2adyjWamRXJM9yL9CWGkXA8zNNHYGvq0eex2nHeqffJ7GBlcY6LpWc4Y2yk8rT
ls5GclQZ0BS52iaa5uOK1ybTayKWduW1Dy+jN8YmYyrt9dO00gLofnbL9Y8BrgBEQUDI5j0MmIwc
X0ORCuE45hFWIMc5XpOdWQJ1In3LbWj0+DY4HZvWyFACcDpfjwzdkdssG/KWBMaXh83kdh/uJOAP
U+qUsExeY7tRJDxo6ZaBh7vVOT0Y3gYQp5TVdAEOdztj7q2DC9bsXSkyGk6TF6gNEGHYZSWWN/i+
TyHOGptgW6Nvqg3RHmEj0ZDQ4k6VXY8pwIQwZbufRI6a38CyOATAe6ZleenLN5JehPOL2wfq+COv
Jyn2QutlUuxkoc+cYVZlhhxryA29RgO4/A1vVez2OXqkcAIfvVShtX+mSOwdQix376619wTY1dcP
0Iqh8ssdscGwBQb5tjt+fmCbwjsbFkO6e481/Aa7FvdyoWHE1PYMLq+9UB4aeGExCr/xsCPHOeMR
zBlxiFMxL3WG6MJGG/WGvscuiBFv597Ddf8y1Fm5Ke3PK9syF73J4abWCr+494LxGnFG3MO6ydf0
R6wSNE2Avz8BObQPEf2my066s8PvENkAV7lBiKEfHHIbIjPGTDzqV/EMGOpO0sAHk0h+aXvzkazY
N1zCxQ5pYdluYdbcFi9hakst/UGsv5i14Yf/9YhvMoN0Mp/45lHebzPKqilIvRqxI5MevznIX28y
2AgUYL9HYF78qxnR1bZNgBbAprSh/6BUqtPymDxx72reXFjUiaCDzuKBuoBHKD7iY7CJl8BFjKSI
az354M32Zy+wYc82/D5qz5LhFyqLiKWgwrOi4meiPP8oV8s0/B2TD07PLalHU80xvRQcxOcU5LM2
Ji5jBc6Fyb0FMl9VS6aZJaPsb1BP7k10OiAOSQYiChsXCheG1Ft83e/vjpX9xOHQ6XsotffFcRNd
2JNkFhLzPegY0Ds28L5nOjtDS6PCaJIihAwsZE7WXiqo5YgagMAudX6PvZ3BVI2VMC1PrgTsumJN
gQqxvZweI/t9lLorIrm0OSRppv5fNPgFQ5SbXgkI1BOk3sBWggNH4y3tS+gNnI7HWRekqfwWx1Af
0S7tC241NzgSptNR2nOk7H7V6U5ZIpkP0moStZJq6SPI1357JksAFV4FghriiyRba17tz883PPpS
sV3f5FsJJbSmscR53miamoBvH6jIhN8d6djD78p3oE2WmCDUXRIM53GBb+DvXJj4jzBdms640uDE
nRKCUvcxhnNuK7j/e2zIVLJqyoYpnx2qgPVTTAJJLJNR6IgT+TEZLthtskzdJnmElO/+ua3+vFUE
r9Yahe0ZGPYTAqoTBTUM0fre3ao2j3I6WDsbEYEBOMvj/90VUQ9TM+vdvVmxmQBfndmlikPHK/pR
DN5zRxCAuY4nJvuMIopq8sBWC0oOYJmg2kldUfi5qL7bQMTxLrLQovSfdN0RiNrSH6BUOV86f+eP
rgTM/vkfafz9ZYijGrvj7tVerwmWBtk+s+2e3BhGNDqpTcJo2h5CE6GEqp6TiWYCUZQYWzTS+ZQW
8vnKxx7uhh6JOpn+estDZaOYg77cr5XfaLpbdYm3wcr3ELoveSa1vxETIMp0mGG2tUefxSiegG57
TXjTrdv64n4w0lkWvr0UbU4LnjA0vFYpelYCQhBTuU0V75fXlsLwmLwyppJ7r+uEisC5LBwIFUFq
QJwIIF24W9WDIUvVXMtT6TuVFPfhTcoZ6r/Eb7zozEjEAkK1LTzrV0ZuO4YKA240D8sH3GHBpq53
YX02LzUAqyLndsRwHOPBNWNrljB9xU+if1VWIo/kn/3Z/zxc5a9GKGEtIZN2Ay3V0PIabYTDDiEE
d2lTbkVbX6AuLFWe6q4SplgJFXiYFP+rDl2D2PJ8Axy60fdRDYUUNnlmvGHA2Xj6wrSHKPEA1Arx
/ddhAxe6CIg5B1TvqbZeVBUI+260Fs3Uq7z6A94gjsjS5A++L5wl7bZBbsdqBBKKIQauOlCgvPC2
5XTooKU3AeYlhzhIskWnhtAYOGwmgkj3EBW/5+KuiOeYaY/TBEJJQMJsY9bO4k+TzElCejv+XMOx
9D4aSKmXIfbyDQqD5hos74rEUoEpGRP7Jagq5ibnPAZ6htuhZmKXctdNIMJ4tlqb4Q5/S8qRzqJt
FKnUsGO+YiNTSyR5w0OyaaHQ1FVdWU/2XgPmzxcgbR55TRx7jo5ppqfQNKoAXjzTzgesYJLdOtss
YPoeLj/DpZtQE4h5TzmtJpElypaPqOsTKKh9rR+06zfPnTPgHyRs0vDpvlkVV06sAo0yo41IrRoP
mii2SguOAaKQ32qRhoG99w0z3td9j1xm10WkUQTTa5CzFpLSZn2OdY9JP30NwNqzaIgEkjyQTJAM
qGf+quas2PQycDjqTOWsjLMLAnLkF1LM7QjZFGydiMFl+Y71Njloq//B4yvxwt/Z+voqynSBYY9v
ZXgO7aOJFNS3xD1oruTDpE7Qi+ds/vicLHKiPM6/66CzhbVIqsXBYe6tID0AO77eSYj9zgetooFF
pL5BT1RkClfOzWWtPEWyMAuQ38isbeWsjJA+U3aqXrnd+GrM7mob6GjL4lkZYBpJDprNV0Y377go
AZDeexQwPhRKdPi7LTTEEIFGZMe3+gAAazfjnN2SXUiiqY0FmbLFOkwatICverjrB2PR22MIX/bc
qleH7kwt+WajQvIyTc18R2XrOm3jnhof9wRVvugBSPx6hk6zMoYJrMawtsRZEZfl5q5Aml44oX+R
pibCnDVpLXnnfvTxOWexF0aUM02uW3vowc9QjJaQ1DLb2Ctd/1g+zmqbRGqVSzyTQNK17En4eEHw
Pz+Q5r8tKQ10gs+oBxrGNnRT84u3hnUovr+/pgiCwdV4IydmGB41xEgT8j19sMZ/7WQnTiQzaxaz
yZ68actC0PuIRnOg5BIz4cxuZoux4bZNiR42wTm1eyFECn+4lHuIf6QTehZVumBuSjXFzCi3Bfp7
0urkX72mO3gedcSB1CG/YnBzw2gYwsRiGVOVqE3HbXjBHTToOHY5uK7irsnPlrL2EbhKpjdcovGH
a7iLbRvO8r6wKypZXWOCQMh9C6MgK/CUF2SY0ZSLr8dpEq3VCxDK85T/3gRPrPBvQtOAqjab0CxR
BeHpZxZZk/LRFv1rspA9G31RoL53pKOt+pNhvwgVZKI0UMpn4m6L9HBZDikShUmCEPejscgjEew3
kkPuswprkv2JjyXfopapFQzh+N5FUwq0Po0+R9K914cQZ5Zl+P69sPypG18kevrjuxXa969LmNyW
mP2r5jgHQuc3hyE5j8uQoleiqdqq9jmBVUEsUOA6u8bqcyqGp2vIqbrxpu06gfZ8NdZOOnsdJU+J
lz6rrti94l/UxL0S52SVCCobkXygu46tzm1l0CtkMuJq3toPOCZbxjcxshaQOc+y6LDpHTTAT94T
25xB3vauj/nC48HpLtB3UYOWNB6VE9FdU3WcgvtFM6n1m+k9geulYVb2V/eXkXO5JNIV22e4A+lR
0i7a3Wy6cqIOHSWStw3wk311erMWAZjY9xgjRI3gNHx3PwRcBIgX0JW2RpyXgEj/kkQ7HozqHKLT
vRc2iTtOMSlwbgfW+qWta6hJG2kHydlyPZlkHoXpcSWskuL0mC12NqQt1D9Kb5YmMAZZLssSWAjW
Ut9msxv0QethHo1qsWgh5MgMexe8S+9h2uSiRNzhwvKnCHSxB0V62RnJuUMyf+cZVz+jzBHoUmgx
8/V26Xop1XttNOyAQHou13O4hyh/M8ydAYNvxYCiFyGCKhqmDlMVNl65kwUp4p/ArzYPbgqvPMLI
6jMawrvVn5zIfiJKOCYQU4PsUzcsn6H6Eml4DuZgfP6RhWXcO5nwxt/lSAbUBYWlca1EBLAkWvO/
ICqdJ5Vxzy8/S31MVQtH+c+9o2DKL4uunyijLxdI2s7WbiIxm/AyLOM4NNSGxR3UPbm9GBJ1sPKp
DblF3G8YjTbirPAsIUwme+aktp0jB4cOXFhZiWvIvO1bTHoJ2QvoJUljlAruQqJ2tw1raVQAXnLu
6cYjKEa5PH8bHvWbHA/EnOkP2bHwfPSobwBrvOxEFUVgTVp3wXr7p7QlV7hbi5jcn0Ec7EDYLdwW
UyMYuW7CJYtOVMvGcL30UwOh1+TNjJw7s0fH8sAb2RUswwlvGI7Nc4/aklpJ1/Od7RLDXBH9gbBy
4depXYqtv4gfguQwYQyE7/r3haxFEh28HxpiP9lzrpfBtYGSRkLvAJXOLGOJFUjPLxrJ54nAs0Jg
6Gy7ECSZ66QuG1DmzrbTfcBrIUOKv4V3eLY6CIJTn8Xx+F6IG6jzfoZUz8hs4AQdoXHDxccxOozM
iw6T5W99ZXmc3qWApgI2A1L/YLO95smy8cFi1Ye087H2p7NlKbxOhhsxbll8/+g3wD5SwQT1VDQP
1nYsGacqFFwahYuzcr+ftlFlGeWAwjU+aOUfedy05yQODWAJFJBopMxC5JrD9MoYvLlegeBr8yoH
ykAKDO7rNPk/fdwDhAmVf0gl94/Q4nXAbAZsBqbcoZqDeFolTnN0tYLHgqKPW7dbP1Q1ZJFYg3ZX
f7mOP4tFPpRcfuNptJx5mO2MuS5k87aTxoIRpAb2w9rwcqw3bmff8E0yD0SJqusSD0jUT0g3PqiV
tYs+Qps1w4nsrULxuEWJLfMDfRrTwLp3igIawoW5/6k9/0yObZrmNEIlJ4BNZG9dIZRmHMdiNt2W
H7q9OW+YTBclnlo/dJZ9xCGMG/TFgJOi1R+iKOlZJqVWyfCYREzplvNCpqxIwfmN4U0+ZUJeVOa8
4MtF0pmZa4/M1EqsK08XVC1wLhkNvaR4cAmk7fvmlmDjhHBi0vQ0giA1jcB83NmPNM+HB6dp95SI
LX6gzhPhKvOWzQcvwkFk1E4NZ6QDCFbj+pg/lt4SpcztP4esNzCca9LbRy/kmpw1yLqQSEjeOz49
yt2VxzMnsNq0HSbBMZKCeW6i1x759qDfCQaXichF3DGDghtPnjJfh0DSE37Y/UDJ1Tl3EQP5VSfm
h7BkXwUwmjGS9ZdiyouOxfWSa4ak4jIc+ATNJVdljSvz/TRDesNlYyu46FMfwVrURhCrNwRjVQqJ
maJ/anYCfpeM+B/1LB147pgZE0xoo8DcGvbqgKVcPLpOjap1Ueel/yC/cI77kOVacYZ3YHw4Loy6
hmJCWmL4XmaKS76DvyFfSHSTC64E+WcEZ+8wTT0wS/Si4usrjSacZyy2raiytQ+OgYBXfwR15SLc
BAOaFR8vT4uNJRng4K2TiUkQOB0St0AuJ5dtnUG7c98yIWa1q0N2P5QdSVd+hAf15kuXOnc85RnY
0KZ9nzKj6JHNNZS6K0R/uWdxXHCLoIuEq2cQ7qe37f7/vVb72lMNWtGzU2SNSOwwDBoIVYHPg1V3
03mIPeqdWxjdDXgmKFLiPme6cqh/bN6nKI9TbzHGivZVdjzJfCPG3KVneziYaARodNWXl2+qrMCe
6ndXscNKgwVPzNT9GSKCiUYjLv9aa0KnDNHkxYHKt/qqzXJDF5YugxeKwHbYjYndbuVzH0zBjMZQ
iBc+43V56ICQg4m+FLn5RqHB7tKYLZN3fXV22x+lJSr836T88yeTu2XYikdkhAmjL8yxx+RYE94Y
LAPjEOCCMZDMT0ovCTNwubrFejekw7zy+SgzZjEFDsHLhWFmo5eZihk0X9CQZIRElbDkz9geXmw1
ikQOFiW3fDKMY0qR9t2iOodPcH3k8vbJW4n4tGvGwsiPhGWRhcSK0PYT3UXArl6xpE13nVGX7iaX
4wh+BR9pi6Kca7w3Pymz4hPXCotMYJVvfiX5dp8N8e94WbXlAZ9h7cXYEqZDlEP66Qu4+0Gtm8om
qUbH+lN1dITtt8WbMqzoPuWlc0cBV3iUF2CKxSfbP2XMas4LPdA4V5dvE32ePpQzB1exe+rTXMyV
5ALwfAzQbVcqCvQ18IdrHECcOSJi4rGCBowwZ/mDUN5wMF3vcfLuxA+wGDEjEvFVgFA+FYfhcRCg
Ti+dwsGbBaxIkpF29XPHhvmqSqBiDaWW/oU0HRtEVppIkoybeyhG6uoNmvXnax0hNcYHEiww/QPi
IC96w5wbVHuVeIV8m3KPUFZpTl+uTq9NvAD5a8OQxxEwhVIrSmZlnYdC0sCf6LJ0gN1UEM12zmXf
isR07lGkcLi64bWfVixXPaZvEk6Oro5hq5UL6nKL+EtlyJlRXOL8S7RvojZIc4geGCTJbNdGSFR4
+WKfAJGUQn8nxKDC2cdA6bYROr5CA6x7PD1PEn6IIVc2soWZQuhockK1yC2CeHSH5MsYn7p6fjRF
oYXCnOlFDhNaFTT7iWVJ9OtWmcLDlAr1z1RVpoq9qQIxtIU3aHYQe37ph0CU2u9VSkydKPzLyy6s
gpEgoKs+quvWcjeIIJUbb9/7O/pvKNcILfKVUouML380izs90QYbDLcllcZFlezQaKf37dN68jQw
qDthuJRanUNM6GBYLPzaZ94KWcNdKsjb+buuxPEhghZlAmXBeoSpdXOCwnWn0UukKmDC3Db2Sj7p
Y1JhkoiqrSVyMheTfG68iVlcRJ1oCukacVG/+IQWy0Dx0uUGAcNWNQPWB/ZpXcFGJRaGeGilOmZx
kg0Ob9Gjz1zwBNPGjt7VlolYwdpWC+QWIrbCzuSdB5HRXcNbOwnlOoKdkhGz9Q1QeT3a8zS0djxs
UU/k5B6avThspDJnWlAP+QeR5qpdoGJh9nKCje6QV/lb6iSshsIeh1effTh3cQfme7Gdr5UgdOgY
0oFjH5oz0l8gd5HfdYtUsnVJ20llPUiwBmQ9y92JvkAoikYdes/X87aWjOqGiBlEPzYhdtBNaPWO
IS0KWPff5pmSTyuaGSuX+tPrjgqGbzl4CdQ2syXE5VGzT1bBlyxjBjwPenfkGKZI/w4J3IKHABwg
XxKs84gQ/p1QvVy2zeoPPZOqojz8XJ6iLMuvlDn3XsF/FvkACXVbP7r9Ou/X4zGANRLrAHus17Al
TY0Su8gFUyOpY1q1o+1TaHHGm331X1/yYCTNvLcrVIiisaOqTOkEkBR0zxWyexcj3ue+yXFRA/pD
MIFcpyHpCkpzU4inQ6jBQn12bAQlBZN3Cjz5YZdjZRIMpu0PP1WDFKuVbz6PJ12x8se3sfEQZ7+7
8i57rZn4ILdEUEi5lr8b7HfdaoRZwB/xWVdxPIkifNguef2UqNsN9dYLc/8JhH8LJJFLcqYOqVK7
2ClBSsyFYsrfkqe9GXuF7hdXIzK7n1LY9XMVH7p7m1WIG5Gx3fyKuwiCn8tPnDkbI3vlVycgTsR9
dq/Gadx0EKRKnincQLSX7ahPnT3KrWX9kQL4/nem14ML+pikb983CZ5jqBSfGn+y/gGaycx6kIuQ
MK/cd0PMQk7quLyI1XqCm4uE88p3RFi85LvHbfhk0U5mLQxJO3XZYKNKdCcdwrxNHLUucPaRTobl
IW5YfBk6TH2kR8eS04N5RDJZDeEza1j3Porll9SxRMuDbpRF1zFVMdr5UYxZj+XQmGKdd84EuSo1
d75jnu4KQQQZ2atoeZPMl7eLil1C8kfyHMjLta5tt39pituyKX/gwedvBi1lgAFqNbzi9Te4noBm
DtBRo5DdPgWZZAwFLqr1tm7dNVS/lFGOoPnFvdcfyxhlaJ/GLYZwXpTwWWqnYBDbGenLGG53fn9z
2dReN6n9PgRCwcbQIYvz9laU2zN7AmKnDt2100nfTfXV5BruTM9jnKLyfezt0asSgqjcKx6oPky3
hUDREzsmYGSQLtj53w0MPS9kymN9Y47O/ftXzztwi9poNC20bT+eCfNvT1z1eKkDIAqKIGgkbI14
6EPb57Mxll13uvH2zepyQ0RHH3WSbivpGLO3plhh0xsPPnyby1wZktcsARmkFG9jyjRRRlg0VFAW
Oc4K3H+EIGCvD0p3tNCYfA093oddlWlpQjVMXL9gsOLuQhfTzgon55ariHAvM+1ogs0lEywx37gM
1nrUUa+aAGr8PIyYAcM91ST1YpM/mK40gO/f1U5AA4hOjL5/Pf3Jl6Q/Bus67NPrtKLjnhY5Dhzw
RWdJsm8KNrN9EL5f7Jn1dkgwV2T3gpyEsJzRKIsYAgqddpm1zJBYN29Ng4cp3nJJZPT9wH+GjwO1
k86HBVNhHLegNE+uswpOCMbLkUhzgSNuPsHOB6BQi3MxdTGOTcD1OFkuIU8Jvzyub4FPvPHg0LaA
PryJyjWdexMJHTenTDkl3AAOANR/YTtBo8P4X1hA2WA3XQaC1SGhX2Q7HV0s4+V0oQZuCNj/3AoM
kxGAH4UpaRstayuEfg3jr/zrK/RcIF1mArnAJAduRLXgYV0SJVnYVCXBAhhM94vaQsjRpcCmlt8I
lgJEQdJ2c+yxJPwJeHdQEh3EtsnFDRF8W841XRVPznpq3c42Tgca0VAx7tR5j8nmD98yMkohU2ZZ
nfr+nEt+uo7h741+BUH5RdS64OqoGzslNFAhmfl9Lhi2S2qRosBMPpAM7G8+EbJiQwj1SIu8yYnv
GgPQExlhmNNkSvlREui1WB0gFaV4Y0viA++MO3hkXMtsY8Qxby/J6LNPcPMSUYCAa4HFnzmm7Wbf
k/NaSaq7E4AKlu3BgGBnabyaEyiBdHSmiTw0rXD5Nxm+k9oYRB+Rr/okI7j/qGOKoJVvpaoNm6X9
kov5r0rIU2Uvq5V0KslVrPMTYr0estn0lK1mwyyh1cqBADepRDx1bZu6IIsDSA1I09Xrq8T3LFfu
qmfD9xzxLN9NoRAamRCnA/ld5qcNz3QMdqGgnN/yZ6RjQGoi3DOF/rNDFAjxabr4APWZGzlWCJWq
EeQCuvLw9GGb2aHnZ7+TPvpi2Th+Rpek67CtajW5NdIC6B+tuMkOlQGGM8y/wopP+Sizpn46NyYT
qJ4sdYwlwGBnqJuJPKRIG68F5pewZFlxmPuCKN+NPiv+LOY8QeswTeO6j5fxC0++J/Axet/XeJcA
WCuZjf0SOYloTqWsVgrNWmWeWK52YBOfuSEg1yQ7JUU8veREaPla4jEWlLh9yCPGPpDgNYb8kSKa
lhXQun3xi7WHRLRJtAOmLcFGrarvi45Zz45jaPUAOnY7W+v6YdA24uxyefIlTPPvX1qDHT/zQ+Xa
YtvGZvPskhCrrsPSoyruYyOQB4MQWMowYhdybSAVyyYSHs61xMOnHGmVQGGHulH8z2Y7YPs8soqs
9IjS4rCXgdMnGsyrpem8FSpAy5yIaMu9bitFRg4DbKa9FCCnbf7Q08kSsdFLpL6TEm8fS1J/RCPk
f8diI2PXFMAzSv2BuOw1SGcYCUpj32xKyf9rQpOTMTdeQTf3tClk5BNj1u+xjQahROtYJzZ0LbiZ
WHy1kC3Ftbuw+AZUStpSrqErcKwc9XIUP/VWRk6LIrNTU7Ks4zSQAqZOu4devtnX5SI3wd/qkDxo
QAHG8TqO5j4YFPVm/XBVXW302pR/HciNQ3D66vLJwz8XtWltTkR7EO0u17Kxr2sVDP2OmIHKmNQm
fAhyx0+nLv+BdRhuOczIFLd6t1V6WEx9FJ/lQ5SKJc7EJUq9QgVHpGsYd+rB99/uXVcsxvqB1CpX
ptdVbcpQSverojbeHtATGlLvtLkg+QzfeLz48VZNFTskKsxJyhfnKxU8AHitV59lDiOhxld+Llkv
kwMthPN7f155kosRoQsaugICjUNJJGK40W/Vh9a3jewXsev5vRbJSSVGXp79IPL1+Hq6MOfNFumR
kE0OkPymv/EJNgyAg6eZABS0OIKCevWJ8xyK6ziaeGR+yYyQIU6KflZtHgY6MAEFcKv1I+hsvl/C
uR+5FG5lX67V0S2WrNlbIvM6p8WCr6dWG8KQ4UTXXhLTW7WaGME+J7YRruOYCAigkeGfP4r68MpL
nJuflS+KJYt4imk+ltgEV2PHOuiYOYAtPHylGUQKUza4hy15dzvAXuqCsZkqlO72SemS9j9LZ4BZ
1NMBHrygTo6EZcnOwDOHHqOlhDMdil8bgVQ+glEjw/gwpXbBlQJ8LLBVmg3h6hDVmMLbBGpp/xSt
QPQ59aqK1c5z2hVIQFh2weC9ntMuxj+tK33T2Q66JLeOROZOGxwHsx1H9KTQEBvv7aAz/TrxyuUm
Li5Z0vI+AB+b4IBspO7GzmEuMz0g/54mkuyrwKhQtVVTK0SbZQmUaBXhOxfNGgBop/CWRpVqPZuE
WAlmrlFVnAUhMd/BW7lrloytpp4Z+72KvYfigoeLQq2kIZORAKG9o3AwiqaUKvopoedtdbz5tA1q
X5ooL+e2kfd5J4Svl1ylipqR5Ky+YTSsB3398UObotGoACJbbRC43HDQHQkhdh4INuMgNOdnPFmB
bWExXbagxfIXR+zNuTJbEq9WquAHUdQohyrI06OCLSi6Nhtx1fWK1lyehZZHGijaYItpkL4o/PS2
A/88dzvrkMiJ/GgWbnToAht/gouZE5+V8aih5TZDO2kzh4QAJzWUa+Wlgk9WYMezcyXIP+4tuPlT
EE+o3/it7nql904liycbkzCI73uy8s+oxJ+ER+MGF0dWZNngcthHyrvAbs7BLJMKBDwn1pKW7X0+
XP1wcXcl0ntJxhc2uKZcx2DebaudV9XqGcMvhfcSpY3lJ6UaE3m78ijVsvzx+GEuZcM8ZvPGSuOJ
T3Wm2Kin5FeVX9BvV3vVsZBrpl1eU5Dfr4cEftC+Hs1ZW3nL4pzvUzsdr7pNrAtiUvhPXHphvCIX
NT3R/uBHZCpQpjr4Tr7jzkOg1lPeiaCO9YyACb00vfRUssQWXizl3Y7iXI8fivfmnReyW5wAOoQN
ztbUvpPfaLk/QAdIcj5kb9EWELiCxMfC6dEwOFlOkTOEs/iSMxJ5NjTShlgpFnXztVA0cJV4rZqV
X/5n+TdJl1XsZysV/4kGspA2Z1vutIZeqMG0FawPjMrjAPjeKgzJGj0iQgQcUu1fUpgaLwqx1XSp
T5O/XQrw9Ydn/HrSNNEGBugODNLKc/OaeycV6g+NWSFzO80xX9IxdoEAbjKsrHiae5vTy022fleK
gJT6N2zEqXnByvpgC6dZGlHnuOOxM/Hzc/xS/oDnlUD/pLv+mjB7OJtY8lIfLb8i8HFNETvFCeQ/
zTxZo+6ULCS+Fu2Q/IqXYi8Jsq03gK4O3IOOXzWEUbO8Sl3TRR/UntUzJdESmeqBhai8+2286SYZ
A5czZJXTO3ZlBs5grmacij14YR1nNefvOJB0UzZ2Ocllpql3zrT/CLWrBG1NJ9m2C2/9KWLwu5NQ
fMV37h0F/PQ/cmWf5zvQHpwm2Nk4BCwNA7T6UiQZz7TrJ0PW646DY4BQZj8T+DocwHtE0+c8vByA
oJGqG5z8RsRNDBch8c11pSpY96gpqj3EvZP4NsL7iFK5wMCUSwqkH4f/66e7/ugP/D8mKzGYKz8/
w5UwlxSxGQDTLBMIAB3eZyW05ruLhfajyfCHzXWF1yR04OKXSroKbfQA7P69bznsS4DWQ+EfnAzC
FwOukoQh+bO2J0KbuszhZzrTtwGrm1E/8fHH3jTe9VTJUwhZFrFycbLYOakK5F8I9Y8PiYbr2poo
XW0QKUV4XHtWMDaNLmxJZ8SkOB+A+FbwpGrBr5jHbgvvE1T16rtp4OXxtanO0zsMWm6HcutB5est
XW6QvyCwtFHm/1XIdZ/o9LQYk9yqqxczVwGgqX78cgtGGNFGT4gZV9fR00N4Opo2JxYnRxsacHN2
pNaGY0fNJg4cOMs6lIN1hLj5T3Rg+vggjAkoUpHimSKKfhdG/R2siaYnOyW7IjtEHm8l7PeTMlFu
QcQZy1vGbAO2xL/90ICRsKXn2XZbRz3eFDkzyoflowdoxTYUm4TOPDSB7XofMs29urkRyQWZcBB4
qcTcdsR94YG2st/Z/8Fa3L+QzZFaZA414v+4neCQiCI59dCVzx2K5UIQ/LjhcxZ+yuyG+Yml0Bf5
Ls46lTPGQSRik/OcpAsikFAHJvACQn0Klvu0ddD2ySYqx71PA6mYUxxid5a0fWuwM8qfx3wayXrz
JwxIVtIf5D7IXDsn8NY/aY96FPTAjJPdUeMRhaT+DbtBNZvMP/r7RTBrBM+g0LDakxdLF5P+Ja+f
tsQcUAuszX1TmNiI1rDrWIguvdBduWmb/lqLnRoHCbHHRQuAyyhrWLNJ7+0K3DNI69dpCBEp53Ba
6C3vhgYXoakab2kOUCSyPSJawPSQ5I60fXPGx6Cg95XqdIuJDozmdBSOJoHHQZqt3xAyJTCRqb2V
cTSUuhLFZlddjbhYIb5t1wA+olU1S/VPKyTVyuJLdHVJ4LdCE7X3tBp4bM7ez+KRtP7cfjPGzAYn
TTWiWYtxemhKeqUt2DFnWQUBdVDJWJD6hKoQm3wvQeJ+NXQpYnUzZN9AbpOFLLm8HMOdCbYHzpTG
nFMAynG4gCjpc16OELCb0vzwvXwUcTpVp8Ym/SDtXc/f5xwgOg+pdIKJoJWvUtIpBkFCcmwAWOoC
V7LsN/Jgk/fqhSbKTuiPf6buk/faJsy/RvV0BglNigDZmuIMnPk/FSvfLtBjUtJav/iATuZa8FBm
PVGmxa0vggfPR8+fzB8+crb8Dj9aWsS4aDDmX7ajjEKvvrwLssd1EIh0EASnuQkx7NiNXpsr87a+
oJqfZjj4GAz7mia//QiDImhn6LgwxgDGS6jLdNVnUWMoPwIPxcLS8d+OrR5rfZvqhMsJwTyLkVLH
WAS3ZuKO6Sj99zSngyic6ULylei92DgfYXQC/fOAxQKwaXFrNCCuvnMN7kouBfh/0CpnHiOCozTD
GxZfLcE4r2Q2xu+P79hJAimig0cbE86al0PfVaEsN9A6GBN+84CQUxd+P7pC85hkIflGlhvKUkWB
C3il2Kdev2ktP8bY69OfvLuYn+/MvZwkc3sF9/Wn9yipW/bR6lzaMd8WXgz96rvptV+P1Wris6M/
kC9f1Vdo5XpQV/rn6yG52MmUGTMs4ulPG/CuIII4vRQ6T5n/LiKrwpBjapTlMXV4xOTDV2mCYofP
E62FrQsMgV7azYEz4Y8co+8/ATZqHOXcrgTNTaBJNmUabm9E54yuWztuYUOhujy7siSDm0emsAnE
ANgjZWZeCfw7adstT4iB6++bYXy6P2AcAe1TOM4UXqYYljchUB2XhHMZy5zwezmjuz+Ato8WSCHs
QIzYptKnvMIKf0dGuId40nASH5io6hL+0LLS4BX4lFX999YsO/1cfpmdPhRNQfJ0sbKItxqvZvYe
ViPowoK07fpiI3M4OPL9JcAYd/TXMi3V7z65cnv+MjozdSum4VcuvIvyKIjnESjwjUXXs8N5UN6p
Ce6DL5WavyC+oD/i4Ok1Fd3PEII+iM7Cj/NhRA4UEu6oFzE0K3Rjk55iouXNyxVRQphrZymWkEy5
KgX22Pcy9MDYFZ3hQgkNyYwfiPYC2BMy4qmaFKJhkps7+/KT/DB62+oVkA7BPjfjDbbxSWSR7469
F8WGaCanrZBQaYpdiMXDOn3xrAfgFzEqb/a+6srXWMsownVO8sRVTUQgug2ziEN2zDLhJ2US3yTe
LKnjTzSsms8IKSXNS0YFi0Rh7NvElQbJt0vSGgCr6fFm4YDio2mTUUUTOjbFbufTkQqhTJ9w8iHv
o5pR8wRbRWW6IGGKKAztQiu76u7eR+iOAn3syyFzn+YcmN7UmPNKZzbFOvY9ELTIbm8nE49pA8QN
2CY1i1T9uflVSBFqwkQPTtTFoVVKsNsYqzeUkacnhSqTy0fPQE+H8XLjQI1eF8fu4lEuWWjTUK9c
k1PRHU1zHTJGLQ3D2GQJ4/QzJqlcxesUmVzmqFopszBw780M4+Hd1aje46lXdbXIS05+ZfpyLMLx
KvHyCiCEa4gV7oufRLxkeGc5Usl0o6/7AErdzUQ/6pPzSyDVAAfsG5IIiHen/19oXpandHaybn9i
3FxX4lFm8TegowbqqsRQXGkXXQq00vIuzEWzz8x937Ap6InCq5vItVLPqretVLVew0WmsWFOsiDx
uBssvYx7h1NY0HE8rYUMuYuncyO52JMrIlTV4EuQlrepo2kZ0O3RgJQLrmR3HMpUn2PxBjV9IkiK
BzR4kfPr6J6WP0O4ogO3HDwLHnFP43BDK4j65/hWdGGeciN+QD9wBjMqb6iGsvurKOSI5nns3c4g
qKkluam07gfPaxVXDXQxbzsK2fNdDGvHb6l6r+2b0MGtbeb2P9U9o//4+wAASbb50OG5JRj2BBKT
FJ3nv4GjgpJwp1khCAOH+rmucmVBlWYSDQ+GZ5wGw5v04amWbUdXOqrdY5lgwxfxYA7kD6FKfPqe
2eXabpch3PORa2GSFKqaq1/olxTKUZwnGNRThy5XKjVSXXAZnHEIoMYiJcZI9XEwWe+ZfR9eFsDK
TDHuL1NjBVcM5SZe1V4CY180TbtW+TXg9zBlgMrYvqKIAHRmqn9d5+gMor/F1zOUFCtvSItV1uSp
sG1znVp7qLODIKj5tPeSaIyJC7y4cv605IfnMirpp42J/4xpOSW4ffxT40zHAVxjnv4qMmKeE8gJ
Lp/biVyu/ps1lSKGTJ4iM4oY4i6FyBQxtcEFkp0thtHyT1cE7IbPZAe9N8UyTWhhO1hl066+hziU
aGQuWpSSRDeaX5bNHp9hnhHRINlumNCcGewMP26IrtuXLUW/FacOTIkTchttgInIg4817ldhbg5e
X71Cggg8NzYQGEvHVkMIS3dmsbfIn9O7a7/3Dr0P5LMV0pasj42Z3gGhZ8v+ha+p0rGAZp/Z8deE
RBYabExWIcIVTSVg5PsyoqnVa1lv6EowKwjqr/xZMWijNEE7EEyaLp8yoVh7BJtPTvXtrUsH8c/Q
D+dKPD8xgIx38V0zzNdHVVlQEoEA+8D4A2Tmo9lyUn5zRvoIoPtu/40CSpGAVSmxHKVLb9l53TWx
IvQiqocYipaaEuK90je41q8VW/syPzPa2scwTKHKVHrEn1/145usy+ebpoulbDV1hA+W91KcWujC
U7Is+q0qRC3w8PdyS+avf/oM8s9FJodMG96FBV9t0hFcJIsNpg1+w6uLASjSzwMbzZJ1Krvisv3W
XGawOpQH7rRkFvsNURJ2qtb+l41TtPP70+CgG6n+UUhrf+4f5GsffTzdZxc1huX0IoA4BhZs3jl8
8j6lxvn1cJwDS4Q3SvHPAcTf0HrkZZQnpr6gs4cqntCTmz4RkV1rFVkHklW1tbbP7LORrVBT7Rgb
9Ka9/eJIUOytqJ1s6YE85iKzuug6+dMf9HD5cGCIxIoRH6IjE4za+s+6eRBj0gTOdQBM8bacxpdu
qQXyGWM9BTRQHsk3ZIuODLDFjqQjysmQQkWuTGIrGG+BddB6H9g1vdmhGGTKqLpEi4wy3YhcXwQT
jcvXDmrfY6pZKjYxNNHo1IkXTcs+1ldOkrvKkry/oqWCKiP0S8WnNXY23ABZvZuhTpxHKLVc41tw
z1azy4DTLLvIZ9DYhVIJvIq2mxbWM2Iznuj6WDo6YqUteHfiele8vKCYZaA/eN1ko41AfsDlu6bY
H6xX/7oVq2Rw3ylg74xOSqIhRWrTgP2//4NRPUaEhVwjkpiiRR6dVVcAL8AYbt4glJPcnYTauF4S
rt2yO3/cxrZChcWgqu7f9x+o87FH50//+oFy1VCcpGaao7wpRCoWVkKMrd5r0ArLgtgcu0UB9XJ9
iUm860XNud4tcv0qaSDiZdOYO06LGtWhHh4m8VN1a1XGYs1Ab6Yhc7IF6E+6E7uqPauPR2IycSNc
iR1Ffbp3Qo1a/eMNlf2N1nPN8mKFkDcJY1XN11ln7DGjPdEmm7UOVEhlJYMslZsCFKFHOmX5owPf
VfQw9i681AH4Xc4l81pxdQ0IDWQ/1QtrYcKoZyyJim8QFyA2Y5g34V2nj0GoKp6kjtFTPGUe6fyo
gU+5WBKiM+xanTv2RsI7QZkWwzAB5l9XUdYNqzyspKvw38gzOMjr05dEhrLN++LTmSpCO2NHe6M2
CR5ADoi/CfWaW1iOGlUdoAxHGRX6xKaFxUeBScqeSM3FDGsnRdGSUftQkWFUaeimDoEYoRnVbM4V
k4rRH4j64cNfHdhtRBFWm+qpLnVgGTWAwdRwBz3zFOEC+xdpmfQUSeEMQsSLSQ8XEb/StXXKiIl5
MbIxLqIaNGqkOWo3PBVn1By5B3ZSMDXj1JmfZsp2R9s6JWLGg+ymmqbco2TWOzGD+i9077XNuW3P
Ek3VLkbO2uzh2Iz8DL8+RQ7J72ES1g/ru2PWssUctD1DefZqHdz2fOgosv3UIFJOeeIvbetVDvaJ
vEngt4MT6qtEcWppwhn4a2ePZuPI50nmwacyXlSUlA1vjTXUYYZEuQwPmwHf4bl5NRPwj94Ds639
y9KlE7q5FL4gfO+8UT8bmD5Q8geW5hzRvqWz6BwyntFgt9a1BNl8v099jicfbc3Zxn0wrHaRYXPN
q+fvYKERxTkMF/P5SzMEvt4nrtB5t7wKuojhGG2jJVrY6O8Rk120Qw3i+NOb5ZlKpdbORcAM4ZZO
CLS+c9OHy5mjJ9u6WbP81RllVyYtj22D6Tub/kDx/T/m1+yScYIq14YNXA39gTyBtIy2YUTy6+m0
xGrHS5bkp2HLGWCqyra55nnGEP0xdp/E1fc6aKnh+a/K349WufI2gN1g+FeUmpJjFWmmLf+Zmy46
Tuu3Ph4QHKjjrRkwqh+uKQ/qZUjGyXqiYjQQTJtpP8UUbI+Jt124bVEkveVZSzNR9DGP8GX2Wyfm
AAQ9IJE216whc9y6+aL156YS5QuBbfluY27aW+gut5ElxHZsMvRwfvPD3tE2+/kpuNNDMbzplNZO
3AXI1ZQdWm4qdWb3bUkJBeseVe26BcPjkdgzCv5hCkW15e4p2hJ+noZjFnmM3ZtDGsZFD8mmF+FV
qSEdapi2Bu2Rdw/cHFNp3Nsb2WY6v2qAdf9f+wfLO/oj1Fa7OEImJWJ6poIMiqcNuipp9ZAk6+P8
MDTU/K5GLsS/i9Ky9aRZ1DD1WqmMd0TUCUIs8UIWPHhhmrkRCGr4McN2oXeKsq509GBQW1i7mtxv
sojjVXctF7gQweD7Akxn1ycCKPiJFH8TuGPA8AecatUAXCxS2c3SkxufInfty9C/K0i07DrhvG5A
abluBMswWq1eg89tVZO8vmoOaD/kE16GxCCMcqRpPv/WD9YWK7drqibLZtDYb8xVrGDgtqDU0XCI
EZYCTktlnxFcqc7ao/rdM/S29i7fbvugWI0iRzL0Ypqh7IGHKEVLEIx+i62bxspZsP6uohJYCPQj
V9cmNC9R2TpNpzItR9rWEhq2BUPZNi08qyLipbrnKGWgPh+hulU9sLFU7VDsbDaf1Qy80coz+Sho
vUSlrZbD9O8azjrsMO97SgtcM8fZnUBMO2ul7stV4m7dMKEtqr5wRFh4JthtfmVj7c1OGIUjxTcg
G4GOMSLic3WeNg1gZjeSEu/g3FgyMerOrn9Ohr3PTPxCpEQtoMqduAM33h0jklX2Z0FWMAI7Kcvc
qHRjCygoa1MJZprX7XG+9Bbr7lg3NrZkW9qT5bAJQTJ2qsVOLJ98I2YUhdm8JgsThtwbbPagsvcK
DimglWy+R1kcv7roCcxd91vffdtepHVwAPWG+/McJEaXtRj5iTG4617BuO2AFfMlaDEC3Npl9ozZ
lYfqpwbI+mrlUoKPg/Qk5PJazeE/fd1Yf2O66Gvi62SPGITBYx+Hj0OwjgsG98b8QYSXTUfa2/Fb
gGpyGT9xoCPHCqXCeJuIOLJQPbsGetHWqX5rF4AXca94awfU3pUWM4/4tTxXD8c+oaMQVSiJR70/
0hQpTJ9x75nnF2gNtWwb6274AsUOtw6rtdPjcbXNyjmDcj4NaySzbt8NZ80yikHTkEZS+EuJ340x
96krguF8C+l4cc4rt7Ye+/kq+tkg/dBAJTme2rNYekCm7uNupNZJpTRyp8RZWrhoZYNM0ZsfBeAn
JGptoJGBLKCfHlztb2vnwENaHOshpzuxYRc/7pRHCzoDNXRezMubCoo8Ny4zYZrqC4IXa1GomaJU
cLZzaULRVuLM8kLBj2KJYBVeQgLKCbNN1ewrPMDSwcTDVGo9QRNiV7OhYRZnZd8vgUTX1gdKWfb3
xsucN2dDuMAxRk2VtsZVLrPJDouHiEFtkEeRjtcZ41oodq5DZVNx1JEmXf0A8MrYFOPmzuoeOyBj
CdnQCov/is3a0l/NoMgLsXswEUVTg1WC09nnpeUC6A5WmjqisZpmKnhG4Ci9bwp0PS0TQpAWd0zj
Xett/WZ1lqvH8Jydat7lFKeDmNZfx+z1QaQS/90hb20W4ojh3k24BuCdcOUzuPHaI0etFOnkJ+4S
JKmvD5wfooCY2YySnhGAAKCvnARdWf5sCjysM2YubYLWEoklZPWVidx9Wo2V9T81r7BHX1jxGeJG
toOrNHuuArfYJ+SrBfDDkkPy5GZsWFlJNRqM/6F+MFWvP9hQPKTaOt0k0Q+KnH+b/NK3gsp8cjav
2LnoUod49qqYAjlFSbzZHTJV4XBPutdT5i+vWBBIjh/vxNv/xrM3iI+7ln4Ga5j4zKuwU/yLzEhs
SfivHv3QzKukOJm8KKafdd1lU36XmInVlkYKNO/3Si2T1FLiLpxr3ifz71gSSYoIxuHezOOnQVic
DMHlu96IEOkS8pt3BM0aSbyAgvKeXXSF1RabLGhOKZV0vbEKC6Q6ReguVQuRB1gQIf03wHWN0kJ8
+axKWN65eGeUFShGevycE8vKazNv4tmAFryUd3G30FGMH6BOqpsJMNRhEd1Ixf1M9nXv55649imm
kdm9nCoj6lp2btw5+pmPkn1XNuz0tLqCI6XAL6K5iNsvggq/067JCDweCMnv/Xlu3L1iicceuLzr
BOP7fjGaKs6eUx7TP467WSGYPe7KX+tyZtLAvOcrJyZ1YbFa7rS276BZMdNXfyHEVwC85mJfua9J
/0Rq+C7qOW+qPi6EZM4fJxBVI3wSlj5wMafLHxgivpv2EZAmjwlv1hGBuKR05LYXldtdmn6tpwCV
RDpGCVB6A7Ng95j8ia6/dLVa5LqXoJKnSTQlYwtrZHaP/P/h7EuLDfDNKACrn1w4Cihg02+ulZXz
cn9Ez0RtZ4WIB24mdvVnB2ROcU0d2dG+3WCxunDLVlRONRLX0P62ZOoia5diik47jFqzD+4GjA+E
cJmwfqwg2MlHBpYXUvnKD0Z7FuPLMM+ZcC8IiZPc92zO+tRb10tyK/2aDm1JHLv3UCHv7E923DLo
X0TDWT25nP04B684J7J5ibh8cDDDE+OhGKNk5AYbAyAGMD6G7wz7meCaY4I4HiisfrTYq/Qz1j1h
md9Y4YAchWW7qlT4aoVyiKUcYLJdBmVuEzmtMgN4i6+WdUZ9dk+fdLsmDPSX8wF4lcpAPr3ySsfz
B9/TbbRCkzoIYSGFd8E6+lXIG/qhXByXEWlcN/qgWveNe92Pi1VdgZT8WKt5OqWhwqL2JxJjURva
vqAKTy+gJeiGG1ByHbh9dBGc2AYSIg6gbOXHLXUYEYDcnM0COpEmxJFG8zSRqTxqR6tdjzGw7fyf
o3DzKGpwnpzuHo+BZAfWnlsb2Ln7u4Ie5H4Jjt8pvW2mBtASKTWeZfnT+9AgY85/q3lrD4UqygtZ
VjGvypmeQATqmXiHkzVgkdecfo1Pbn8/qQSOSx8bTOu9TbmhJDI4j/3SvWhfiNfLfcrKJY+UlJuU
LuGxV6dv+1OnZIF18mCOuV9vnYN5GUeNkYSATNiZ2mrVteJm0c1nem8vfgJj7T2I6Z5tSX3Nbbhy
hZkdLD4xhtUYrxcGDSJ5x8BvCpW1k+kJJ4COLSpzn5lycwltdF6KXk44qNQlMe61AdnofJDCONX2
PV/bsn1LMFx8XENr3coJ9dxXlwQXx7mjp84NcBZ7eFVB9ASa31dtrtTC0/0ZfTDcn07A1qYU92Y8
RQWxUUACYhC/jvcQBLb3CzFPyi1rjwLAWrVJhHWVgmhHqA0NsOqZVFEoZzuomNFG2vstcv5I1aEg
ezIMnJUKbRT+5YLYydpNFArEVZ91fzXIrstwYBx+VSd7aPRmwwH9ejJ4LjOtxzlc+8stI1Kkye8L
SnO2U/wwJR6cfp6tJNRRjIdyD1A3SDiam0EgSo2te1a8dQbALKLV0A83SC7WGoV471SAj9EWBOCV
TA2d/gDMZOzLlo4MmddFVHfRZFDgte/p++dVw5Cfhc1mxrU9XxZqmhUCoRr/0bilcAlvux92fso0
LzNwr5gZweNSi7uI1Di9w8qW+9qrVEb0ljX9MQXO7Lv05IVBGsqRwSfq4x3koqEg4MRlx1Rku5bO
TVFe3Tf3gYwlYV40i7ksvPoD14VA28F3u7ArkEdpYaSaLyUnp9ftRKQReqi8PDwGGQwyo4ndaGue
FqoPF/nEcl1AvqaYHcRTbgEGVz3KqcXCOA7dLZAHe946aSzT5gglCeZnjMAYSgj5coVGGfa5buYD
XqHURL+Fd79gsjaXMZKkDvunYi/JqWU574NF4gT2R7o0zRN+8aqGRjzc5L8Da5ZEEJFZDxjul/Y+
qHvb97fkFAtuX9YqfZxMgYj6QRYTsx687IGvV+Kp/IVQrr3ygqTxx3fbX4PCiaXkTaa1ZFPYHbWO
A+lHqxDCCAcZZXaPjR0KCYtoGvCRzgmQkFtzD4rUG5GfBk3pCU7dflmQgba2AxouxhZuCZaK4I9B
RNypLlYvaNYzn6g9DbfzzB7njz6ahG6wNe1NfPALNY8aEtkZM6jG7Ik96OtdgdXLS1jIoq63Bc+u
T8d6dPVKY6sPU0gOwZtRRsy8u2PfuVQ9tQpBC458ZGfODHBhoP2OolDD6c3le49hpI3FwaalBOJI
XeJmcTskK5reMp0UFbI1OZ9z0hJedtBKNMMOCT58GUfYevi9q5UO3etuzHxuEPKceDOctiJZD73N
gi9wVmSZhlv6m+3oN0dgXI7+WG4zyE5n47ClVs+De2nvkDNn6Wa7ovj8hzKxdM+BiY+nnfh/buJh
9/6gg7cPSWmghKIlAekLQjKUJpUmXQ1zAzARn+PHt3IfF1Xo7YaoAL4HSI54IR6JzS7bftPW3aTJ
AIvsNbZU1HURkJ/W3mQhohfO31QQ3mFR76BrTq74iWlLrOG/tcomDAwSPdeFMWou3U5IyG7g3WHe
mm3wYrYxa0dJvn7I9nxl0hhh+5Wp9EYQZNf3cEFpGSzN22Sb7oavhyvKFtWUFlJmIPvN1hdUHo0n
CylNLarfMxLwakj1uxECNaxyxTtXotS/7ZCC006FRSQPM4q1JHf1fDmSaWsNv+HH7ziRvkIC+pla
mb5hUpyOf5lY7rqMZp1NEoAX0MnF31/P3HDeVamJjyT4e6wXQHiwoDU9/oIYD+9NJA/ZWaGkBWU+
1ej/Zp/RHYPVLMJbom0mLGl3ilnJ6ypkbi1DeGXoP42YTdCR7+KYDY7EUY7xZz+D56rPOpAM8wpR
onAVlUWqku0GmZC+8RshxpbD24tkZL8PaTXJkEPsoZfOFZstqqmeyFISY+nu1n1UZNFNs0G8ncXp
BE/+u9W1UDAgBDuPro9txL5R5V/QGx6kK0/Jr1LQ59G526IP204jzPVcuZFGPbODyngpshYMnL1p
gnGE/5ufu2mIWoIV5dUIdJFjAmZcBU345TkNkzEBIjzGMchUXLFdAM5/vRKKDxXwERF4fqlvVIP6
ow/9966lsH50lchpe/Qr8igmes7TdtCXZ2J26XVc6TKepOppm42dVv0oZ0scpTqxLnasq6+QjwDg
ywb4WR/hmkw6WLu6aeFw0KD2IQRWY5CExUiDoHr+cQGSk+eV9yW4lW/GBboXkbFBYVXTlWDeGWGx
mTdVpZ7PrL/QHydjZkqBENAmz5/9W2z4ynFOfqq9gGgU4XeutDoKztWwMOkDHSTWWamCKCqhq0uQ
5QsxzMG2dfYrhYflkZ29xNdaiZE3f09AU0HyQOeS/2Ht0MrtsjniuSVKNE+q/e3MqcGiCCGDqwuE
ewNFBk7N9s4kV5lps7KlqFcKPH+V/8THr95l6prG5+lrr3zJQX2hNF+jnPextQBpZliOEvRHmrIx
nui7HcBhMfCptvB2jkP+2wkp8r5lNENnwXAp32QMRJjxtxJkgEaqFwi1sTKUqfKEu9Ykoy7dkSH+
/foIW8ZT7jwIMUdmwdWXpShIqHMdEDPC3V9OG1rO49aYqt1G/z+Jv1Xl2d0Y2Mv1mgpfOIlrqlM0
+4k1TYShPruMzYPhVsK4wyfthXAI4XFHlzQmWXyWbEfZZWvP//bDSDrQJwi8nuvsOzd8Q9n+Ntsq
zqgnIpA7CiEGCF/p3+Id8awjR5Cc+ts9Yxcp3FtApSux7hKnAEDqsn5UHdNHBqDn71ypVvN5/cfb
KLm4t4gYZJVvZDrifefr1j+GfB6ca1aptcpuHEAaBIK1ILoHWwwFqNaRd/ysvLzRpSztQ6+AJlCK
oWosf1270bGrUWfBhQJeqHCY/3Tixdl7OrNd77asP0Ho1lwyzejqz/uIwnXAhK48R1yyNVV4WhCm
nDn5FhTI9oGuoap+Dhhu2aiw6qAfcgLQ5fLWE8WDPmMep31eGpd+47Dn9h4kGaRQbl6OgicF4Hx9
ymDAzowd9ERaYKzmuLKsP4rl2ub9ii+eTHNXJTJIHNOXXzi8lSMSuuCYBZjwR6JRst6G/Eomecp/
JQCG03Lq7zN/qK5NJCbAJsQdsANUB3xZns2OkR5xW4E/Qz1m+oTC/MEGvJYn111k0WlUwNcKdecz
KvO+3Ej8tN/bx8kSQzPgojZMhvd0FG6DZMJ22OQmy0crlart75PpdxpKdyVht4+FB2fiJXrnCmAi
yN1qu1cg/NsCK17LhRCLKjvl9WdSxNOw4/zrchJuR0QYpUeCB4/9YtyqogZKLfUT9k75a+g6/yHn
NetQ3Ldhtg6m3IFAnBcfLFwKIOH7M9n3drPS1aJ1A44Kd7McdUjzTEqNRkMFU0iXGVjkW0thn1lo
h5jygq6DLxruGI/burzCAK9VF4EL/HRIrfWfr9/MMfYzG01e5P118y6cAsru9UEbx3f3/YRlTiS0
yGaiiZUEO5xEv91JWI4JSCU0dR9PXnlcCgZSc/Hl69JfZJA72crLmH4LXrWTK+/KKcKNJqeKd7aY
xkTgL3fEiBvmutM0oVGc30m1J4+vjhiGD4IOyF9XHm1Kq6E133SO8b8dPwtT8+zeqRzjZZrq1I0f
jKvTwJN2ppO5y5Mh34gMw4oeyWqhq6bChaUBMhrX4qIUUJUcTlCl1/e63JCn/8YCYa3H9xekUV1M
tLY7Tv8BaLHfSwf9q1BykBqK4MJA9/lWgckAASP00D6h4GYrRvphHpKbqcUCJXoqqcmWkflZ1kb6
rrc6XkuzI/jHl4KfO2knmjB4KfAcs4Wv/opn/t+wQBKDIeNN9mFRCf6oT7sjYN8tsYdybpieNJQp
ip2Wzjm27RWLmrz2l9lb//dg3zmUKTi5Vw5qAzoB1hdziXF7wBhZReLwABAFiumFOPlVAjvnkWZy
qIRzW8YhOzzkiKsXzFoS+6AEmVzV74g58kPIqPpAkxfI20cA/OXP+7EpMgKSkGGruPopDaYJagcm
NVGvHL6sSPwQVwcmze/JNNFghgD3UXqCOZr31CYOH8Ge+w5VtgBWvZ86+BYetNUJ551f57gHfw+M
5roIMERrfmy9MhzBUNvfzi6jQPfH08AIdQasrmGm8mE6hoYMADd/EVLHO9UvcbNCwJUFVvhKSYoM
r7vDNorJsp4juJ1CkF1mDxHkM/gJjteeiBKV0Kv9AY/B05kjL1EWzbADMIhllyjIoGAISum39D7Q
DXBR1fi0SFzto8zbsk+YJqBSpMarJpgc6Q8KPApv++V7O8GmrepxUs/CIX2XLbGk7OcYkrulvUOm
ez62H12iNagbb+4s2FUzuKcr5aYbje7YB1941GKz4fen6xAggRIc5gzTM4CNmKd98xzTTaeWUZWj
zPAB0FLSA5gnQnmhLgcx6QfKdewceoqEBLQ0t2Evp2gc+PCQg+YMfNe5KkAWxi0WkMU2Hn/WpmBN
dtGuZa2OKy5kyyWZD3dTtQFNI1EkOHavKdnHf5f39tgt+Mf9BBB55jRB2xqp6Jk2BJts2mYm6Qdh
U6fQ9IaPTnPb+6YSYwpl+NgTAtsY1yOFnR58ys1FxB9QQDJ0PrxULmy1mjpH7hZlnovtVqWiMaXe
SEE152Rr6AwIin8TqoCFcIs0SvzXvicx0Wm22VJIdPR07cEAvSHe//76iusG0l8vH5gRHF/keZko
sEk699L5bLbCHsj4OXOzcJKhggiqJUQoxQVOAPqaMzYOCHbESKB0nPmLv+cIirwMlJU5V6J6RTZP
gORgoSpZl8iDdpSfv5+yasbzUZvE5TiD15EMuLm+jrRk/DA9bWrrGFrklyrrQ7Ap6bhOkKXyw2t1
DUTw8xz83PLyRz4S3HPxVoy05smiBWahl7ENzOBxsUBURcIghpYseA26dTJeEBa0tqY87p0l4hmw
FktnUB9PLQNyWvL4yqqoDTSmlvN4wo0d8m+akzAJ6YjarBZGYB9gCX20hI3KhtrhJO16NkT2psSp
v1vcGJVID4+wdmT+SnNJXPb9EPZi6o7lvm9RQr+eiZ6HR1cS6Hxl/X2SNlZZ/XwyGz7AzReBnplO
ddwpW0/CKryP2V15U/oWSZJ2oIQihynSHBoIkLBjulplq0RcNX3o6kNJBUZXqVwgdGSoX2EiOw68
PPGpGq2sgPC+LyDPcEn/LxEZbDOc3m/XxbFjpBz1U0i1ma2viUAE/TtfmbGnjmcWYBdkWdDCboJZ
GdpXRIp1UYO0AvlYL9Qxfh/+sFE49zbG63kHHrkLPUAvRCuv8OJiSbcdf3U7WMxo/t4vbqdkkpBp
LnahBSUUUEieNt1AtMtoXm3u9K/5TbfhNhuCNPGiM8rlMo1dX8XVUPSXwW3XIlgPSrLBR5zukOtz
HpsFcW8qN+NVQ+jHmoakBXgPu7XzPB3FarIDdV6VoAexhnAp5+XMox2xwwCfi5S0Slap4yVNB1et
dXBYu7yO9p4REE1ACgF4FT+ELHaeDNU+hIAZ8U0vTclFHLvLCHCLBwOzwuQqvLA6NeveBfuCbju8
oJgUYdYJtZY4tRkJOWlYL5qL/8wLV+Epbn0I4+uJXaV0TPm+duSJO6s/J6nTrJLySV/NUY1vFMN+
3Xli4tBFfmFVzmHWb6lAcNGQTCVDjetOHFNoyu/mtBicfkO4hwjlynwB6wBWS/C1/2JbUSY8Hytw
nAOssEtwA753qyqg1odB9bpzr/kGCqmIfv1rE770tX2qh9kjHb/jjke01MmHcPJCa7IEWoqRiTMC
5adBUzr2raY3+4j5F3LlyoncLyaXtYEiczz9UgfuClAzT4ErU7rwd537OsuZWoySR5NAm++/nxjS
OVi10lFkQOUuITfWvxG820y5KeDYSrCNGv2R4Hvu+2zynx5ov6CanvVRuzuv/w3Qzu1oTajSRk7G
K4eOHqVgcNgJ+GL8/AYm5G2FkNZyO0hjyP/1W+VwlgeOihHgj0zsnZlDXvCeHizABhqIgjVKKE5n
Ln1uDCtAjW8gzj7TpRgsZnOYdhpEJH1kwykAp2DG9tIKNwAMjUnA/qK9nzKcrZ/3aGL+K3YOzu/M
cf7+sF1RaFQP8B9Ef75ZONOnlrq2HHYuF/Z8enZVaAVqvCb7CkFCplt6kwuqaRAWX6u3dxTv5hwH
469NAkravROTnVyckbn1Wsv1PzzunOViz3Mi3xIbHBFC96ySWXj3twRd2yGSXztfpB0dgx2uE5l0
ORhIAfVBP9/ypXlRvHUq1PtC+eLS1G/YuvX/qppSekKSJwKB72YFlKJP5mXB4CE7GNKi/Jqgyc9Y
qiS9+EEXTpzXoZXizSrGQKmpxk49h5gpJUygLu8GvVZzFQ0RdrKiQkAE2b8UGbIRMQv/LJyQkz0J
7zsExTiwdKhj3NC4Gozypdg22UzefCFhhjOhmnUWI9RKwKKqYEDDBAO5PTSw/Fs5WYtUh7hPx8xT
GfxJBlWb/2Smy2G2kYUylv2KQRSxLE7aIFk1UpeyAkK2OTJgltlxM24IwW159taKmOsXF6g6N8wu
nKxUf799iOipWrwHFEueNzAI6Onb3w+Y2L+8CLNwQ+3svR5DIsdMapjQi2kUFDHFhjhSRLJwqolF
tC0S5sdpdihs07ANkaUE66c0W6F4B7o3G6ufOTmQsYa7vWmLVThiyDwwj7mRUjYIlUamqVh82+8t
1b76mh8Y/TEvayoMrLPNj0ITAlGc6WX2s15xOLP5gxev0/ckkIKA4i6Nas8Z1TgUdNW1smmFK81V
8QaMCEY1qi6GUuFiFVubu66//qdmoXn1oY/xfAq0NkKXweq8eqNdFvepjHnoFP3e+cuzsOgI23W5
DUB1KPRr4i5qleetMgb75VUjA1eVDFCjxvbhI53/3QpGEUVB9dT2qMikUw4/a+ei3UHPjGoVCRIM
ktzwT8hxI8y8rXFwtpHC2PuWVYp7bOY2ipf6uWTh+rFduc1FaFAwyRF+qpLu3mWo1ebF0CBbuI8F
IhnzzIkOq2KVIblVT1dH4CeFspSF5w7vu7Ei2vqIlKDIsVgWLL2mJuCqpiA2gWkYMVGmlCDcv2Ix
SamH5+m1MpHBhtD5zf2VmFxF+HtmVK0SWcIuyTQuSYJYyFvjstwgLFq67U0+dKoI6NXux0HBko1s
PI7VeD3ya4sV6sf0kpWsOWeMdqErwyt9IQBbYHetm+LoOMpbuBZH2N4tJG/EdUVKivnIa8oIkSqC
Gj03FOo8Zxz63CAM9GStRFXbJnfEA+Wb+rAo6/IP1AoLEUm8Ff9HEQ4I8GJJDWsq7mrZQQdp1SUL
wzL3YYDNQabNdNuHGHf9/yM/fPK15bGSiI6tVI/Z8ga1700Uovlhl+jWJvYPb5/espxB+TqZ9r2a
rlKmcKWxsReQ54tHoB5fC2O6Alr/p7glswuCJwE4VsSxlHQZeV4egMzLw66+abY95hD9X5n0Y+zW
c86lXGGWIXay50KoTRwdxpQJYeTmCOjt/6bNMuKpErRdbjQDF1WE6ZFptPlnc7WmNVMPBNm0jxPm
As/IMujaqwKmUqHuHInI6P7K3h7wr/ugVIDelNbn9OU3Lrom1RgfEYgW1srVC59TQAfAVEGPY0ql
deM4y/UV6Ycfe99CThl16nLfC5AASN3t4a1/Bo/LWJ6Hqh+K3mnGCpZwF6Xs3M2K0DqfSwSMxQjq
qbYRO8PYiaqxY3UcZCIYaCelsdcXX2OHIjy2jB3ExPwf7zE4VTsOOFi3XmpXuRBNqgTRiCixPYsk
cp/Tz+F8jv1IS5buX6wPRpumhuhIuxcp3pgm2dbMjdB3GttXFslFG4Wb0tJ8ZRcWJc10V/fRPl8F
HR6ENUTxngofhTGVy2J945faZs0z7C2mpmKlmm0bPlANXVPA6d916X0TbFNDuvAW8pECwtEgwQnm
jZKFtqIUmmWyrn27wNg5BsbUEJKolusfiJsUOyBr31dNXQBMMTa6aTYDCSaa9eQuW2KOEM2oh4rZ
NN0nvMysSOQI1bXbxw5VrCAVVwgDvLhoNy4GvJ138aNkIUkZOXKOFOZY1uJtYFEgcj8K5WtSgtdR
OO6LdwIcdqBKDZJyBud0dtNrdwjTtPAisg2N6KXxn4qqCR2jU1u92XTAvHMtxyu7wFkZIADuAV+H
M05W4B/wcW8//d7xV1TjLOQMPziFVUcvgBYM84mdkpXOm4FM2ULkLlE6j4wNPhOdqqBh183ID9Tf
NbMffVNW3eOxV4wrY9YwfL8NEp6+CzpUajf3Wlh362h7vUSXItfVYwk0BQacT0Kl+ti2uS9ZBA6j
6p5Yesu+42Y0q0zTbuN1zZkURDf2LMqBE23lZvsdGMADtQAdyVMg1nCa5r+RGXHxVPHhUB51vLxr
9MRYmnTtd9CPK2LV6wAJLCBnDh1dkFna6S8xk//LKvxhORHglCq78aAL2+peB1PJXDRW0xkfRK5n
zfr4oE+ftR4SfI27JUCYDJcxLMgLcH2KPCOpcYKkDbwRyxtI+rhjdYEXG6g/0lQ0DfXs0SUHc2GO
q64tycPu6wzHWgvqpjbGt2FmSMfQ7B9sJmPpqQsw1s/rbEN4Jb7gi0jOKcfk1hrjPqXpgz5kr/cw
uv2acCjp8e+DuGyrm3LXnYw8t7NUb/Lk17TXcJnoyfPbyb24UKZS4ozEDbI68gtlm8kibxtSm8LG
heWt65Tn+twDkcWp983E58Uqh6n4F5xI4iV1HMEUBpE+st7YrCoveJGpZ/Qya4zNA4DgbTLZYCIt
6rKj5crzQ6Y5LfuPU/bPEs/Y7uNxOS3646iW1G+ICYe4mCaLlGQXrWLOZn2Y3ag4yKBNbmkQgnG7
/WHFKz2Zcbd/yYK56oT62yMB+KqbCuYLuerFLKiVEtabzQWOsqcQoQRDbyQH0bUdTUZ6CWV95KUK
Z826RtwcMdZAx1oHNz/D53vHAnsyjRgJhn2iP3pDbf+hysbMl33r3u1ZpcmmxbcOeadQVg4jxv5r
JhL4KQfyNTI75BEsHXt5HPdkN2IxZqCwQu+nG3jTrxwv2M/jI3lqhoZfSE0/TcVgVaFKK1K5Q732
srI6j3T/Ghj7FCwex0orKXG+nU0qE74tAwqhqtEXZdRG+haEr/geHsatRQOKSBHYl15rx6hJazRu
VKWKCOmpE1/xleIlYNFWUPr2Oi7Rmalh5A/dwQyW6IvqoHa8Tlk+W7G4E7gT/7uK5+3b/yiapM3D
W3sE+V15zN2xDMo7RCy2c3CmIVbdsS/XMPPYOUusiCHrpyq+PTR7R79/cRyJupet/rHCvr/p6/L5
VVJhuJiZiIzlvXr/hIOJGMfQ6+5jnQvunx5WcVxvFSbKVbf8vQwcj+mZg7JFcPLiSpYHXFf1f1lE
XA/LkvQ7nuYfB6V70cTCr0btuzskTv22PUmyt0mviJ82N5ey670AxhInqbuRlch0juLpm0y/7Zwd
zWOEe7Ke/3zh68xsgg2FeDmU3+KuUYndbkGWFefpIGbkIsi7aFnxcDuQOcQ/G5K9YlEeBUeMHvNt
G+W8XKLoTgS952Vwy2M/mcn5ev8pEj0vxTDrhYV9JSmnp0SrdvXAgpWdcRuPPQbRXb2nSfBG/27d
XD7Std0ts/cH85UlzdH/bRbBrM7bQs1/UDzfLBWopfRmNYMyBEqCJGs1yeIFRyTpbIHfVd3uxizO
0WQz56n5UCQksiMq7bSEQPvQRWCIOeiOiKQkBc5V9nsBHHJevhFFXsp0QJQbCOcgPfQNn7pt3IcC
4iYXddXSs9LJVHCiVUg5HLmbvEhdaAxJOGvWaDlvCrHskzDFEq9hr287f5AE6pj0m96W2TJjvCt+
oQW0SCmaMMyrgOEOfu57qJP+77LWA3/jrnbEL8X4lU64bBl0hOJ2sjXCVHfTC185ZILBsGZPEWLa
KbCisWScPejBnlQPId6fKK2P2efw3xgT1xog/E7uzzF4JFgdebESqSgP/SU539w55pucGkRy1miX
z0SFAmae3V5k54FV9VITYNuP+kGzl9663RZgE2zrcA6W0ESueco3Mc5twEVl7Y1pnvMtffaQiudZ
v2Kc9x6sub3dAbL8foYlb+pVtZhCX26eehUOUBX1+a/V97B1Z1JSwZLnTeGr/V7tOtm6IVAygzqc
BBp+VeGCx90PuVEQTrd7pSgjcd4DZ1Scn9AWtlEz+S79cthrPMlqTbq7Axj38FHCeNN1i2aPhXKf
wRCjXUehj0DkutpFltdi7Xnvy9ehsQ4YkpvFrKyac0ZmY5rD7UKR1XcyxiBno7hpkz3XBe+w2cKT
Oo8B6ifqwiFfTi6QVzmQWWo5yDp4k015zAjq9HXmfBQXMw5Rze1lFyHlC3PsSQDk40DBIeMe/spm
oDR99KGaTgJJhoHFzbdfTzQuL2hCd691adriYcObnva5yH56angk2hK5rpGhmlNVjH5imhdFjWnh
sGWvvEuOhpbqAA0SkmyEFoUNIGOqeZEVdME6XFH12YBH7Fy5ooD0T+6L34TTL7eWEtg1Pf3pIYSR
ZcCdpDtzTWjTYyg2ar0TzuxcSf/vJzagPP/SwImhiFwYLyOt30dY+8ImrwbaMSLrQacdy8u2Bj0/
Y0Ms/BBf73y3Z8/BuwfGDWnZWx9xlY74mFD480cb9rlL7qbcRHcPoaenem3idT0Fr62vCyJSVL/P
D1OnncfREtHA1+aaASPt5JuzGVgeDAbyjju1PD6gdBj3OG18yTVra0PRF0fVQTxUKdKZYB2BpEJT
0P0GBHPPL1t0IKAXlgoU0amu1LSZaKWF//aXpDRh3NXdgnwfwZCIYnDJgtRTdUwleHN8r+Q3943+
HvMNYcGA0VZk5EEa6tExqdvYeUliFdmsV1S9YdzJ191ojxBGkLMseS5+5xDJ8yS9utUXEeL7kc1U
Y4U9AnnWtCl5SPiqJUNzYRCwoACSOT28SsRWbFzFaRk8du12ZgEoNNwwa9VM8Jt1twkvzJXYsLsd
wFIvcEQBDFsHqrPqRtIf1S3d+FXq6g/tXVYIZ9nLUUbMtWetufeSjuZNtX8R1t4XXVpjR0gVoOzr
EF0hE+6JMTAi25XFtyN8rbtenIzprHyTrNNcJlsi8iIDT+88S8zywtIOObVtuVeD9d8ZPCpozx01
eieIxkFYJB11eltujVvihnCw69rbui/StSF+lo2NfKLh9nc74fPLKaeIWz373e3QphXv2X4AEgYA
88YSr7crtdHUDzUwmS/EZC8dRmeA6GTyiem7s6tHT3OWw7gWmeWPDN5tCTXd6Oez/opKDsRwSH98
So+e81hERe3r1FZv+oz+aPp5hoqr3EqxwdId01Y67l6ATlb6GjoLpjk8qrDrfXw0iPbaY31FUskP
uqiHwmlSy8yVN8ukN1X4WXdHWg4CTotd+XLK8MM34V+VFfsFPZrLFNx8vV8R8x/nhjlRF+XlgkSC
Val01J/IwzYNMrO+a18wLfwE6xXw7ruxN9skKzJOkH9PhhfaIjgCO2fwSJ9984p8b6z3Z6RCYcWv
yBITL6uZd3lkp/HyzfHX9rx1q/N73x063bkzY4kV2dYesbwY9pdUkPvI0bajlDmzU3OJN10d1r08
OYSA8etDqkhI82A0UX1P9isG1AlSQWNZF/b0MCLGglJ8/kczhabYNPVUeox5uVII6gsMWvTN3loX
7lRxm15dxypjKwd23frRMwRfD4hbcXfnR7AQgBGmZuTd+XXriFgvbL/nvkS1ltLujBCtWfZxmrs4
lE26MBk+9YeN7tt+sbFe151ETcWAADJsZA7MgKflXIt1Zqh0ZYd1+L81GrHEzH2Iy10L0imn9TLO
WWJyYMcUepugya6kPL359ACzvvq4Vdr3CywA37DFKszs1YD55kSEvHOd4AfAZxzUW+w2J9K8jm/A
6f1fXL9rTU1ddtOvxeLQGPi2Zn8k4DsYpmcl/ItLQbYibJMM1bisI0ClrLDtG++2CvWXDYBYPVH6
l3ewkU8uzNueqZMYjbFxVTDmtzm7IlJLZ9j2pvBoR77wubWXge+FRhHUmzHc3btudpAa8EhWHAWH
mEHu9594KX0khPOdPPWXfZuVbrloPLCeQrpOS5OTR+v3K8sfmvqMJRAx1moLm1vyKJML9ilYr65c
2J3tvOSU571jLrCIJ5k08Zm3M6A0czJbZVMLL8gKvtMqFz6GU1kgcD5RzY8XAie/C91WJSzUIwI6
BMcfjCdO691WS97mZhbTIjwKY0kEslNWPyb5A8tUj3pAlgdvHeTkBu9/TUs49DxbgcYqkkApNlk7
p2YKZL4Z2Vec98//7cbCQjis4HnS8xjHNgRMu100o9B3wJrbcrP+3edcCHhPZkZOCc+GxkFgHMJI
7SNZVhKiQFels+duj98BEBuIqRGq5PL8DnW9z9F0KZ0FXuGkm3UhNlRB1zgd70/pUaEPxATnkRqX
kzd1/LHvaz4FhcKiYVnsU0a3Nl9HYNFvppnM0PHAQGuMKn30PxsoCYqFr6AyWUnsReeSSDoKKdGr
nVtLakrwXOTk0DJKiQ7GCTv8oebrNvLY5Hy7HaQHUykXJp5bNuBq/znrMuUZxY8C7Peh2iLeoX7p
AWHLx4HGmWRAU0LF6lifs7T3L51UecrAU4FfycN/388nMEGd8HgnZPf3QkT4Toppu00dwBGUDCHo
g9OcrADpaq5bEE7D+D3joRjVyJJLKxKxBXjXSNnltegQ71EOMLKpEAUfkWLBYfUcXn9vDInpj+lj
lKL5F8sal6mgWJTAwUnud4xE+Y7mpz8kEgSGnruQorVAEBsuuRSFQcyz+T/4PD4kUtS2LRs8M/S5
MoLgfddr9IeXQPwTF/eIfTri713cmX7Sp0lU13UoazYwbRkLDU46V5mGf/aY/sPxmxtG5ItQnuSr
fRPf1BrR3veliYGgldyqP/sL/r0di4xgMiXpZVZXGsRM51dpj+DM439Fz+kSdMg79cnKJ/G3h2HD
wrGim1VSh/H4EExMDvayuVu7Qr82Wo2lGVJybtSa2bv1jE5u53MuxiNKCMUep0uHagupom2lN1Gn
AAzxaejhfesK5LF6pYLQG9bc+oseBc9R6UAG2oHBcEBNxBZ8yc0h7yPIdJXacruXdp1Pw0Fyf++q
ZhZdRjieFQTUDU1IhuHU1iiFvPT5wDjSVMBkAgcNwxOmZWfNigRcM6nI0mP1INZPqNlcIAvEvsPY
x2PAYqt8ZND5E1hlSKCQPN473GvD8OrRo1YxdmU4tQLYYazg0MK+r+p4D+PJl0KDmIDp/JvGk04I
7DKq3stXNWBdnboGfdUOmVxFcXQhXMeinvVTF7UeUOw/VsiiuKkaL/b8VZHZN34zRT7rARhUavHI
mMCnrctjLiLfEQ+UfQCV5qFK0ehxyN4aczlSqSHwgx5KUK5jC+S6jBkZbnUvBOJejZxZs107trQO
jtVolexlRQF3qTAekmi+2jMmDE38S9KLNIcrk8bZ1rUeqk9Wbg6jKovC8zrIw48V30iffbIPx7UM
5MA4W3Rxz4vZPHU5tpeuJGJk1QUdCPX20UNmY7gY+hGFZeTasR4lpZGVKra2ZbHyLrj5PSEWyMGt
3s1fq8xAOBLx+xYGO7sfptIpf4ChZx4NF1XqhTD6jjs4iaSDBtffKfa68fgh9PWCGUOTrLALjd00
eKn5zQdpt6br52uytDkuKoI0LD2uoITvhgF6RcbleNy3k6Wc/kQbP8FhrCoBHFUhKwgDHmeqmahw
7U579hksSlTP4BjzWz55DyrmnNNHnCyprrQAkw3+VoH0wGNHK6jDfXI/CTOpSejZ3fV7yyV0WUu+
5cQP/gAWpngLi/bGQ6WncKsqoNv16hmiKon2AM2FdP0SGtqcWt08xpgQwtKnuvpDTnBZY9AL45bi
tQNzYGG+H2dn6FcYbLY/xRNyPshEEGWir/sGiewt1lQJCVoEPAp6eCYiFSTzm0eklq7/dEOz1kZ8
p93CiAgZKWxihQjw+VJ6QVtmz4jQC+j4/vNY/A7/Tcwnz+Vdmvr7Y2nOeH0vqbsBpp5bIi799VKn
jiqGEAskeVJjnolTVFlUVrhL9IPjX4W1gIijFXebD1/fg5OOu4cqhk9SqiOkqPME5iTvUx+5w++B
LUsy+qRjwUJVVJQUlm1ZW4QFit4xKA/cWcm41pwyAVLgFFNagYTGlHCg7ak8TTb8+gLbCLiEdwv2
vX+4YJX8QRZbnXKlk1qgxUXEzGfXS7D0lALt0lfOnoyRWtMfsAYof4+L8KQxtqvPRRj3qmVgTcH3
NFisVHRxxCSaOds78hTkqzJxVkKevj+o3CvR0F9DMeTBJ93ySRYVmAgFmat1WSqH3zLVBAwF0Ibq
QLQSwLTIx5k3mypsIkbJNXB0iQ9/WNMV7AjzkmwRAoNiD3j3Dt/AyiQ+3CZpapwDZ+AEnVFzTQQp
Z0fgnYdURLM2wqH9vKKXe0GXmK4ab56Pl6H9HlRHo6Csn8kVc4Jw22MCQcWqKikGrcfxeoRwmzKv
pFu0a/+uU6i95hwDl4eSUifOp/qbXnOXLpOHVUkhFP+ut7M/LglbPE1iEigAtolq6FmsIGbDk5x8
5lGqCfiJlwdndRyOx9IEW+6UDdKP8sSA8dsahVARDBTgqkhYO8c+NP7BQoJUNAC50/ArPo3fK7Eu
4RCNXh7RFJ9TLbp4H2CXfmCWmXTnsN3adwQY3RDbTYDvJLdvjXL36YhDnkHBZRWRy6UEU/fPe2KR
AmdvqPXhQ7u5Ms3cJPvi2ZcHgLQWEzw0bOcT02NugILoInaNQ9did3J85Vaw+N40Qvj+roXzVeo9
Z6Y4X4tF1MFMQ+9U0UPyh/li7O1Hed+vV4g+yARZlbylyTEqlBQwIwZMifLZjLd8GFDoHC5yK5Wl
OPskUTJ8dGiQ1XN/32nLEwAQBnnKMw1IrCuHLBBSyqjRDgZxRcLSBtWA7prsCbH5+ePy+i2FzG23
DfgCdm4HhCoDvYdozsRNrTnfN3y6uRe7xMPxZPWMzJuRcKY8HOmLbGhI0RJbVx5dN9iEhe+B1FDK
e5r9+TMUWxPgQZv+Q6EIa74q+OGocNptIMS7A2mihDzkRC4xgedAlb35ILJtZanNBBgkvjdVjtSM
JcVwI+XqaS+/WeQm7S+6pbGoX4fppOiAaF/fK28rdKNzMZYTM9OBczkc8Kxj8uXmTavoH1Nckl12
7OP0u0fC6hGlO8QfGE6OZfyqXOQXR3qlUFVafTo9GHPRlcOb/REt9RwZp7V/vrZVJn9YgHD9UZ/k
gRaxBxzJ3504w9Ug2FLPeMOssf0PGo7YY+kmRaCw0pBHliLcOpDnqBhD3R8H3imB1HTORx/s9dxc
vVq9ubItTcsuAdr4rEQjTOXbUVSVuaaF8Ucj+cUHSjQbGcU+IktjGyT/pOykiO/PeUsmdV4kOnKW
XEaKx5KFt3RAteIi84xgNzNU5vQnMl67e8quwAqH3I9cttKqAjeuba7960tPhe0YBbWR4eAjPp+m
Jo/WQEDEjvsdb1FKHjKOJBvjrXS9bfi9rQEcZG1DhPtJW81D24Ot8zuFGpsLFIC+N9oH4lVjiIq/
lJVa1aw6OlJnQjDsVPsqlB9C+Jxr773iiqtDc3yVOigmWkSTkUkt2PSwnpJCok1UiEtscW0zmb3E
InOCuOg45gwTKDNMxvx6iUfpkoy8U1d8n6dEWYL5mq/2Cx1a+tPPcomxYe27/naTbqQXeIwcnARV
zuzcp9MShn2fILUaU7+GA2zuYB5DgvzQQtje9o961t1zBXyrCwn+qRPopO4XvMsMBXtgefc/8w8s
rqo+ZXAwTjSTZLfh+T++yMScKG+f8pFhwiPOJVT1MzaNeC56GqB+2/Qs7BzPjYjoo6zYqglNA0xX
NjZK/46f72Y/2t4jlYnMLm8kIBUIgp17kmoSkbiqoHJ9aLi+o1xMRPKPg9Vc1+oB+PkrCAMNT5m0
vsKhL87IbCpFLPT/zfdmeWILBNpavAjaEbtvQXNmqv5B7xEiE7da8EAYhc5ZO8XGdPdazBfJMOrZ
AdAiCUH0aNM9B3dnMEfofLwIqv0c8diBfU+iuOQC9D/sTOyW8B8FxzozJbGIl4HUG7m5EGG2iql4
tvuOxP3YsI3eIK0QGYXcNlgptdkayzJKte7/GnbBPbnnW0MTIPsffnfNYlu4vthSpKjLhxPopWqY
CgSH3T2Lhn18TF6cC0DLlwf3VgPxfQ4Q+uBLdRJMp+r7kGB7cISiLxluzQ8/Wk4lD4o7neVVnKbb
GDr+bbJ099GlUDWcDd/1q3SzKBIVO30+leOtepHl3zZyOZtUMG2zLmjcGGL/fPxBqCskbTo3rvYt
fkP29N6NuXLxOLUClFKVa5AbNAqclBpmg/r6W3ZGkIHKgcE2a0yN5+CPz2ZEpwjVJfXF/QoOfI4s
mkZ00ECRik36ONBk7MLr14v1/onauAOgQllTg01TQhX3hQMVyl2sd0+kkx6CDE2OfPKTUolbqc0p
IQyMQxZjdvz+3q59LM5+/e5+COa8eZ40iVZZlGSGv9QbZNHtU32vN8l3agrAXTfQQ1rxB4ncsEvW
kTL8P0s9GaefTs2+H8fq8I/Q4atGnfzJOmPvfqs5X0ysoe7nSDgPx21NCryGxxKR184HBFlKHhKl
j/c+6XE+/SzA5eVHAZkxzMbrerwy8iRRb2YVl9+1Ma7Pfq7TXkPWTY2vxBFI0NuBhTXP/nuDk+Gy
PCYZCKyUkXLBq5bBl4aYZXMbO6vSN24mMKhsX4zl4hA3DhK/ihb41lvncsgw+1GnyBB8unV2Iynj
qUaxgO7gpoQJae5nF3hheItGnG9BNDqpXsdrDVZpdvXKYqwJAksjWbPczqjIFRU8Hddl9UujcKMb
PPB0aZvSscuM9e2eWIl38cBBLtb+JjqAIXLAaX68G2niMt0A83m+YopWSkzKhq8FASQZ72F4Ctcn
cLVtQnuHrLQ0jnz44HWqeoKbPBGoT3dYF6LZDXVgLpBSXD2n5FBp0+kBykouOiNWMx1VuoI+z20D
OdMOqnJffxpGJzKVenVjF0AJo9oLwhZwBj+YD6j5mvABjjIcLBGPyQcG0k3rDxzG9rbJUnlrTDWO
4U4CbAHpEVY5zLuhEjWrikJ2rUHpAJM6DSU2z4rXudoLcNISbpUOb/3iDjcT+Ho6c6jciO7k8at6
AgBqovA6OMEe/ToufDQ9aEsPi7DTEcFYEgjxRGYcj57G8M7fwlb1aYdn+L+jowUvcFUWCJuI8eid
iBKkK9y3UWStHH0ArVqeLoLh36R+cGN2pUsl1zOyM0pFb6i6GweazDh+KGUR3eK61I3tesk02FAC
6cCLswKAyjWdIJs9r2f1NtdU55+BYxwqQWziVeET+vacNE2bOVgLj1J1QbTv+Xi/3nKUCmeOJftI
kV71Hs2RSc9RK/0i7+32KXo1Ma3nBUGphWozJBg5tbTf6Xe5U0CGLJ1OBhnZ8a92WOQ36GYQ5miT
goZ0hjqrhYqX6hdc1g5rv9EB+Zd+QHI6N6vg3i4vtbMiJ0gKukb/zEnWlUy3Ov0S+0mdSMJYw3OI
3NIvesSETXJcDK/y60DAkakdUsFFgqZ1lUW7NzrDoK+3BkAxgb9RuJwrvX1f06GnKEgUXL+WAErQ
6SZb6wP/nVLKe28+oa75FFCc0+TkMkuXFHIiGGdVsxIzUJeDFE6VXUNUhIU14jdroqMyhWLzL7RQ
j9HWF0d+3naTkvYiPcHzSKDqtK3znb0B2LEbbm/asbkc3sUmVSnDql5pfAgitHLQhUXQzKTOn0/E
jl5Zi3gFN6XUpAzmRxW1Zlg/Nxl8zBZ3fFS2bD0NXhvz/E7mfgHvwH6/Q3EKH1g9WRV0KLBEXlgT
WDshzalLt3WlFCrS4GuS1j+d/LvxIJAC6yoJRIOXza7JmCrBKejD1ASpOLnUhhhdxaisi3g3BCij
aTqWPLs27NTV22GzKb32HUnQMtPqZRN7dYe43oC2VDLLyOmArcZ/9zbQKJidV9TV4DvAzbcC6yMv
hc70LlzYL0e8OB35pi1QTzIJO38iEU3AFWA5RzK2jkw3y/JdmCBnBrz9J84PPUTWESScYMm2tPCA
XWq1/97UjKrTJrkwEl4NUJxBjh+bvVx64NCjtCqLBQmF5xnjEn/P7xaHLzAA5ZpFRJwCHImBCFHG
cH/Bpmdg4qEiZUlObfgFqzu00MjQfv+H9f6nB9qi5vlHHF7uWUGsuaSUss6qvUw9TLad6dNp0f41
g+C7Nff5iv9wrPIyIer1P6Et4EYJg0rsOLZq4lxAS7VgVIGuO4Rn2/U5C05M+UQtW0KK4PFoQYp4
cn6rmrgeW9wO2vKB/AZqe5li/eq3TF+7F5e2vswMxHy7oYDL5xkyhpV7TMR3+e+63xkmh5qdVLOJ
rJeWZUZdp3fTGjz116DQCDnVf9nq5AH/i4kp08/MjREyzDm42g2F5qeHO6FtliFsoeNqY6aLMGte
Vu/G81//EFPFAXK+Bsc/U6owM9nzTae0477CjLRIL+P1NGAT9RFRE1NEuk91b1MRQ0VWH507HX1z
jFjrCuUm+tB5m8I9h02btHs1t38yUAFZkAd0CALRQoGtnm/qrIg0M3I6FyxBFZDyS/SMd5WMXx/L
Gr/HbmQdaArQtkhnaMQjw23rYf99Tx6emnXX5OlL69x6kxx9p2qOhVIrAkBYnjw1Xxg0GLW+aCQ3
Qjf/1LmDy8Pf2DVveL7SyhreMD/0vytj9wCY/KqJxmNbDTrZFgHiY/7m8qo3l3NDLwAa++64jJfU
3Ibc2cvlNOcJLf+QTLGcrBf+OYbLJPs/9OoSuluOXXQFRxNFutOEUR49Lq0v4slTy2388wxWX1Ld
Mv/hikRKg0MpMJNy7phpRXfiVxQhWZiH4nS6TEKXp6asDuI/Str/K8jktn7jQ6Npi8uAX6ktqyHd
N+Zmj6qdTETEGPeINKuUeX8P37/hRMF42CtClW96prxQQMt9IQJX9a9pXOwa5xLZUOW0BmQ7G2nd
U23jBO/ZrYTRrMa0VXC/Is9onVtlNy4402HT0vTlH9e9myonfGdcwszGsXmzHklYRfkY2iPg5MZI
penaRJ6Y7ueEAr+BsMKrOMNWYfX/Zt9oaXuE88DRdopeXNZiV6SYFJWN/zqe1SfGjJCZ6KJNT1wQ
dHQWy26k8u3JuGw519r0YA9S6AYsjjHT+AnjkMWrdzP1Bo6LfwDtDhuYCvnU4YoDbUWXKjb0bwuu
rPXBD3hEPAi8klz9q8r1vlrp+8bzPIIzWLSE1CviGInSvYunQPyeUFa0AZDd44Cde4Vjzd59J1Y7
roDfQSGm+x+H2tchORdAjzV93+AvJKYY6iA/WoOXrpUA4r5RgnW0dE8JicYpsty2DfuiVj97y3yF
iHNnuS2v1E1UdThkrJysvH5nN65PE8Cwzz4VlAk8EF1782rtNQ5HsAoffxGePo03nCuP4KH1bEF7
y7uoBVWKaOn60UQkhgNv9Wz6IrYuSPN48jdz8uAELzdLHL8+of4FQxM/kK/9I1eSmzsIhFchWofL
qLW7boYuA7jzvve44EOzM9K2J1Swrbb2OqB70sUFVVfnjhHO+qADgnNxiMlvWRs2lmBvQCfRmLvN
sRj9EoeU1Pm+hmZSFihGp78zYG0W+GMRG52LGSMpki0IMsCKJA0KB3FhWXuvAAYT5LrqE46euKpf
X7eaaso1YE0ynA501XkfqOKeV2gM+4pXRY2tLQJZlOM8jSNN0ZkcyztcmXJElSnynaJTeaDutDft
eZw1m3A2bDws99X4MUyX3OW5NmIrtqtVwmP/yCioyOqS+Lg1iN0PxDbv+PX4giWRuqwvSLQvbta7
F7PAljHcYFBSL1DE1b5V+N9W0PPWTE7Ivxrjgigxb3pU5tKp733y4FkrjZJ97+Yw4ep7AAgW5de2
hL70f+J/bAwqtCyBXtKiDdZgCFyMk+XyaEEbjHeqqqYSb+/AfV/NHGG5mm/+LBh7AZPEcB0fabHN
jVqxQfAyihvuBkVZDNJi/zPglq8qYkyPIIH/E0pk3H3Xd0H6AyXxguQgkgqQK/LBFEWVdbYAG+nY
SirRqNSyvBU5xZpWFZZjzwV6sKAk4aLEPCstS8JXIUnqA2sAoWn2/Apq6U0TT/optiHww81IsEyh
mxdczbcqz38PoOrcrrh8itE6XXw8CsO3VBv6B85+ZqXFU9E3OyU7K0VfLOHgsKVOKLlqu8Lbb4dO
yd6B6eeEd6a+JRplXQQv58hg8JmPExWOfSn2bwxYHLlh0aqa8XxrxVxBwejPlBtNVaQA2d2Sj/+q
5hVNlgK7ySIt/WMx68JZzRfA/BRK0L6Rm7XbhZvb0xYRTHt0o2xSR5axe/zGWj383Y5y9YfN6u10
Fd3XzFDSFDOQ4h7lEIl0O4K2hqUflnaPDyDW54u2MyLkmLYM0Xeo9NdlZ9gB0WiMBbdWfdUSVAWJ
gIfTD/cGD8lnpJu8O0+4kgZcRaOyz0tbb6QMW0ieAG7E99GoW63aosRoPNHAUxoyaLDAfFIyTBmM
qlmONgGhm8g+P1kwwU6zpSOTHT4WWd5g5KoYWrkkaC5T9N3H8kq857/7pC+s5+FqRfsfVNksjcdy
kFY0cPY7Hll23TcVADb/Ul9UCBmni0HJRvgjTmxAJYiYwLTh04ix+jjdAcRzjCCaJVCVJmGY6f6c
1v5+wrJBRbsy9ryYtyGr2bNmOJogYEKmUJR0IW85XAmmtUdmXmUxyRG+nYCm8HZ0zZ+CjCs14+iT
5YSKHvxcOpC0NNXMg7qDOfEC02wwmA1+NZzaC+JzrwgsEv5SsUrWikjZZxfmTOemOwQ8Uv0kGL/9
FHALOrmSvY+oJLR6C6JIr8tgSZ6vCUX6leAt1rqcXfJhew7VVUEIMymGvEzKsCh1WhkPY0t3qK9T
f+NwIOMYyeNrGKro+DuX+5KbHdHHHZgCHAJRaPKaNG8ILiXHe+QLE75mfRGtygTowHDhhlWYi4i7
r+bie97Iedb63eFb4YjjIOzkXWo/CkvYMd2ZKoq45hMYuL87824E/RP2NlZrZtpBHsvNIHgLEHtp
MlksUXPronlkxpAM0fR3SzSdfMyPC/PGSfmi3pGhRziiw3XRmb4zRhS/BGsHWENIHHLrIENd+LMc
3iOteFapfhGMDPnraBkq2UL1BUBgm9A3cPZpJiu5rwBuHDmo0i62Ma5YmlZniA+7xi23lcdAQc1N
Qt7Hz2ucckyyCZ0a2k3X9UE1cRf9gZpyomIdJt5xPZ0VQgEqvkGMP+QduS6QmKWmx6pa6Z1cUfIK
VKiYcHtgS4pE6cIoXlotNAvLrX07hVNL2R264G6/L/DzPZrs5ZwSxPxjtiLD5AuSz8/Lb4I/zaoD
QxjeUwr5C0XHJjFm7HX/pk5ivCbDx5YtLF0RxOrF9s6x7SlMYG9yM8jIFB1RlaOp9b2T925i0Qi7
c6Kn/nPo1o4148lGeGNlaeZwD/YpfE4G7fG8IXRVwHxRg9RRhqN09/ME8LyIWYM98/5qJ33STKFo
/227EawxUxuW7hCNN9wi90McNWOqyG+WdtgqfzysjUaM2/YYtaixJg/WmyCzQ/FBnY9wjx+UvuhV
RCD9QSJxaHaHqfvypDNLGh6Py9Sy1y4W2hOYvkekIq2xkAQhE0XuY0aA4whDAu+wRvNB/GUjNWs1
jbqnALWqbK9U//8/w87gudAj6RDj4NytSEV+h9Zau4wqjzgmD9Khnm64MHYP58dT7ECLKTGreKRo
HpfAgo2JpwAkdN8Zd+YT9CC96vjcpU7hu3m2ZfcKYnIUBZ5bCfkewHtO1x4nvXIf8KvtEfj6Jbjn
tQ3OAFUuTlbGobax9EXH0/FyyXp0vT39+wuTPp1rJiC0mtcN8AREGwXeJRBlfGygq0/3nCuT98ib
WslyEdQLm4z8tHcJ+BXAXCijJfU2RWQOamIsH7R7EHNd9q/KNyYLJeRP6m8AgSGirfmlXbXPJsNk
l/kPI/zVac9BOGALyPylrdiFjaknUvy0OmEJsFwt3rkIaFrNLqP1+wOSNBQnr/11pNOsRe36mCIR
6XhxVGEFqmoD6BytpYAT9F3c4OJlvw5TOeIOS8l02il43IR+Ql1hfs3lNdxsMTW5ynzcnZ0smZsY
2n+/ls2ytMduCchfK/WbVlMB5B0RBkT21D5FhBKzOnozMr7roTtAbIJeSc6SIkVhB3e2LnEdo+tl
T6vWNj1SU061i3S2R9HM7iKqdIEHMVExFxNxaxcOMw2lMiBZrJrQXU5HA2whTZSjxq3mEPJUTRTS
uVMin7GWySbWV6+7DM/Lxp5Ha7mfRPHtAfG+8rKyLZ63Gae+cWmrJ1JMPZ9nH7wlx84U7R/WGhsW
wQ9czdjSi3Lx6HpN/gyW2SIdR5WueQKlSWVes3/Rn+6n/fksyMAKjIdi5sPFL/L2PzpWEiJF9ntn
hHCDotbrYsg2obYGofqBexcgVZXnYIU6GYWSgyG4uUPONSIw6d450w8bR5WzQCjW330Kj7djWFxU
gxVGc1Trd4WwvJyu2ns1/O5ZWRURiGn4H7iiA0wnq6N0MuyX38p2nKemYbka5KwLOxyh8qx9ASOO
SJBH0LhLB5yllyDUN3AXzOWAkK+tNOLFJgxqKvSpaKldA2xkNVC/0UZLwDL3fqmVWI0RV5zz6xz2
V4fTQKVpSyDKLC77D2SCsSer3Jg/MG4iZxIcCYvSJGgwQhX5y5xVdvBfihVMvRBapOoDLZeLefKY
CUlknit4F0pbTfIXoIaXVyw/MwbEMfOEVZ4Bi7X1xVR157painDa6u5IH5dMKfDA3FR7wfVdzlx3
ONdfYbo/H/BTkRIAFGFTPq3aVMTY/APiwpPlgCer+hBneKtWvPjLr0kuKD4iAPMFMVVKUZmeeUFh
XbgUOTvK1BtMFgM5xmHI4pw7NBuZib3ADNnRdXKm4GDq85nZ43m3X3ltJaIHSehM+hkqLy4EpJED
kjIQYyJ8JY323C2v52KAGmdSqVgSmP0s1XnYd0JH1MNsuF6cD+yAAil2jMmnGpLPYBUuwOASpxNs
wYQrWoizDG3C63N5iXGHgWkhjwdBn0mKtNcQ8BoJW+H+4Hv4tr71bSOyM7BNOoXRgRCd6A7Qe66M
rWzSejmZiYJTknngODx+hu1eltJ5AVQsCXxhl+dAVLVJHzTbO7bTviygqQdmUtkczGnL+cKpCDhO
HIoUJ5ZqPm74qXmOKkCNUuR9tf7yuZHS7Uc43EQ05mMrFF9PydXhFPN428ecAWgZ8/fuNCCpyBDf
7XVd8eXzM7Wj+PddmAqX08cUbtjtcGuSStE/mPvlOGcca0tFxLQeTRwxlu6L0squvnhAxdPgWXm2
PyatZibl5PcV6Pq/b4uh2YEaypP7tIvYsryntlBpdrbLlhspHWZfJ85tKbN8EWc2NGV6nikvL6Xt
B2jCodJ8zSP+6LOt6NhleIfktxPIcqiNF37/I0xxvLCcI6FOfQv5mlpihBIsT/zqWkU9Tb/GQ4kr
zbxG4b86U9WWhlKFBXrhqggCdBehR87U8Vs6W25ZUWJvZQzg+6o3F2Mp/t02Fifv3/R4gxSaZ2Y4
LVdhLEvIlzbDwx/G2I/hyX7hY3RwZf6g/tIJFNwHwRCVHIR2qbQljqjOSvACDjDH0KG8drEgsSa7
ZsVEXQbXKcZU7qYDHBJ+FwxK0Rhppjw9uO7HMl3ibZ4jFaElwbkH1T/ze27iPAdvDcdgWenNVTDi
4feAkzRU9GapG+EvVqr01vs0jo+I52NYOToIQisT4G3nkNN6tjuFIyZ2KWCuMRRDqVEo3P/Fn7IO
Tgwe46XIeVPYFtUWf5XTWTZcu6on1v3sjRaB0KsW4XZXbpWjrubqvGfzyiD6bcG4ayiaHyvidT8c
bM5ScGmJizKtuDNudmaigVBQbqvzp51O79OWqLYwRFI5g69hjnNeOsPeZXKE1WvprGYVkv9tiQnO
lzyxkz0rslp1hpYrMKGxPOkvpIjWyYzLSL4C5z0N9S1yuLxsm7DyLniXhLtkTnrotht8b+mppIHQ
A9c71ahOBcHFUyowte7F+l9vTcCTaqn/gs0zO72czx5OWohJzgtoieE1ouZNcUyf/R6UFTjoZMDJ
zvn9mxTlOTldyLZV6e0WHbeda+y/V/TVxInUBalzX96bC31wlwfIf71aELsP1R0v1p1J8HmsBtE7
Vx6r+k6pZ58gehmCmKDN4bB4YKAroj4zVqh+zCjsBevxwZDUOWhbdEYU239Oa2wAe+4PwbgK0nCR
VSrT4akwPwDLxoy4e63xEwB2GnwQ+C5QMnif/roXk0mX+KZZXPGJOKt072D6G3bopE0c5Gu8AEFq
SoPDVQPZLAO5RZO6bRZX+IBaZyi0fw4+5T138C6Xy1dqcTGQhVg+a3BjZw1rrDYpInCUOOvkTbrq
qINmV/BtrTYjkqapVkWNgXaKmp3uBF6gzzhF746AnHRs/YvK7s2YxR1oOsE2EVPSk9ukJYF/L8Gh
t+AXZkLl3lMxQIXUC9c9w1VCHLUpqjB+0pp4j3gUIXdklTCJBEAYr5PuWZtmKISHqyyfpXmilwsm
39ZeQeai+dv+/nSYa4kf2q4k3pw7ONhTgI1dn1Ff3AYBOoPE7ibmTawYq/sQ6tiezcUShehFNpf5
bodzMxGe5kmXVUksYYntj3Yfs6phkBZxvulFRBqK3w32kHqEreKWrjmwetclhPE6ta+nHuyY0fED
eLb8D/C2gvBWSw3xvRxxt7KsicRc9IYx5Mjov3IvvMUOGZQ5YZLaU5ocaHwxcOf/wRAkubCXxEbb
X++SnKh6gdMHP7bowKDr/IwgcLIni3+rwtYwqSTFr3H6OaWwepeIDuL5mhfPdOj9Gnwx8+cvWnfy
Z4wg4nHJzfcvZeUSxKTDm0nUuOxWaK+NOq/p9n6Pk/6EnS4wOkFWmYe47H2ZnZWXYc9jgGiCZx/o
MoxB0DyN0RHfAs5uBIXseLmarwcZeJRE3AnrGfCzFvYEdfBCebo0+4ThU5M39jldwRSE1obKGydg
EULz0/qauXghz93NWWx+ok7HlBkZdslt7NNvrH20zcnWVIjV9rVocYzrc5LmM5L1TpT4f+TNkhF6
hniqYhjuyzWjApaycHPSPixo7Qiw/RAtW6L2yxlzWdGZkz3zfnpmyB6MHu21hGJA+/uG5NWL5nDa
Na+xOtElTkA0Vze0L2nNlsFGdQKacg7dxMBTjVpZv8im/YySVLamZsRvHiikILxpLL6mVi9Qy0u1
S0QAolLfZ4dT4gWVYZUitrFUVDqtavSFgCdVy5FvkRm67cH75l+gWjF0mVnFITFjNXkZx7riPKPf
/bBByF2TYP1DD/xB3/SZEU4XPIhALK4v6IvDNFDhlZCa4BY/RB0PciCzajb3jg26odjf7wrc6saN
uB8beCwqqcFEjGUHX5Jjn2gEZte6fq+NMHowyktjPsIVTm+Kk/gLrfkdV7AWikhUsLbsGQCHUPPN
+15ezsL6WGUw7StG4wcK/rhQjL9ILDmXI5FDyzW4/PE8sa+seavB0ySfeCJRdwpoQHVwRRtY2H/+
oF0EtYKGqDhKS/4EUJYLDGZIfBC5S1Z6Yo34wSd0S8lY4vB3XzaSZ1jqZ5cqe0WMUVHfYqW8GF4m
pzRuRLPRS4J1T0ix0ZO8/fvEY8NCgE/aPyXka6+5vzS6zboSCBur/Hly3eFSaskQvBV7At+A2+mz
SfUWxtC7BG4T+6P4x3v6c5YiAwtAff/Was2ICw/WVEStbAyjzElCXu/7NUm70NCMUoM7A6BJ3NuE
h2/VJE5I0TKmVlxAzuCZyl2bEx/Nmj2QmjIuxn223rOtdNc3e5kyWqbZjgAYaoPvpX3fyRMOI8u1
1YnG+YPJcSTM+L40vg7Goysl8htPgxpgzqiTsBg2KXJw0bQ0qp2C9QVWMA93RtCrNRflZ6ruWa9w
jA0cEy0KG3yNkEXCsHKFqhlCmDfmy7JtGcK/QUhPjY7usC6i7r5oCeX5su9UgxeDKpuwclXc/Nl9
BFv+g2qI4Kt7N2awa3IjAXXNP2wV00fczpk6Q1f1qC+0FCBScjScmRf9QkB209eql/LvB/EDGTP0
z3SqaquMcu8EC2L2EJaSaSLH4xGP/VaFFvHEJp/mA3wzM3Ravn/C+RD63aQulGVWkpylCX0tbwcj
VmySp0vC0pOuv0CDofr3QiuEvEiv+uOygw9Tv32EcQuQ191XeanKi/kz8VGpMIY3pUHBk+yZwxQ5
KBeRZ6APvBjHOXdD1smCccaOBx4br2FTV+fDo0JoxRtWUL9d7gX7FO+9E1D2yX1JjIMLuPBBfMPx
SSCZRO6UZNbgAoNA4+9Xe/eB3I2ZH1wnXTtf+FCrEj0WBJiLwUqfIOIxLA54Sr1sxoy/kIy0Io15
to2ICYFlYOpPHOnMfCHSQXdVToNrWDcglphO0zsDQUnUn4i2XEQyDVcnpl2upKfdhd4/8f/sDdd2
yz6ACH5qbTnRL9OJfz7QUmq7yk5xemdVf/lH+6YCr8vp5W/gmRjXwKIOvOWI5xayWyo2jQjiEB1+
Ej1JbgOddGSC0CUbs2rRPo/+W13Y6CZ5cljkOZKBY2w7DwYiddcHVlmJhmKzPc1qphpDGssBr2jE
kdWWBh4Guqjz6y+orBb97qojlrnhr1eq+uPi5zSd5rZjwo/0Po0l4BwKHEsL5FaZj3eUZYaWX1ms
2y97qdxtYBcPaerEX6xoFh3/PT2WAuor/GOga2zeAGEiTvcpqemUwHz8VcWd7R0Pzv/X98IwaoU3
RghxytQ/WZy9kSmzsK399+oAHMuBxEWQGNnuQS1N6mahdSrbFHDSNd6TRQfbaKSGRomHO317NotG
AvvMeSu1Z1d++eow3lEUukxuTl8mwOip6fv3R3tZeaUPD1O3K5wQxg3Q31hmLayDCKediDFzfTCm
+1Z6Ng1K6CpkjqAAaUhfLsmrRZc0/+lZ1z1TEtGFwekLzdkX9dxU/JZogotRaE+JhCchrVPhc/Pu
iKHRl3fhs7w8n5BbFaeMKF9CcKtQs4dS6k27qQJ3LXyf/Uutflxbfj3eIyxfjsEsLNGFFqjdxSHy
ym5VuT8v/RJYnumWvuxFnMSqO2qAJNRlejUXObHxrRnqMjp5dlYZOm42GgYigoMzVTs2ImOHp61c
94mMdKBQXTfXvQ+FicAF7YPiLN79bPzMF3+q2wrXP8CKm40CQOLN8rlIYQRf6KrUresJOhVI6Jvl
aZldOuDEOT4530SYTyq+H2d9GDPg1UemVjf2Vnve0Mn4NJztOQ68YAVLF5ErPe1rU7xuq8F2cCQs
qvGBsm6cEOziQrVDwTAjE+AOpKgFog9kbmkQdqGcyZsreSdvElAyqrY577vpsEVz0w77gVl2JsSN
Yk950E+/odos2gLZGCPKNPdAgSyMzkqMnWLR+WS85rsqTpiYrYuqmIlStDm2cgpyiZKUJxJ/Bly7
zR8Ai3Me/y9+fwtx3qq+W111VIPPCeYPIAHT60GyNl352hV2Hn0ErfteVNCM0B1U3ItsqNujX5/3
ns+eG1+4vxdDAGJqtIMleAeWEL2n2lFdiA9JrcPVyp6xr4fCLmSZXzA+LWvVGMlMK+XEE1Yk+ny6
HoY2g5RPo9m88RD9mbCSZnPvsJ7VL3poy4elfZiWWr5fMfykcCW9p0H0gCBUe7cZYDygufkoNRkg
NBCbINe4tYgCR73WlfkPGCezelPinkBYhFH1ryOYCpvBmZKnuECG20TtIzFqc6KJmVwcF+OdJqTY
XOi1LxmQ0QuOBOhSMaZ83VnKjdCwSqVE8bNdDN2NCTGECqrHBHLQwD+HRtiLmtqcD0UTYidHFlcr
XCgSEB4YeGoCAJ0bBCbbzhh/N09Au4xnCnA9/IB23d0TJBVLy1BzfAz4tK9DjKKr0WZdyv/Veg9y
QG9Wv3LDAKpJEAMCZpRMGpEzdOSiEZCIs9VZAYKrTPJdUnC4GyNpoNf8MX7/OCW2GGymTpLHR5/F
ShJ/T+VBt2KpH2uVl7K/nKrPd7FKxKTbH3dy2xllPWdSVt8t51Y66bWnSi8TiTn1DmdmZfvzBCY+
kviJ4vGQNeyzEeSKW424ZjLr1EXQiEh902t3SsupljolXgmPd5zjVdszl5/xSUz3g9fVAMDrec4Q
E94VH31uza7yrNFhjqhqIj+10M4z0i7QcKD79ji1EhsIaybCMQigjD9vNBJL18JA1Al2yRRkLepa
MeooSCORKaM9L13Qs9tPhK7uvNh4CoT5m6jVhUZEwgV3ksMEDSQ/llRFBgvzNIxArrqZSslDeiD8
3WIVXU6Z3f30/9ntMV2WlnemV2SxD8vwZDTbFg4xjjc953nlWCXwwqYIcmG4rfjIaaqcAlREW852
JyxMC/St9jN+WWypAWH8hrcrpVvqU9p6H3uYZh0F/BE+BuWq3crxPLnXB7sXKiJ22EJDtHnO5qls
DMZ3Ay/bh1Nr9iGYGYv7ak53rp3QSR8C13UefrM4f+SohRYFYFW13z5E1c9ByXEQIt+xVOD3bzf/
8O6INF/Qmz5j7l9+OHTMsbwmMnN31jfW4LiVksxPU+V19e6BbAVF2LiCkYgFdrf7vD+yz37ztC5m
NCfbxgzk/curwFzmOUCVm6z33B+9+LhIErTc69m18LuseZvV68ZGLlRridTDSfufq9lEbRxthugl
DycS6aZEjKUWSh54Gv58KZUv+ThfH849QEgzohbl8lW93IEqaL12R9ynUdEOpZq/wh86wnF6YaQt
1ynB6R6fLqae386e/1sjRndki8IjBSqnRmIIXQJWYpbhv1Rdmr16+zoXW7cVVE6gMy4dCaYFqX7W
V+be1Ehu86XaSrgiCYMNXMLNAMcy3lLQ/780rdRCsmaoIZXBygTRf3mVgSVx/EMB6HonXC2ITJzG
ijYCgcbQFBMJsgAmcsSuAyhjJBmMWCpJ9rlSu5pHINf9Hoy0fM49ni8hoXF+VDPFnDDj7OhmNbLD
7kSTuHkoUWdcxbn1FA47xiHUj5BwNMWvAhhFO3sY2f7bJu0ds37hg9AHGsp+WmU+l2lAr6eYRJjR
CpGGYTQmJD9pJlh+JMVGsFBOrGZh03VJphZ2OgIuAbZGaKHgcDDVP/InR0X3AZWgK9dTUWTKAOHH
NyCtDLU3SYYAbR3NUHva39HEYB7D7Kd+UePhp2nj/rX4zoZ/+mGZi0DG1FOfAcpF6qjS4OcUWs4K
RX1OA8DMs5DmgsNuKX1DdDIAir/fr+qTdZMjiUmiNwlG7qmBsyTLxm3/bScMUm9Ztw/2yYQ9Hsic
JRbwfjVrijn3SCjackiQeYQgqDvjwF2Wbmd7feyZbjk2qg7Le8uIrims0dnvCtZmhhyQHfaAIS+Z
Ma5HKnNhQM3y1IcrBVShWxzauyZQv1L60YL1oOnOIchrCLtykseg2A3+mulaymiiadb9bogAucIl
Q39HZaUiCFITKzbs9pe3dY7KHhAR7JeEEPF+0gKrbGIYuJPWfBJxSzBCOoHByZTDeqAOMwm0um7T
p8l/SePgMTXS27qNUzwRz2t8hhl7/xsIRuK02w62mUi4FdVzX1qtA4ZMIO0MNy7xO+FoO4HNSZfY
xj4yRSbueCqHOI2QTRwG2CbLWSbQqW3/75YQlEMWAib9e8YjRe5AarQz9jldRoF6d9r0DdIOs5NQ
OhQDivCEbr2TlMq95e5YwzSGTRmziFdAZxYPOxgR/7R1gh6/nTpfUs9/eblC4xXo56YxobeBUnpL
fAtiT9SJOcbMkvIEG1fpeBMrUVqHKqatR+rypeawjPTQzGIVSd3p8//qvypHtLUQ6ZxLys6Rqoqj
RUOi/Chkq+4gSbRPjoJEonh9cm6Cl8vaEm2rvRStwgkfbpejIgsG1u1fEHT/f/A35R7nqetKSHzA
O7qwlf3/LQquG5/tj/dD/lzwQAjxqI58d7IdnLAyZ/GbFF8NRyCYXmNpu0DsoukleXAnta/bx/g1
ruGRgyVZaT7Mbpgq7L584KjUdDax3iPKIOlR0vA0uvTbbPvZAyUV+vk1vmkD+gn+EG26P1gYH/ag
Ao/kHtuvsPrLT9eJCsAzl/cHx3qS7/IYaOvojVhbrNfZ9lpaqOjWrquCbD6Htf3IygyasZtnqFRZ
JCP2Utl1FdI8JFzZLCXraihEgILBI71trLmrrC94P7/MA/8TXUEmJVXMCJTu3B12+505arzixGGb
d9gtQncfLdB71kkCqHM6Ab5SjzYadJLuCAv6ec0BtfACaeBr7O3zHqpwLipHKvKDruzXcF+QImbK
C40OKefnKqCu7OnxNF+PKb8aXM0p7QUzG3etzs2SQiKCSLG3gzb4/PePqo317WFnBwphkk0mWxyu
2YLZa4iPxAh3FXPgsBP47XQSeqfZZmg3RrMe8FTfuaOjA+i0i9mkrmyRVPlRu+YI5LknSJoqwQq9
f6ZIwblug/+YB5k6JS3kagghsJC/DfoEr1pKDkQ+jZw8ddDzOv+LtttNA9IFKk7QJ4edV3KqElcs
muM8hI5crkPt20CaZlRmKgv+lu8hHtmM1urLrAkYP0+Rt11WUSVWjSp48BlcX7lkaUxJ4TjwnqbL
eNaBf//BJO5TKVwtGTawlL9D8ovTSgTyMhFr8/0gLELrS3ndYr1RT/ZBgNbxlY1On2NQX3bfxCPI
Hq+SBm/EHwin3SCDbQqm/ORgiH/Bt55KND8lG0gwatt62pfNDJxkbG9o5aKbL6QE/TCeQUQi15Ju
Fhreh6TFA43Te/ZYbtGuMnjfhi87hz7YXokhKTRvkylPxEbKHUfvaYqjUXCsCMtVAs9p6L/0+IFR
eHi1QDp1367p9WolajCSPL6ud8v+oeynkeRvyTaEa9tPnuR8mFSDdafMHp6d6UJH/9OEULhW3kVN
IEiB5x0tiv2YGlQgscALr3rXtrBNvZxlyIwnFVdM4/vf6S/mju+oH7gtBYO7gPr6yQSqERjeySSQ
C3yq+427XMC3jyVFP5eSdpwyI2XwnXT2Jtj4GXJv3Teo8nGW7P5fpUFseEFGSv2kpvdNrQyj9rbp
5Nss8Umxbl7E9jqbCvuHDcbD8HCpICS7h6lxgl4G2aKs1tkyb+Xk+ClaQ6Bc4p8Xt5VxHYwz8uih
i8Sda4pSa+T27Asi0CJTL13kzrIaFm6T5pQbu40EGuJKf1otU+WwfeWQZ5PEF6R1b5PKLucb9uIk
4oZMkpRANg+jMmKFIPG2cq+djVX8x6fxchS/Fima1reE9qE/oip8fsnCtWs0sdeGXRHVmDttZBal
heAuyPJLvN8BM+MnB0VkN35oGpXd3Fc9i8JSfMKTrKtBgkO9tArvOowYqOQ40f08TlSeDQrSa7dn
VKvLOzdZx14KjeB9nbpyXTxOtIyHhsZv7NauztGqldyflaRd9L/yq1IF6/mWosBHiysgQE6XbumL
poObD+GvQR9QvZlC53uMLXDhm0l/9nik9l3aFd00J5q/dx06+qmyc9eMOm6kBHcl93u/gjw7p96b
qGc8cLRfeiXdDKkKfjYKiZN6pP8Ugq/UuTaa+jPdUj5QjNRyzq5e2/nQFo/PzgnkLGr6N/OdTGNB
siWnH4zl1OX004Pc1Op6ocPIlJsHReXe5XSaAlIRCshUCcPVhdljXXFgRrFVt4CPKYd0kJFg1XTp
/KvHshwPKjVPPrS9PJXnRdZ9KR3E2+HEBQA+n4Z65ME0odgHgZnSbQWJ5wiXxHGAJBeTfWfIs4vD
fRhpEdHnMNYKA7OVGAN/WyjueGy0X7+CUtY8zAd6/VJwDkVMGZSel1wXJ7Yux6qlgnnx7U8QGhJS
Vxf9hmXByEtEXVW08YGqTn4YYGjSqLQhn/Y+Y0qdGXajh9iSXkzuZ/pteffatu2/kYIeAHj/SRtH
oqIFODTeK+OtkRL5nRW+33ZD+RBS45m45PqfUOsLJnCgCcucBceywBgoFU6rJYZxdjV8ACEKfip2
iiOTjIQJkIs8NmAEIBIWlec46+PdH7O5t9+T9wTckVSbkeDIWIZ4hrmMXLqFG6DN+SbKLrlYOeY1
b4PzYnxINY/FimRFoO8FYSUEI5K2Rm93Uc5n29D04tofVkt0jPOPsEoXaTJd2m1mK2tysKo1XZtf
9uWcSi1BArNQ+kgS13GnjCrgvyqv4IkjM2aTAY3imHllRv2/jCemKrSgdYbOLT2n618fWUL+EUA/
ZaRDNVf4uk7I8CWNSxjV8z++oT0NexmtMOYGbugCQUEq8qPKEZhVp5fE6clg21zQTt8Z4QVWPuZm
4tzSY+151UW7C+zIoq7Kd7jOazlmw+GRaw75BIPntd1Sx4O6/x8bUyX9EF1h7afY0ypI7rGV45SB
QSHxTnO6mH3Nm71YPGsJz0YGn90z2BllQ6/TkriLS79ziemnoptk3kum/iZ7p2devhNdMLofGnp8
yC34tzcewoI7VMlxkwXfOIYLU6ZndDvaML2RJPrMHNDPfuKmv7jnlbT1uF7cJvUcGJOr2oo5Cs2u
gJmyL4JRJ8qT3zcl3Si4EIXJ0hkcllxPQKY7IoRNSM4CxnKNzlTcEU0O72m3zaasLtqEFLedssRK
f6bYoY+NFPCwWAyj+hGIf4oBc2w7EMfxdwJj8nm6wPDNygdlANB9cpplO4pQpYS3J9iQfHKk8pBE
/sHltqlfnNOd19TT+2GgadjoHyuI2dJpMatEBMuyQier99T174CFYnsjrS9T+eYl0G6Fzo+9lI33
C6vR8thDayzsu26CSWSg2aHJhwhwGrXUXQWNDT81kCrPc13qUqK26WNleCuF+rUQWuPeabtIQ4PY
1qeK1cBgBAxgAm2d1XdPkbA8W6G5R+zRR6wPLFKmJwROeEySUJQUnyZVWDvLfeh8PB1VL4zDOyZE
U4gjt2o+c42TdyfWk6wzBIQtik1ZuexUw6mrYKy/gHbqHss1IcGWCMSmtqG9pbzFKRaBcjifqbgB
K+RZxIQ7La1NNo9QV3hkyJ5CqhN7O8Lg0kVeZVeSiug5CRJXylA8USN+jKGA83Gr3ciVwrsmVYPy
IB8x3AhGV/QtVqVGO3mmZeXoDGpR/ErA3hDAfx37ipY1SrX9VVEclVBuYUQpJfHqXkgYpW0f5i2v
zrc+WnPstL5BVPcXXJqTUvF3w3YrRCR26LYGXgabag4dtaPR3anGKqgniqwChQMjSjjBQ7QLC3Mc
fb77IWN5Onk3uBuTwLW8NfTsf3MsftMbWf2f7KlF8H/EBdd7pnKomOZJpJFFp/Ys5bS+uLUUT6/B
hjNdatyNF/IUFTrZk0ptxBHFERxKT4IkbfWX7n16i67XGpSsBVcgNYPPTCVHfC/Y5o3cbOKATxkV
U/SN2kXDIiJPMsODoM0aT6ElcmpKgQk99l3M7X0saLQEUDo02HWsBtF57pc5obizuhEoOAJ1tZar
qKlpweywRmgyDT/jAQvB2oGu6Fx9l1fSEqKo6Qf1r1xuOgdQrdO9o6nLTZjrHORdU0MOZCg84uRo
UkOw5sd0oCEMk4ieDbhHEHQKH4HbORZwzovFK5jFKCILNpovLdFe5xDF5ss0jI5ve20xJXLUhZqC
csmM3Y3whiVHF5XTdd5LqId4puXdTAIcnPoVoejTd3k8DMMi82UeXVWWEyO1/eAqedq5mx/yXAWP
9dVX9X3n9FIlXa6Bn1BEPEr4a8L/zI2uswSQ5S73ikGhql1bxPvo9bR2cvOrntZ23pJkEnXuU1pS
8/Swzb9h8cyCncbAL9xoKaNF6IGEMpIZlN3cZgE5vXoYQgyAHNxgtZe+1gJMyA20lk+lZS9creDr
IzJG0TX1seZFKy5vQOnT8WZBoclHwy8/giv4V8v0OrDH2WkO8h/Rasx1GeJCpEzfvXG69vlzu32A
HfLVk2pjSoG1Uiz68DlOQqzT2xuMg+rj2b74JiqsRbh0BpVXxTaWGGowyjt2NdwOtfP0ufHpQ2/3
9ROGrs+ILbWq2MJ28SfOqEwXe5rzxRL4uyQjlbee9R573inEr+atFboexRepUcRU5UV6CtQEYRVW
0rsK4w489l+sl9l+hv59C+mHesK6HPXPcKEC/62N2vFozrYEOnfY6ZMIBE1xA5JO+dVn3pLy2KWI
fwsBWmqqCuQUQD6AdbHimCZV/d3zaYMIgd3lz29PDnGbCMEIgVGRERuRVIMKPqyXjrl9bibalEH+
P0nobNQT8h3skPEayDvYZA4xdWdKE05QFPmfFv5EGFdvutHpIm6Zz+RxhA2yb5pLxhkkVC4bQV2E
hRPXE881Vxb0ga5Q6lNe5A6ozVKOPJ+eUDE0nm/AdM3aclhJ3IXAbSBPNFk4F87xotP4EVR1cFto
PPQrQpIKGYEdTWJPiz+bKXdAaLxOtnuDjScMgTP1Py4FD8HRfH7IzAZLsAQmow9tGcfINI+wnWUs
v2g4bL6kHU0FGL4rpgyy2gWO+wLZSGNYyBnvg1i0LiFGbBK5iN7xemfLB7Timzi0oLrSwoAKn392
5qydcanQkJhLKlpxEBYdVhx77+hJuogWHg+9ISNXEJQF2Txw3tr2U4KnELYvw5lpryTgFWhFUZTu
v/js7dM7MQb5YxhDFhs3doeRppmJDA7CZGO2L4vg0uMzkqqN2rABP+dSTYejyFkssK4EH+3bE/hw
YKK1v9bfvIdV95d3zgbx+ltSWD8J+kZv4HgOAozEvySMTHxXmWqnCKx6snTOr3WjvpL5GesInOjs
7CqTar6x+b3GHC1hGxqwgRmVjFUlzXlQB4jCJmFGtVKfQT/8CLkjxePuxZ6pEJMEwStf+m1PZ5Ik
ye2Ke10+UE6DFgEZssaKgkwKrWFa2huU/esepW4ayk+SeUWonwQPU7KRXk1gC+3x6eFsl7D/bPAI
BMnkWhz1vHmV2Y6Iuvr1XoeFzEqB8HzXEDwvt/crVhLXBKe9DDaZ+GhUCl6UzwkdJCpnnb7OtACX
MjA4VMiO7xtM+jUD/5dqQpnVsEOTJazSqw9UMoNXCGchz2fNmMb1zljxdXyE7KxCczlVP4YiDhzb
wuJVjfRybde/um4l5EIlbQmTJAYFleofWaPm0fRWJrVbVia5SFQ/b+dHGssXITqp9V15PHECvCL2
k6a80cjExmIryLZsx88D/4KFNuh9vaWRQbkdN2/q/0/6MoRPv3gWZ30DejClCZ76pMo9odUzaZtt
ammdEIduJgDW28by6XbyqMSo+XUWyIrDXvFyhl85fRPVbGnk5hKsfGMJkBb1qYtt/wngMDKoc8N0
86jM3Gt0M+Y2tfHk934NO3NrxTwNCmQ67GeBv0aIkXoij2zdXmeO8AhY8f+OPxukb10Fh+qMIs/1
8w9bipYPYXD08fxmrydNpd5K44nuzsCm06tthHlC+2YecCMF9PMUXwrdxYXQOcmDxKdLXJ48wZCQ
UNpSFt27+zkuRozvfuPi/O3d6qpzLqxi/lzE60GKIGp8pFWTPZsu5HB6SaiSlCg+8mnLml52Xe6d
y2+iCBjCSpZjD/UHuMYXm9X+5Klvphc6d9oH6WHWFUZPakoF7b63byH+4JLBw028TDww538We/bB
9bCbQGv0IzJ69f36zrRozQRBgKQNYv3t/ufGw1crwIVyakgInc1kOkOicyy+/TC9wiPfzokuOyPw
BH6PXcRcCW2JgmNqvpngXMiLGssiq0EsFChepFBvefgrWZXSmfJHfF/sQ3H1wUo2UbXITOOEgdUw
zVtFUiDosUs9OlmUjr2vjlFTKAXA42BDo7Rw6vmn3umkx94q0AE7mdkfCfjNnty+MTFjuGZwuhqL
ZgwZnpcA3nrudC5KtFhmMakdE3YEmV0bKHLlZggL+nojRFy9QluP/s12/qp2w3OLqouqEW24SfBK
6RfwmUd3tmvu2guJdK/s4R1MWCOE11i8+bt8FRrSvfDdnG4zpc0M6KVD0IgBGKeU7iTaJSLKNAEz
QfFZf2O7bozpVqymmLOHCVkfLHF1FHWlRXskE0ygbETJMA7tA0BpmSWvVkvHcUNPN3rz6vX9gyIc
kguw74towsvwwPlu96NhsMhN+nvxasjT56OmsU0WmB9XVqWqLX4lM50CVewqZ1/VfEb5MC6DpwTl
60+qrrKlBB9BasPGOmEg8szVGYFnQpIN+Fced+HMHlv5TSYJh8PuHOSE1dSu+KqKZ1TgZMkC7Hw/
aEtDSKH6R7Af6V9DTiDoX9MQ/yXU/aa61g9+3tI68fR5kS9a7ZZI09MANAt/71nU7pCfGNprki3p
aWrb2b/jRcNJmOzrtaQUGsEiXGakPJwC4MIgMvFjxYHFmGm666aZca7OsOfFglapcYrUQGMirnvT
YZkq3K2AsaZMXciITdp5p0bdLpRQiUOQmamUoAn1HZ7InCCSwyruHPbOfJdWfm4nQeK8st8LFRpH
DPegKhNQBzL8LkmBEsE4G9ij0u2ss0W645spnm1stDoQlamSMOzYvzjOYQZaoQ7ucK4YPsULEtID
qjmsNUKMkncRBMHpGQKVI9JqckWEYw78UjwioJuNgYj1qn1Z6J3mrf81K9NdITj6V3R3fsppnums
18obwWzgyM9z/knD35UixNOaSJaKkFKt3vArX9G/zNF0nINjLxhVSioVmbon+zbCh73hciBu1Xts
Ocq3FTvZe/yYJuSDX+qumtwohpvf3mp9uPKPi8LOVWpN4gw7cZyMX3DVgDnvM5woG1hqrdEv2U5c
AnVIvnwc6WHi3p+oDSsbWg0jErsrDoIf6tseA5l/OaA0eX8euE74FLmogin7xu7C+t8O1Y1U/O2Y
1g2XcIkS/xLSlWjYSfDizWaVwkcaIM8v8zLI+8zzwW0FShkVI71KsKJhRi243rrDC0RKo06rUE9J
UaEAm33v37idE0C6UpsD4iRqlfvHPrkrw2brVGTzQAnt+DUm9m2n/N4oNg6zG1gDKwMPyooiMnZX
jDj1tXYnfZ0rqiy8ehxroLjwr3UicVdGnvPv0GOiB1U76DrGKUNJKCGjzYPABsrwHKANkUjV+raj
sORDVnTCmHKJ0dcQO0Q1T0oWKh8EfBypE/3SZMXUKHmF4Z+9D4PxpJNziPFqC0f9WPAB4vtT+44O
LzqcJAUPR4NPcNVeypG2SVmDH74P4n6ENe4y79TmUSickSGi/AMzdYeqnHsoVkU048j1Hutfiyld
+35G/VHdv3qjqJwxVblijEV/UJ4pHv7QdzEH1r5vCXg+FytSjIUdhq8tvxUZFTng6Q/lMP0M+K/F
z4yq1h3zmkPhoHlGXLQvy9n6V/g3f9upY3oZADDOR4FRtq3PeLtMo+1Ooz5uKBUcV6P95FbmJOHQ
oB5TWkk6d9Y37ZWD6JHjpAw3rDxWP79KEvRoeTy+QKoiKlKCXrRjVMaCZdxU7DsnO41DCmdlrDpU
Fgl5lwATiNRVDQ/ewysXkw3OE4HCKeos1SMh5ClGH/ZOGzpX7J5nKnx8DNLYK0iILHYZnR2qrYxp
4BVSsE00KfoyeX69yws7YRnFgcO27SbdlRyyhE45prKKmhYqrJPDDRm43JSUtgZgA34Rnfze4x5w
PLDNLBaIh6fLcCxDi+2Rl6LPVmryIS9kMbovd45MeSFdIyc6xq9zE1I9qrehlrFRg7EzKKXPvhXn
WX7Yz7yfus2eO1/+KhNPkCkn+/yry/2H/eVlO1nrW+9owLwuN3Eo1bfa5/ZamxMprmaq/Zb7cOdi
6IEm7YtciOaYc6Nq4zMKPQ8TlREiEZCWUtH4IMLnEJrw3irR6H5stOH+J0L2NK8D64jESxnpYtRM
cMdGdul9Gi+ZZUaCeYJBKz/O1SY4dzntBDRXPaqtPcO2075mc1tgU6D8XpgY6k4k4OilkOYJLPKl
sj497MCL32x19ctD5KwzgLIG/HHFFVNP0N4DUmmFSo5nVtBCg6BEW0IFAZdzyFzUms7xbv1FFvOo
On/qpBEe7TSovBjiWL6L4chn5/ciHbAYcn9pkqjcvnFqw9ZNSK+csF9Vbqhr1djoMFXT7CUJXpt+
wlaYgKEnnUvEnIqZnciN7vNAiulLa65mtY+2P2xCjUGiQKXg0s0QgqOE691b2skCgyjjud8peKX5
NpBtxQgRuXTuHIzCinGDtRBZ3nrEgHwYpJtIH/2A0lyu0hOasiEGc87ztqTCahFkN+V6Xq0pF6R/
zrcQTMryZvw1ZyB3CgtIT2Qhb5Lu148P/VYBboK8V8DrCoFBT6FBSE9zZqkb8tSmX1gp1aNDJ+hZ
UZI+KLH+XQ1Vg2QqKgeTrAVlz9188JgKTtxUOIPer0jIeNIB9EkP2Qa9xIjY/aQC6clh+ZJQKRi/
n5eOxIh9CDwhrhZT3H7nD1MuJAcmdM08e3pj2v7WPYzye3OV0+Ryxj6nTWP+PwSEB/WGF2DZM62t
2J/r7O1wJFhSwKhxdanNbD1frsoxQtpuNf0hOpr2ZldXZ5Lq/PEmZu/++V197oTgrRWHjJu8U4NA
nCN8BcMntWQf6xJjZdZKS4zn+HBp6nfIPtRWjkj58p/IsUKUI70su7QH64UkIGQ5e+9/xBiJ+C9y
YhfZEKnTEIajf3AAeWaVIc374C8GjydJeFsiFMXTJ/kRWS7XyfvhjbL6S7VEZrnH0VEvoZ+fZwa0
vROHQIZMar+nuFSxFXdDtmTwdvy3qOuwkOU6Mx1eGKzuifVJHcR8O/2252NTZ1tEp/CbBGfOJDuY
ViyYcgtzXOQljP/k/g+fzx0+/QXnNsAIt4DMKGiuTviXjvofZOm3yM55gFP1dlq7RwT0vUpBp8G0
Vu1mqSddym8dnZXP8E3oZZO/miOL+sjBn8yEEKJPUioowneRqLTd4TNqNrINLdq1yDoSx2id6IBZ
NxVXqKQmhoDDTTvikWmwuQ29ogDNfL0Vp/yzbxTdb9XLZ29VioMbPuOSxyi7m1c5AuoPVRtgioQp
ED5MWyraFTObOWSnH//FbPR2TUTyGMBHW64gvV6H+czumOlFM5toyx1wjszkB1c2RydnUgTFPjl2
XbKkndfID7AAlX73vxpDjYEFo3IekiS+l7K81mdWxCSLVFXVSfZDB72d1dpUd5PvNKhtPBjiYwO4
yUdjo11Rkv4JJNliPY2JW11Ni5thUn+DkGi7vHO5zg0Xa9Ceb10BBYcpoN8ePW1S3rHJ9LZYLjnW
XV8+2AMpscf2HkEaCIf3KkXo8JncWIU9FtW1arA3LIT6BrRbUkFVlf46eXVeXOwz174AyqiXZ7ei
I9arNpmX97O2ArsSW2RaCDTdaYtCJ+ExOCdZRVORB2sH1EL0zexeorElv2C5ZH3rjf0bX5ZZ4CB6
tfipVC9k2y5W/WCoX3kx1Ut9zm8242qeFTf7RAnJcR3dlE9FNrOBCOodE9HWKk/1oqusc5pXaUlA
NZbdOjvkRS6dLJpyK9XCBPcnOcWfxvbJQNd/wE8Jzxx4fOle7pC5Mih7zyd/ZB6cDY/Bq/iL9xNv
rn7TYS7C0KroxOiTxE9RnC8MaQ6pseLWF2wYBNyPirgzLcs84IVkcBtS15OypV8dc0FnQsHwG8xR
mmMVdP3tzEWNoKVC2CJu2jhClMd0d+5YIBbnh9rJKhnu3MBL1e+J+0AvCiner8nmNSBRK9bWUbFF
5vps8HG8rCsROrlDbTAe33PIj1xqDypBU2g3HbucWrtg4I8DZ2O+JycPryNbmLkF+pc+B3bd+HnV
9OjZGAwQUjCY532LPyViRBLpo8lygCOgunaASW1HpEidAwJ+pAAsCFppjDk7hYfPgpkWwX3RFnk8
BU9Ps7RWndkpW4Cw+mCGfPqpAkJJFuAecHkZM6f1SEGfeQkHVGf3WnB48O8okh1RJIhr0XQ+JbDk
Y2saBtAKkWcXldVzVOdy7bhX3LkLq8c6gKyP2/yqYUzYiO7gkrSOA5nnj9z+p3hl/9JO61wctdzF
84PR9zecSRYZSsmNp5LfROV6+pwF1EX5nI69Hl60jAhl0CjtJjAaxojGzyiqeF1s1frPO1P19+S2
lJFonGp7Xxts4lnOJhhlo2+tDHDjMzX4k9VcLiq0OYFZNi7rtJ0CX8khu84BLV8ahkTIQnm3vR/t
G+hcoVIf++xpop7yJ3fzpA7JDFv22KCf8WTOg3VjBXnKs48X0CP1wtwd/jgRfn9cZRduTmG+asId
5tD1qfa6TiNJvQwBfE2PXiXXVQJkIVRpnO29Py9BV72Sx4d/NpnuhwI4Kc32F2BVrg7isT15bYil
r1uHSuudcwgwVBwvOf7Jdyz0QUxJe1AtvgRKZHpqOJRt+NSdZg8WmSItQK0TgRqyki83BwkzVFLZ
mobpakr37W9KbLmM9Lngc7/6JIN75gM4dYmm4jZmBDE6HXxDG+eP2vteDOMLeq/nabNu4lsZm0G8
Cj0XnEz98QigZLOX8zmnF+PjclFFjG0KJM+tb2vqaxHuSy80cwccLoCb0fkRyZmHrVmvX+wcqP2k
fem6+xOVx75LR5h2yYQTjjdvdtdQKP+ATA6DzrJrALj1MiMRptVB0/hfQALOJ7LyXsas3PJZFHhz
9ia37+cylZZEVApI8LFzgrlc/ptL+xEIp05PqImvznq9XUokLcqSRvNCP8dJBZjpnjY8J2LfzrjE
o+1mgZ9TjSpUxrJ26Ng9ABiC6whmYnAapr+Xhv1hm6SrFj2iHYe2eRmIgrCgdEaYrpwbeCvMdmbJ
6cgftwhqHz6F7s/6K0DOhfUMgFJx7bSwG+l4Xkn18Wu8FqGNu2I03GOvXLTRvQXqkLL57PVmyTYt
Z5+YRPxgFr2lXBu/kvfxFi4FYFETFxxYm8zeSa8xO47Z4qFZr6lg/J05aZPIzQJwTOnWniK2fCDU
7ZUjuS9XpGj5EXb4oFIV9tvJ+1XEhU+iIacaW7rwgvB0n4cf38UIdU5s8LLtnNGK/aGzDoxRkLfV
62IFT57wIKQ+hLdEBmCiAjNjXLuzeqMYefY3nCJ8nFXHDi3a1ZogwjvoctcTcmSRDpNJtMwet9fJ
kLHzglCpX//7wD/GDtlUnti+Jng6AbGUc3PrOptbsq1wBkqf59UROwd0KrH2JZ8rdL7n9QIrCsoG
ckWo/dkoQBAkt7Cpa5ZXk1ajivahGtZqE0H9uoJ4vlzeS8l09pVUaIDMth6ui5bwGDOmldJkEN5F
v1akDA37QfICvxB/ZAnOONLHZrxExOZXg5qRFOKx9j4RZBmQTXtt+VeStOxWaLS0hI3gis1IReqN
ZTO9vJTU7KT7EfxAvUWf8UQYK6lMRm3wmQUL6A4c2UCpNSOsAhL+iOKfmed3CSAZh3EpBKvkND16
+ofMzyl4ScWnC1Vm9x9PxBtI2IizBmc4RetyIPj+jOXN3FYs5/mXbqKflfxDDQidXva9Cju2NRIN
OyH9tOt+kkUrzFJKgHyZ4OAtcCYh+1bh4tRMoZ2UZJVgYg+TGb9AgHKFgYWxS83eq75ssDTELWP9
nEAcvHdBlOuXsd3qj9mJ1dmD5cvcSiLKPgjCD6PXY/86T9xIbJmyRbhaEfIHAA8L85owitHMtyT0
M/G9qnWa8HLPdLJFIp65ForscxEr8+PW4dMD9f0228iQ53xWycwpXlqKtY77n/daGghyUwzRlps+
0zssJeRblTw++VTdu+WGu6n+gHAmldH3ka0Y/bV1tXUeL3gFJdgm44uwqr4VrKkWXaaefFln93ou
+EICQJcdr/Zo+OMYPhqimpU2w2jijHVYH0KDtWNipf8/4rknSCeiD6O2ELH9WxmdM7ijJ1jBhp4O
6t669vljkZvoeNoUVTyRAH07VxvFqNJz4uWxkYObT3UZOYqWKql0shmWgUJhswWGLo33mXaYZ5uF
VlLkIhAsJbau3QKAuygwQ3eo3tAKTh4iIiSDt++d6jTvj2UuxYyiAP/QPc0pqt8qDQdgSJtg0m/N
v83FcXy9ldn1iNq6mB9K0GAZm/qeh3GdqgqpxcyARpCR0PQeU8NpkjTs61amVJfIp4JcLvpKzatE
FsSfDOijiYbZ5G0iIAklq4B9z7KLPneZnJOiSARVaTKAj2okcf/U/RIyzQfLfLCxWtY5MtDkauvc
2awqI6FYWTu1umXFJxge7aYIoYKciEcTyDdKFzhC8VbqTG3euUM2vmf/C0nAKwEX12V//JVeKYzR
2ahR2yfMZL0sOBqdareAYH3u58eNFS2JWzia8JovQ9i59VkjoeqHfM1ceK4yi2JT01UGCOBH5nk7
X8zg5KCUEprIdZIytQLrKXsALjrOsR4fsORNfGUBL8opPdeCRkXgZV5Ma5XaMJz1SAERMUfFf/Dq
BZcCn0dF7XKA3cuX8dPqEyQPp6E76Q/uOT1ZX8BfhJZriiuMMbN2B45SwoAmxhzJgSVnmDR5qv7M
5X+E+Hk3e7eJ4abkg81Y4hXIKYGgjYzgd1Fo9QRHKaVyvr9Kt/8bwKgryqFJ/xGLDaw/Dn3TULLU
+53ZFyA4frxffi3phnmUtz2HAx8136wfCpFnfZVYloCZG8BjiIQ+waxw4+Q3zW4W6AbpjWlO3dcl
CpuzIWG0PIpHQn2W+SeSDf3teJLg0lyEJFt44DBbDTHipt6v1Iz/Wn0Dg3pSDqXHCPITqAKTZI8A
ms0A3RvnrYnFCpLAgpFDvFBELzl69Wbkd67YKK5JGNJTPXWXo7Q0IGvLdlSwI5DyiQVYCMJ/fe0J
ZaNrqGafSFOJIumpzZAMCazoYe3B0PF2zApnqs4xTxkY9ijg58k3rNvxNXhMlNILE15VASgJsEOt
aUxZKiQYVgBJfWsTKBY40z7oj7c5Qx9ilviovj2vJoaMhfCk/Siw0F8LR0Y7vnV9ilfYy0APq54+
WVUESPfGwKQ6PUAQTXdfZLeoUiZaIBr/spvrTOYmIUr4jvYvcfUq864sXzeu7aXrXoUWpvr9xxMT
g+pQdf1qBbtWausmwy+Qdb69mbee88ZuM/EndyHJ2Hcs+8yjyXBLgx6cRua7v35Ojgah6HcRjebQ
ezEgElzqL2v7At17k5CGbOi9rjJZCTEgcj2r3A7+0h4rrVezu2SImMEHat+hd59j0fdDUX9t57pK
+PslAx+FiPLWvY6TrVY9uf13sZcAnIaeDFkJk7xOAmb7z5bT0fmVEiRBNQG0lDgg0rlgSGP+1Q/5
9yPAS1fV7M5DbLjmtyd+jmQS431AVjKqTI50rYnJCi9iCEyDGQpepp+PrflC3sGEe4x9BTDGw85c
bj85XZd7w4XlJEIZfkzDm7TPK5uMq9llGz6ee2RXNrDRks6+gkeEonq3tzAMIt0YjaIzLR7+/5Vx
GjySf2FPEQt0VAmhJ1hw0+3BreHIEdjGDlDJgfrV9OgAT1ZaQQuudgGUnqJHJjwzCY9gkHniKNDD
Fn2N4Cr+mbuWlbkfRAhVnZvAbavikjIjXPE3pJY6Rx8kLQv+/dWwcQNNhfpr0m9mmyEbJOmBM6ua
X7+JsyQpZ8zHjR4SFIf5alqo9IGTFXqB+c4zUFthus1Y8TgxRw1NsJas0IoE+VNLsAeCquKhv+Ml
NSdQuHcjoKjM+vPcJ8fT/bHtWE7+O+Lm0yrPZp9aQ54an7AOKj3QxkIcpM+OttSPfF54yPSX6tcf
3XtOxQtxRvdUmXPLVlsHL0q/LM8jFONF4NmbZ91F1rNCMQPSycNolc8jL/TIBA9dxDvJ+U4uhpYl
dtVgxdKYUSWaVHXmocU2BLsBGp/n95XRxIGGf2zY2fJAfVy4BDbMADDz0LVFK0DUpWzi6jA+Q8gp
6lpoqkZ+AyzhVBdRPng1kV/MvmPdiExPSCdWKXBrWlLFtrsMSOTvUrBS3BSHFvCPXgM4NAimSMPE
LYQmkplVbeEwQx7icTKFPyjvPR270QEGEn2eiessScIfdUZW5DaUJq31xIMJtO8rirdwrkJcBRFp
blRZMn6RA1rmLXf2VqUwWdMP6WQsJpYoYUA4YPcP62Aih/wmfr3E5B+iOd+i0nvcgIV+ay1WCo//
wi5Fel2B1SjTGn0bBrwHl6dKmwKf+cSOLs+tLDY2GhHF24hL+c0c7BIZC1d7JUPAFkQ4ZD84gwmE
avcV4f+EE5WCM56lFqjLXvYzl5n3Q6tLQiQRM/8tvJOr1bcJj+yCgpgCupVPp3ORtLLb6dIIibEB
+I4B5uT0AjA4z+91bYDOVx1KySRIBl1XOYNRjj+feZBGH2EVLH9lRnXvMN9lOoBI4ng4MaFnD0md
I5ZA52J7v2n4S9DBw1Jmhhc9mkIKMKGqDXu2H+jc+j+SwFR7UdYbkQ90ggv5J6DyuMj7tdsdBfiF
Ax0cpl7VjbR3v4J3QF/ipW3XoiH7iqIAvdqBDHGoRcUn8A3LIjsUrOSeffQxorIyAaMdxEhhpu9E
XhNVXzh5+GvreEsR5X9yVws0BuBr7hwzTMasYaFv0uMwr0+3uRg/wxV6ybCvYY2Rqr8QJhfDPgJC
F8wSvuMRYPOKk4Fd+ZhXylcqbfIyz+8O8wUZhyMO53jl7vUEMY03KO8HSOiaxMYusHAq2PwWORWO
tInZq2A2OG3ADweYF9s1L0QmOyZ1PBBN4yu39xDpFzta8iMyvdRU6UjtkQPi17jg8BgKDgdcwmMA
SsdbQFmfeA+xv/jmZlqQrJ7XyRU6+B/CWpSuzpUcJWxWVJLetZURgj+a9/+qqeVcJ4zX7wN5axhg
+4QT3NGXtN/xYtWpj6Nw9EV4uuw2xABIAzQOpGosf4/nBecvI2R1Gwaj/aXkGKWJc18ChBWPolHF
0oK9D3sZNks74JvjdwQNvsFVSF5VR9Iq8OVxSbLsl/TxKIDKc+SguiKNJqyLCrLGKyge+x8oM6vD
TE325k4btgjcgQJjlhMhA2Q2zHhSpmiHJJvMs4RDz12EqLfBL9K6qyU98eDZUsiWaH9M+LOFZAnb
17qKIyj0SsKopdc7VVYhKGZcYbiWVuiy7jDg9HEcAp13CBnIu43YBUCTMO2FZhd4HVFhofelfvuf
VyYWG1zdleNQxKj5xcWFp6SN75zuaxGd7O1r3YEZC/IFOi3cPb/NZW1ukNhj1dx7Vys+vpVwjh5n
22+SNQ8EcM71RJnFzce36LAJG50uza+KwWUSoBZX7CwZjZatY5IynXolQx+CfpLVm9ljVBeNoOBX
BBIuUf2v/n1d/fIYhJrOxUXkNRW/9d3GTP3JwU0Mo6MXaiiAVMj6VIYRxBsfAcPIsZG2cPZV+wt4
r2zupaUvHbPSox6huBBsmGrS7qgdSL+P5/0BHD5L5okx5HVmWGjZ0havggUKOR8DHazhfIyx35Wp
+25PlqZSXhF4YumO6qfR5ryfQvHKWi1bvsr+tNETvyCVC0Jc+zA+mwO57339bDHeZ4yFvS4DRFQV
9nHPM0XfIpYckRM25WR++PYykPChiVBP+2t14iXGdsdd1Gol3PrO7FmpdUVLTCbzOaAG1eCOnp2e
+JXDDKRVQEh/rh3DkYegc+cnH8QIYLXtIkj1a2Hn7gbjC3RWxn+trmpJhNSSJ8+8oHNPPaL2ATDb
OTfRbj/9iY27OObw6fL9vIU5yCDuFUjj85Z/kv/tWsKq0+1b5Iv1Yzwxa3qDRWCcsfmuzD3118Mw
YuvEtV1/WpNWtSCmYX5dIBRDAN3+6nPZ+srdtazmh+wXmmZTAb+SACfE/fL3JZkR2vGbb58168+F
dwSOcV01V+w3OS7Ga5UZmExSrjEw/YbHbGYmDuJfFX2uY3ghWixcoiZqaQh9RKdSBPitQBlmTd8U
CqIj5iplIxB9qn8E8Iev3RCt9ZcpfbIL9wWVR5IpwRutieD9QDMtycqXDEsZKUlyJa16Y3xwg2CN
UNAA0utwyiSNyeR5Inc1IdnB3LYTU5H5SZVVeBF+Kn0+nXh5tZn5YUehvGC4dhzZj9aKRSjzfraU
U+GsupiFMoxEN3tb0WTBfszw4ASW88rZ3l6HnKugv02OxK8GHBRtvVkMJnxknzxRlw3rj9bcoDwv
Y45oypWGRhVQF/byu0KoWeBW6O9HFVO68nd7cP/2Yf8zRqZ5Mr6zqecvBKZKjyJ8hwNg1Fgu8XY9
Ho9tfzisQaFNgZ52SRWb5hXz+yAYzquWhggkWYLKnf9FlRjU1OSKxozB3Ius7QBCFRb8tL8v6auF
QiLm5PUTZPkAu4hg2ZxCS+wf8KLx2/lfYqLaqk/aRly+6XUmLyruNgLMMCnPL6iVDPA+av6Zlc6I
HBeuhX0apAkxOgpmUMlQiIcY7Sq1XoX2+jrEj7s2ua+20k+cTsOTinspThLbqAQGckcht8vOR3QK
tCERIwRiNnOn7rajsLm5SKwgFrPiOlkp66ldNGafSxeLeDOZIcM/hNFoeJrM+N9ygal6lzDJ0u3B
rA+P3Mwg1GkSGOEwvuI8YBb5flOJ+XSdGVfkiXv61zqiNktUVJpWtFq1Z6iRiN0MkNqzcVFMtQBg
mKNda29WxnG94X5IyteS3Wc0ugH2BQiJ9+AfpwTaQcgE2eJGx+cbqj4UN8xaisNpcM6h1L/O6XDx
335rhAqjdtWZARFxvHnqqMBYg1lWNuvrszSecuh2Jr18aQcldoNtr1cwwBY4vI7h6iBqDXcNhDJC
7zVySR/PV+qQbKUJrxsQPpVCzAHqcID16W/T8zfOTEtxpD+P6jsgvyGdMUM486MLcMxK9Ep0w76w
pxn2O9Jf8bhGpM9UziIThdHCpEIaKLx7kN5t+bLw8SUqqGBlLABxRmmu3OG76rJdMOCT7Z3XItMu
IvHlKwaTjYP3lgx+efK428ZBFlwwmcWr+B7EbVxrrBuBPRw13F+vjpgLgVoIs6HZL8jyqYHmxcjJ
ekjpETiVWWtc7x/tO+ONLfpTeYikI4tkDrFDiWeZWcCI/rpsuU8Hmwslw8vK6weojhoFshp6Ub21
/F/0V7Ki8ikDkgxzh34gWq7cjEGYCWygeK3UDP7mxlj+r+6LLT2ApR1kTAq7fa9PMe3ahR2b6wgQ
+MdDLKqxK8OUaAvOXFbm21lUVC86W4f2H1wRHH127HPZ2ePZe+H8G4djG5WWIjF85pGDU+Zu4kd1
US8vI4OjqtrBWj4EsGAsKnfhwG+zN8EIO33oS1NTKRuETUx4Siz4gLQPxZrYFPWdJp0U94gzMK6/
GJhiyEzvLw+Tq6cJ19o652MJBtLst27k6jDymOoak0yIVa/OGbOD6oYQQaW5KmEbVj65sbhc2F9A
Bv4qO5MEGGTidLhj7MqF+7oPylzL5hYhcr8WTNFjuzF6yXR+c9af4bHyf6nXdtpSfGxzhlZXg4hy
kLi1vTrgtVeT6b6Gc1769LM/6KwSMqgzSgRH4kK1pjqWvWR+RPr/lBaZ3R0yeFdzJTm6mqrXEFvA
/5OUpY4s9qGXXDLpVoFwrPKJWZcePkJp/gfe2HSGTpj7zgYVO42T4FFwpVx1DxPLmQyy8OoA3d7O
bmonjjPO4AIn1OM4SLHamsg7oSjQgifGiHxkwsElEF5RX7LfruoHOMdB18aMKaVv9HZugSWd94WM
I4a5WQODNDu30ARlGT+NIfvXChSdC37/SkmDK6I+Yh0G1skNKH/yDPyhassNwCpFKJYtch3cIybB
ovw7C90l8AkGehy4IloI0/+JIr8gg4PTx2pWCyq4Dv5olRq6FcJtF8DAFv2l6wI/MMkRg7oWMuFM
tejMqK+hMgQCgRJHXpv33QT7w9vMFvKVF4kQaP408nsiOLnPEg7F8f5w1WtN9ylgBLm3LiyBOl5F
6mGlNdB3T2C0LRQ9w/gi9a4UifTwT9vQkNC11IIkR706CgVcIxiAis4vPZno8YNxaxTSFv3cy5rz
i9Wy51vDTA9wijfI1fy9DNl0kn9U+s1q/layT45tFFaqn0WyWJyPkow4+LzP3xneVwYHd+F0YqGT
GlCIdfvmgg11MbOSajAFFh5tZDtYK3/aEJxs1Bb9X7HN0TDJCLrf/O69eooMNf7EkzFfw/EfThgP
9gril7tU2CC3bsVMlQAew9v3C+3ijcgR+UCgOtHI+2LqbpRS8y2CrEA42ouGgl2LT0xxoqeBsGDb
/rIlhv/vIBnbldrJ3pZYdNErSJ5tGZ5FDRs1uPHE0nuy2oMlK3fqAoj8u/wi5dX1G9iU5f+3UCn5
rNtExBolQhPIjc7ApnUhZ2PeOj2TBWf9EJcIAH5MP49OIlbWjGKWfU/hkIpJYDi5D+eqLofqF0Il
OlegIVYZlde01tEClWcannkmD/4fGVwANy1n/edsvE5EcZ7QRBb9jAyJJiy/Zjyey3a+Ti7CQy7R
IyVy1OfcF46Y+tNAmG6bHV0OsW0rEC6xWkkt8exPK3UgM7HwscjB96gRUiAnzfNPSuXTTM9pGUe0
JO2I+dIGtayptmzQ0SAnySkzsYVZQ6TD1IwjJSHgaUsYp5rZluoAzraO8xpvxStj6lAhnriOt+pp
EtHTJYbCbUZV2CydTaUjf1MWXtArE49GcijUucWCQbC14GWNhqI2HiN1ykxlz0q/fTanNj9J0gqJ
p8pJmxARMhuMl1wjtICRNJ+UKemyOLCKKrAi5Q7IqflZqht5VoEu/NkrrIz6ZzOua3scjmjq6T5C
H/ArKvxODvPZGy7ncKoiQb7f1c8F7Xh4p5ibD4MucrGEigq6M3wAnPp2bXjZv927QyCArPw/h/cj
4P1znIvrKWTrLXR3QV1gBo8n5YKJH1+oHFePGnaaZLUGsMJSRv058AUQPWHbmKvdSiDSSWM+G611
NC1uKuLLm5e6QVSsm2tctAko2MrEo67wV9UpfVyU79RWho0Y68g/NS3y+5ZqTEONUAVJfG4IkSJH
loiySr7WbH7mdK5GGSRJXF0HuH3AiaXnQc9ISjM9I95UaGGnYINstkG5bUqtocUqXM8npseWHDKh
p2K0wVjBHdC0EfO3ChWW2ZBHIb9lJzPO0EcIoNrTZwR0pDq8AnYW09c6uEJoJMdCpHX+rZNniqXI
7DSIrh1bOGhuUe3FPvuYZyTaI09y2Q6F5z//so77SJcJRiyNxFj9MZ2BbjtUx10CpLDYRN8h3YNU
2koWYteLnr6oyo9NTdWDZtJIKJIPY/HQ4hsgK0Ba/OWLxn+gRV1ia+Yfc6d0ubetdIrauOGwImTq
xuihXymToDahoaVHssvqV8j3/3QQEchbObZj8FWNtuqukdcIBFot4KlzR/BqFGjJTFjbAiEbjH61
WZE6lkwpchF2yS6P/JXh82w7fJMQgQoqN2SpA8wKpYjiJGgKg1rTAT01E7KrWMhrcUXjOta2365D
QV/4jndBfodP1r+BycAmuIMT7bMLb0HZtNvK2vbDLc0rQsbm35Whmx+1IGXEdOnf7l08ov+hz9S/
AyGqwyOYZdjJvEkfZJFfwSeq0qLL5ulChCB0nJ8ubXiyFVPcIY+Hj9gxNY6o3+9Ax4+WmGQBdA1W
XF88JlMv5PEsJBLOr0nf9Ty0IdaM5GHzYoNvoGtv1vvJ2D7Eohk8FoYFQCG2h1+fcoT2tQOSciYM
w+gcSZPhGjbhcQtxVX6/p0nT1Pk80Tmhm8g1SJ8KBECuU3H+0xByeSIPtFLChiHFg1llUkYFP7Zc
I0KgIKoZZaQdmjPVnl8lO4N7A3g1BSVuEfNfGf9pvaf+TpQC2CblRoQIpeCgarsP1gA4L4DcceTB
7gjSSzIM32KJeio7guE5Q8sBJ9KO6C1aGPYm/nvrCwV6tGC2gNPYLMEGpraGFGbDjDBm+v0JdEnd
Ff5VdD9YKXcxYDl2aug/IMgdH8/PTVI5SyOYjGO6fspY21QMFpbKD2Zqsgj9FFCLUEbpygBLPTW9
KafZlVPuSWIK0LK7kVarpzkXdbiI+Tb55IayCHdZqd2wLsi2N9xzvNuUBYIF7oEc3WrdTC9ifd7j
TvxJFaODQI+4QgN5/PYnExpbZQRmxt28p96mCSycxpBY0CBltHRvbQ4P69AYT7Ek+0ZAFDv5hCcC
RLXc39AYXgtq50aJH/fL2YQ0UEPi8Tz3v9RGSMV1C+q+LE+vjZRGmwFPyrpniu6SO9dNUIwLxax0
OLSMA1oNoloPIf2NBMdCKJOl0lRlgGmVoehU6OruK6EdbVNoTdl7IUmePfPQ2eb/qstuJE2+j4Mp
awP659e1xv/DB6/0lvhTf44kXIPD1Jeoz9RRuRjLhY6PdjrBhMuvJeKowwrvBEGLpchwO38qgsKp
PFBnelZr3BLWdAjH6b12K1GjRRsunBdFipeRjawKJ08mKxpufj3c2BqbmdSwRAGorrBnQaOlpAZN
9hAmb3ZnPfXVUoip4vVnTQFotUwRlW8p315DqFmW72p8FY2DfxW7mrvo63xIkap/+mnLfrNxnKHG
T/ZBaP97B8VbUxU0tkbmg7fIL8dDOcgl7zYhBP9L/PJOj2MbKQ5EtKCgFNRL9JYf7Xwff/tsEog1
+8cAgQY7dsQ5WWk29LZ0iRsOydcsQ6cycKZB+nf6+v08brrcUwVsTM9ZLExjiziHIFwPh5YblYPI
zvAdaqj5lKwbfBKXs/oCUQQwe+Hh5B/uy1bX3aV9fNQf6wghUxcc5UsEoVC+tv7cvD88vlK+eioB
ONfxJrYt944zvs2e39PDN1bayGAGi/bzjzE0spCMrUb76oioVtehFDySHtukXiSlQdP6dqVxnhEX
aEZAN/PUcfff/0VpbglPsepfWKV1+YYXtZiVTN11S7FbxJ8cZaCVOhzu0cL5qhdcvRl5SMJRlOMm
nTRIQrYB+CrsPKd/mtVD55HkdglzDOkHH7xbOK0kDhL4+HFQ69J9FxS03ne2gyUu+PsZ+u6QzfuD
RqQUQbZ0AIfE80ILoOs+n9Dt6W1njC8vNokym4dUbqPS14u3ojepOV3tTRjmlHaSnJ2pAqrhCW0z
HdUwOWlWdBWYe84zTbMBswlKsj00N8dcWWAPHk+E/1k5ECo1I+F9w+1bDZjyKWDMq5ZzrvLLsprp
92P7zsuXuSiBwEpCKbW8YBw2GP20DGqgrDgu3jw7KZIURhJzE1xY4AuVVqA/lqx/Uy0fbKqnv9z9
Pf/MOjYOcSEp6pcmSO21+x/pVIrtptMUsIzhO4BbNo2t7FgvEDjIIrD/WhmbV3uGvV9zHW4DN9Qw
mYcEe+rMKGKvSpANZDzM1/XicS1LZ77EUIxM+xss9iQ8UV2XSlLniL+7JWYSxh2tZJy7EcriFNml
C6nf4ZcNx2wdr9nLlzRbo2bwROPCWiHzaPrMRzUp3T6oh5PFbAMHZ6LOa5HSQS+piUFefx3L0kgZ
tvo5XEmDlCmR5kP+cOveizV+UYZigm2u3/RkqeGmUbNNP1S6ROqs/aywvXru0vzEnzRr1LD2OuVE
wzgJNixUbVE6O9PFOFRJiTlbh4E96h2bYXuMGjzTU/k4OURgLfwnet6sBKe8G7KPL0K8nxVAyyoW
s0fw7YKU/YHN/2gjNvN8chD1HoBcAKX3WZ+uPLctfM2b+AJgXMRJ8X858jAZ4+ZF4hQqrO9b35z3
rQi9HdI+Bd8ZNAwBZORlZteYTfWHX56BSNqIAFotQS+Agmn1fmMHfGtZw03RuG+B89hyQX99jPzI
rUwtDq8onE2xmSTlNTGbUeNcF62DZFeBcGidQv5gahy+IpmW8VwozTz5t3/FNlcB2aGohvMwenz7
9JClSp7Ylh5Ikkui1A68C5xfz1wBIiaetFv8AF0yeXG0ztc+FMzpnPKk4h0PPqO9r61S4lE9cxsU
UaKo70jawCISx7IucJRWuHbkSNp+qNTh/CuPf7WmrjzPpoCnWodaHY0owgN8cMqkxZQzhITIiVqh
/PonkGk3yG8CBGzODN9ymVaLJvBHjcycxSZGQ9fdkJMilW8zVUimLXnhd3ZeezoJkxnjIZC5E1E6
cgmIBiX0TRzi7G3NtHa+JrO87mkEc78MuuigBF+mnxdHv+B0QHp5S1jt7iKkbBLW60fMU9NHiB/y
6P31WJM32M8taK0XfQdR7Glm8mKFuZJfRnJ4V9frDXCNR21z+VCF5Qh32ygkhyrII9BizxaiDmUF
uOYPB8qgrz1tNTAOuXol7nA+0ymKfOlsrD4ynY7tm4nCoiSPnzi3pYpbTNb2Kf7EGOWKZTwbVfTl
QdhVGG9pRg2m6CCJmsuGK1LWuDO+xoJWgKDEDlvccSwTYVK/0pZLjui3RhwcFHvZ/oWEBqudT8ZY
wD0xfiGotQo1ykPpEBV4nYqjWOrF8f4jMyutb6UD6JM1F7L1K1rJL7b39Xs5cxnnbS2G8lYUjZlS
PSUIjfCB3A3H7TRVjolIrDK8DA2RvB4UavFB4D/W34sZ3S+EYE45W41Fbi2hQR/rt+RAyNOiwTPm
kW5Cwah+JzgWi4/7q8pX6N2s/7HEXwjhlzJ1dJz6RR1PzgJxfOISSnQxtghdEFRGOuJJBo+j8kr/
cqa0rrTTovJC8+USWxehksB6ZS7zDqeyDijPl7r8bsEpmhaES88oWf+LaAD+H1SbQWzRGneMcJ1R
1aLbLLHcJaD06xe9KM/eYY3PpvWOeXvvWgCl0vrkdjPSs4+0xJP+EKa2f5B7VpW5aUc6qjnO5JPB
oIE15g/tYc2l9rFKa6L+FGRi/vL7Tn5abiDujAgrj9yv8bubKXMRdS6JLzIzK0IJ63J5qyhetX9T
l7fVLjSRl1M5CiDJrPYnHnblWmpyx7y1mD+mIIXYv0EOvW6MlD8VFrH0KAMr14nHYG0zLrTYHQvE
G77XUY5fHe4ynNSVjaMAQgSfi3vsi5hieKTVUNXQxn/gXEa/1Uk1mAEm1JQoUlvDKCH3zUqLo6dg
s9UC5H0C5HJD1Pr64KaQ0S89lwZOCJM8f5NKH+rC8Jsh3LFE1b8FnorYci/2N+8xlRwocebKiA+U
UQtWGyPcj1PMAvv2GwERUucwGablZfvNjd5DZ8M3A0gOihyhy+WYjwI53bHSaZ6zybYhFsl3NAYE
edojNYU9DK8Nt1/8fA4XQrCHOgB2wguUPaSan12CL+gGTep4YGXPTx+D87oAiqUzihr/5w1xMzNH
KkRlFw5FnJIRghVxVqnF8YKqvMWyLvwJcul+VOURmJXglLYsFRxI5Wx0xGdhcsua0AVOLm2Z6+Zo
p1fNNVc0EiYpmsuGBvXE8kpeuGwpKEHmBr4yBuaEUFY8eG688lw3MGyH+/brrKo4fDSaHQrrBA75
iaiPJ0KyQxpCB96SU3FMYjLYQ5U5aL9MUfBfVpntT5QfleGHHBt4GTYvQrVKA/JoBle2jN25ekHu
L6GeHPdy0FJKerrZYGaxQbl1p/dq7qU//u338EXGHJgM4Wy9s8k8sIZ6ZG0h+dDHyXJ+DD++mpVX
FeQBjA9BllXfyeC+6LEDRToIqIMV1Vue86q6LM+IFjjygWKmZVhF5nSKWH19/PNPdWZzC2Yi7pfo
2Mm7bTzXAOrNTkrgPcKcxETV1dk766gm97R/v1PaqG7ztkI1Hl3DK3SPDpMUXMcZmWSnTzgwV9zr
kV0cNuegbQ5LsZHXYNm1C+mbz4IdEgYrorpHlslIgtcj8A032KdF3xVudG2NVArZ27iTqhbllJ68
Ucs8Ww+kFrp5ev5jwrbFx+GwREjIklnoeFUFv6YDXq/fEXzkLNytY3EV1zUq07jpHlfPPR+so5eg
Fv2TSl3CBg2WTHNvzQM0JeUNuwqHaHC05rx/8z+/57vDFCnAk2etP4+mg5tOYaxKb+FMFV+BKnMf
FW6mP8F1V7vLRCW5sLgghi2rPAA/wjvkti5eUNkEMM3F0IXJr7lUZhwLfT+tcl0bjps4k0qOV5EM
ZQ+9oR90a/MC2IAsxNeODbU/Mo3iAqbKWl5iVYsZao341sZA6wTJSPdRxPjhq9izcErlBsvCPPp/
0V3G80ZyXseQcnZGUp8h7SPxNojmnWWX8AoNNAc0LPxtheIS8bDGUJwurx7kE3czsUc8e13wBMEK
fS0TZjYfQsADtaJIkBYp67uv7oOBEiSwd8+3AS8jywXYIhvePdGCLxI4Nj/wo3kZgv15J+OvLpYJ
D9nYITk7e04bB4+4d9+ChMwvlcIcxJmCH9khXgEL+oe3bxxm1zBdWJ5CW0yZR2X3SSgMMl5cqIbn
iPEFW4WA58nM3i8a/jEg6rfTjIRvGjlWzakn5eQKwvIzOLvO5CmqDzLPxuCxjuQIzw94nJGI5si+
BWbJhaPtkkvQ9P9Gbk8+LwJDo7qLtQrSky6QEllKaFJseL0BhoEUDoycMY7xUZmCTNe+L0BeuLcx
8o0aWXHyttfXjTc0LkfiQIdBoyFrztLF/fJe93BaLmqMlOz0jsdRwNgYZWv7UIu62067Yrf988sA
76ztng9CzSTp34yxkkIYIntKQeXToxXlB4zKqmWHseYjpsaIOMB1u18+ZgnKzsUbmFtU6UCFYirX
eYlHl7fdMOUR2k7KbxDXUcNT3ZwfnBbIr6euGSdkLFgAQlvrTi7cGFBWEQmhZSq8Ggd9CeG/a/ma
Nf03Bbwn+CGF6XN9SUf/qYrnakyjhLgk4d++m4aYALia4836eBdqybKSh58pPUz/qaJ3jFeFz1KX
y9jBTi6QF8rbOnz5SZ29O3XRM9m18h+2w7EvSsowmEKFgsujG4+wWuLAHApcZ7N4MfuFvtFECwhs
xGMCrmEhBGGNm36RsNcbrd5HguErdZ75UTvQdkjsI+YHOBC5/LptbDJWruUe/s98eGJgBqromWKE
cUemmdZPZ6PAAZijcG4xwjIszGRGcKDAt44YiVHpRAUT5xAT/fTMbONWLJCiuxmGPIY9vVwod953
kGvI0wdUi/jsMpDe24p46oCWZNNp4E9TG4Q46DWiJEiMTJWzusAdFfk5/LwyKLpiI3Pfuzz0KeTS
Z9S03PYBZ+NYF+l6+UPLiw2/loMu7DQ6eS+R8bnWY3C/n0eh2uxAXpU9AKtV0Kfqnfk0fypFdbOu
vVMRntv62wDBq+QXwpiB4d58Ik6g72BrqJAYP7Y1OjhGelm154/wul2SdIkwo5I5J1rxoPFP8ZCH
neQI6v9n4LpbSoNdaGB5sq41AHgbYW9Dg6jFIQk3E8ZS2P/62Dnipv9j3uuGQWY+mHgnsfrlINsC
NypSu9nowu0RvGzAb42FRaQrsn2fuMzcObRgowf7R+Eawb8lMNAakBZifUd9a5qMMgWpbZHkL5G1
Wed9U6adE8/DyIUSWfi5sBsH6yXDYil4oasxOJXWLeiL9jbWtS7q2dlW4LklusynNSqR3XFoDbKM
rdVg+Cc5cjzNjVgVNK8H4NiSt4FGw0ITSen6HYVuErKoIwgBPZEAomJBuEM8V5NmzCojYpDzrZEK
yTaQ0uwlscmBFw34Hvw9+k3oqf+5cVjFmumoQvlQb08TztQ9kcGKZAxmTrxwH5nHbFQj8K1Y/g98
1QnPJ1RS2JgybL0Cwv9FeU2OLQkpXl3hONIaFnX5eYin21tf8rHFKtHZMRe6wbVpNB1aQhQyQpes
xAp5F3+pMW4VG2nrna5Y7fh4QMvKpzlxfdoFPFD8qqwiM76kgE0V0NDqflW8h48mtygfkaeBaxDz
AKknVmLT00xLDpfnvk4xjhXJMpHS0nliSfk/qZ0HwHNv3jtEj+wYzIDlQ1sFMLi9O8trDRmk0Opb
U60UXrbYs5/1pet1CekwszeeoUOYW0HYlMotXc2qY7HNmyZiSPPqZwEXm1awTJvZpCQpl7iC6yiE
HvecmQ77lk1Yrl6bFb3Pkz+HxAHabMN0zvPelnWIURhh/9IwtJt9+4kCkRxnNeyBeX1zY0KicngN
QKnYj5eXtPJwZJA0nlvS/L+8nvBFYIGBZfY0wM+efA1IG2EjULVEDmJ8YO9jhNlOcCO5WNX7tQH8
brs5PkHBoltFPUW0pv9kxYg3xL6lPiDzQLr3rTbG3XK/BE4hFhkOpxvLjiZtg+tuUIVgTeZvmhjX
+38bewc5ZQkfE/XkdtJz5u3ezc+R62fd5P1gkO0kABUvOR+onPfwEJayWT0gx/ujpub3vAM5kbQS
7wSbfZCv81MU8Bsxv0ltQJnvHtDLvj+bdYUi35rsF6zZBOVHEYvHsBa4VNh6l1KRaK370vSq1UV7
Xt9iUti38aJorEVXCPZHPE2fFnTHBHvATOM5m6Mj81WPMNQ66IB/cnaocAnaOxZGsSTVJ9tOhodZ
S2llVfWQEUCGDNYwNFoH5+6S4MJCZ1h0OAByj1pW9HUjnCBkkAretfvMZp+taVuPzMe2ebZG9ij+
VBdVaEMzNmQX0+5WOpH1pSbaRwoXfaP0o8zfqWWZA9ay9z6Nr2oUalVxtQEME7+4C/TcnuD1Hymq
42k8ORbuvfzDbogQIcqqCd+/WwtpMr3YZTLgmOuN1XA8piVOclvWo7JJ1RMCT+nBtRCSXtxTrDVK
4Kx6x+gKcByW/yvZ2XL5Y8LTsNoubc140GSuj9GHzVnXLHaGvlCIMNuHJgf/Rxz6pzzcVYD7R+UQ
2TkCskeBWy/ajJn9YHi1I/sx1VOW4OU9VPx+BmJp6E+GWhoOPjbzMoYX1jaExPwuvWJJC3IhAHYK
/DG4qJst3C7Sipolg0ezQ/AyPutSRYjrPHIaPU4ckxysgde7S4a6tdc89yX6epbYkrA7/gIPvpWL
WvAaLtnrGzgdwP9fLeVgQA5QqtcaWs9WQftloWmRStc07GNutqlMAVsg+BGcFRcH9NamgOzCqW/v
uuji7q/stdmztHfgDI03DVlAl5QjteazL90DIFZBc0ABjvYC2WVDc5fhz5DgDnOP7c9HSrN/8T3n
XVSVyIp1+Om7H+B6Q8QyxUI6kE5wZkfaFTKPrGcSNO79feRayR73nqm1kUM16lO1uKkjJzoq/RUb
SdCYbkkT6k+M3HqAF2086HGaRyoUwyPK9WoViIMLK4v3lOuc9a0VAZA9JvpWMez9C33kzs00ApOQ
oTnfbgcYjFiZvMPjxNxdW0LxqxpZkVSf5XqGJr8xMDmHRUyoPISv/qJgJzk5nJ2f6N/wh9hloq/u
xDwVH4MsTgBcL318BO/ago8KRyIPlvu321QFo8VTiX07AF3NrYSQMCSu1Qzypv0/c8l8HZ6YRu9Z
TxDQnKaipnNvs5FyqX5CYFt2yR438PiFjSfSirOjCII2FQDEBavGazEc5vGegjSpjGw3ruSbvMPS
+cACRBAGEb54WIPNk3O5na54rFyuOjrNowcTEQ/S3ZUmlSrREJAT0jjmfxfSwvbUP129duTxAZgy
3iP7zBn51yMpuKx/17Ch+AVPClKQKzoJbl17pd5/EZS7K9pKn5Sj8++SqzG2T5Q65MmbZV3Dpmn5
x0TFVC/Yvr75ASEgqMo92K2ecGGtdWsioIi43M5OELHko5Rfp7DEhudrpRD5BHSqwAYxsX30VcWJ
M5pk8C0VQaqK+x3lun9H00XABJ8u5o4j0vlHQtK2jCZ/BXHtTJ/jEk0wUR8TxtFYqu3Z1iwStDcb
wzfbIqdfQWfhXM7r4zj0PNHkqcAfIy1WatIB63A7/Jne1DOCqsmdtTqbOx+SwLk2KUxhGfY7ye5N
kDgxvVFyDt/k1kBJcx49oGAlcUErSCPXJukTPcpSypLZs3TQsMWj+LZIoZFyr6JfMjFF/+xwAuzj
/dtL5Py8CnYfgIDnrGYh1wxjo54FatsuhjDLFfDbvkFq0aFQXa/h1sixcpnd3YKdqGwPPZ+Sizj0
aDHMwtWpngUNRM19Z6kY2oUijnX0htEZL/zR8RnrKjyFBUR43YqZN3dAEIgOs2o6kOX62/U0GjwG
TVHsc99DYjQ6Ezm6TWQQlppPTWIXrdJda6criZItlc2wKMgti5i1zSBLTbgugfQcmq5rdlD1Dd02
hZ0C7a+Ow2z8Hz12vjTIsXyiJ6u0g6njm49BRnqKvgnJzdsip8LVmrywMOmcRUkSSpm1dE6IDtTd
t70mWhm1cPaQNq39hgfUvEKJvJRpalpkyMjcsU7HrNltsFmDYtkFVCQXVuvqH8VuFBfUgGvwa0fE
LBJZTRU68/dvypXXcXY76ifytnzGqeHeT1rZWd7p5Mj18FSCB0Aa8on0ytm2ax370CslI35aFBjS
tQl3l1pt6dzvJIbj7nUxYbdyT7HRaSkgybMko/Lr99XtC6n6+PZqi25xXI81EhCkFi1oZPYUbHsW
lbKqe6yOUVboGs2oGtQhkaGNkQmCjxs0NUhK/BuPgjC5xESg3KIVPDa56OCA9ZEYf9OUutUmtrT6
owfOVmq2qOLBV6MdUZCDYs6Fy/OAiGeNx5ePbzEWTMtw0hVdgvI/So0dBI4DftJkc7cMtA4y94ql
B8b4/mbHCrvEn8sCGmI15OrLe2v9tZds9bO1xGKuM9T08CM64V8Ju7fOGfMnFZTvYMI1+W4GgYoA
acNHmJlyuK/dk7KbtCi7AreFQ9XF1cKitH7gzQgIueOzIkCNiUlFk3pCDPnjz92q/npGKHmEqf3Y
25h8C04ebZ7hsS7rZhTaqYpG840sZSymLK6XPnJjrTX0xPokR3OMkU/RnKrEOtayEx0gUyZ6wp7J
vGs6eirF9u1AOpZLR8EUkRUQ+GXwIpZgT3udjKdZ+to50aBQxONgzWttEh4scAKldENQ5epT4lha
KcEufYg/AunzET1oz+KZxiKM0VNHdyTBC8s91tizN1sRt8H5BXwmVY8FpTUHUcJH8MqqE5nLlkRG
9Jh1QOOK9cXfvtIVWzxxOJdL7R7WywP3oNj9RHDoDO3BTsUluJI0jFfhuQQge1dTHw8LLgjAtrZZ
VjohY7fUNl7uxA0R4M+GNXO2gEzIhvZiBWGYdNsiSrA3YDrTyNm3loYZbAodCEhFYBFD63BWWTl1
/CgbvzpeZT7zNMq9HDYLOavPK6myfER0EipFW6WzVMYXC5vrZ0FW9O50oF267JpZxZCHHaX1I93u
DYwRUV+Eb0K3NVOuQehikJ2fTMUhd8YcA6i4MPNcJzBRgIvuSiJHi6MO8lAzFwndMLabzunNnJLn
np4LNmCM8hTEL2flmtEGs2wOv93OAaDO7xjpGbcl8NyupPbdQYbJ0lhr7xdGjc0H9hWFTpTW0eMM
F9YmaLvInpk7G6QvaVXd1noFOGKls0gbtJv+4KZgI0PW8P8ASGIaCtJhP7JqAw0qzglSZORwsJgR
z7WM4Nu1FOPquAamQctw5VM6pz63uSX/IV6vjfF4VPuXHXgCwO2Hp5rhOCY4tMSORDNf2E6YlQbK
zD/xD3s8mWH95OFZ2eNpmOHCRerVskhCaBLdQB4AlsIHMd+xyy3jCzGYBij0wvHiYauFTB+nMe6v
WGKXDE9k9ePoY5inPc/XqKntqgJLbEQBjXmUIO+yVuvgnVwZfxfpX/xXaZDMwT6ql+20cOGxCOul
zMEP69b7+yHHkewEeFiW9a0DY1mE1kkNYBWgH5qhbFzyp0lg+mHlXG68BTil1sf2XUFQrE+i6hIT
mGYkzk/2Z1pF2ZA9CtBj66HG1fjNxxkawWzH0/u66pfN43iLIaOtKErYs4T8MVxCnwALbTdIiYvD
umSgvclQ5EJJpPBxwGJ/fYJAaL9kFnBa2Z8e1aUNM8b4nYGtzVWnjpI1lamYjAilHdafPs81TM9z
cKtrQbWL5c+ZtCZ7s2bNZH/fMQXQBaXVttJbFKS6CUhRLAoI520JtIFYCYCmpgdCzovpOcFuSoj4
jN26LjRw8DZWF3YNlMrlcUk4BfBYOhW8y+akbwESzMjl4AlH3kZhjgsLn1I9f/9ndgqJIlnTCaSX
g4ifGUjwNVZ5d7EKCQmnACwis4pSgJjnO52WneExAfNOGDjG4QMmHqtCdBqe3w8Qz04BWDMm8ggM
5TiUBE8QJhoVcibIAiEUr8z/w5C4oltsKp451IAnvGkiadwhklO0AfiKdLSq/2xs0HCwW51HHWFV
42Egz6Usv/sOphQTvBnth89m6eWiML9Vb5PiJmU14al0vPBL+BYgyplQt6w0Hf+1vgZmkLBNst+6
gGzhiyKA1r4ZdJ9iaitJZHq2N/sCyLgO5Otcjek7ILaA7oC6bIZIs6Nc52YOI/SKoudqB5irMbfG
l4bea4cf35wUoul+Vhjyk/pOtygmXPwy6q+ch/A4+z1A/KVPP18MraER6d6APkKFIN7pEIXusawy
lPXH3/bPbh4+kuKS7vqI6C2KlNi9GBhB+fF6iqXEbkMwR1tEBWAyNmn45ZMkmcoTpiFL7VbuzmXo
6XtdB7+RmScxfO3G/GaG2xBIOjDZSdZctEg0GwuflYt4XP1FFsC6JhLOYyGAk7Y/agOjaC3sz6al
6wxMHQAP0nvhI/uu0+64QMQvHFm8Dps7bpNCA4Jf2iClTYEd9WWyD4Ym2hcJJMBJd6uVV4J2RwHv
qBTGONy8jP4aHDk3yVOyphbcThFjJf6N5BpdwfUvinsOZ7AMNd83omyGNrqsD/+wg1nXaxtiRnBO
2rFwFudMbJjfZH1CnDDa3ngXxZfR8SrQJBYFCeB7PS2OddSpHo842XcnbOoNXB94G6uh4rnQDFKV
3GWZM7w/Nwlwlq+LzIS1Mne9zOFVdFjrn3Kjryxxq8pLwc+vnyvVD6svRgpaDmefTNLIQGjZp2fv
lHJ1Zbr35yr2b1hogf+VLrXHCOjPLRudVJBVYarohxsp6s0VvWf5JJychAQtGTLZZbw0v6lzlPo4
4ff5Q8PAMYqYxN73pZ2cmCNj6fsGagNJ6vz1cg0esiG4iixOfpoBnIyEfZSYnY/QbCUQqutFI7q6
gi0l6lB8axI0ulAVfvg4kxcpBoQDQ5B+Nn94+3eRV6tsFi1IgajJo5QER7obqOrkepBkbmIMxWJg
b4WOH2NN7Df8JTPPs0n97oUaaYQaCeVRFSWTB1umVUCUzrsa26DVs92I+X6/r2zWDxa2+h7BBASW
ecxImOCkgj77LzY7kQ0/y57o+1Zen/IrdlYTc0G/NYhHuod93xIdVMU7Id3sjc8J8R2txshnDto8
0TuHVqI+DbgQc/GPuT42nD2axbJeD3jVnRMoMA+fUcw13RGGZBlVUm0p1JZ1TunYKBX41mmQ8x7J
LaF3imEeApeVTlHFaFOd0q0ZVqWrNy2hEkukngfqbVct7wEtrDslzvUsXM7UKwbbaiX/O3Ad8fW6
oKGbXtpvHjmoxN8PjNxvjVfn3fbT8pCbmb0bZa5bRTADemGKfXebnbxBZNL4t+QFt9jTcAdXHO1I
zkdk+p1A52wRWd/BDR3gpFsxjMtWf9xm+dXG0TZTYcSjQmavfifZ+BUkj4VpUTRXxPWDx6nKbL/a
F7TdolriHVkL8klPywwl0WVyN9/chZzc5MDY+XRPSU61Ll5xXRRQ43JmzZBXdHPPk4jB8cLHvY+c
rnfB/hIusHoB8MGpM97Kty4Sizdt4Eu5S1G0AF6Eh+48/jJkOJ++8sk0ryDYTMx0R54ELjo7dKfc
7VgjBnjWlgEORv1+KSZU+Z0qUpyHuyHbWZZcb7h7xWFbmhVHocUBHgag4GqEKugcLqqN3dToHqeT
wzxIoyWqFxoxTB0PoC5O7uWbeci6EagNNaDx31VPpmAAyn9OX39Rl2uj1k700xytTctZDthkTmFE
n69v8wFeDzCzRyNDDZz7B/BsyF8B4hn2pADfa0sSXB3vAdORDoOsmbTAoMZgewHwDi5Ytk0Iqw40
oSM3L1xEY7kqsHWqbCTVDOKNdRHqL21o1vlTEcmsZ164TXi1eapOkD3DDMg6ZwShoT3cxF8TAfgY
8+0RRk4E3NmXQ828gQuNSDNONLbcXrUn0QS8sx+rlz/UbqSHTzbX3wHoFfhFZnnU22pw8GSyleni
ssz1SoJUVVQD52vvDNxPjO0ck51QbiR5B4SyJvIbEK7q0Y1kTnY2EIXLK50GqMFbBYES7er3fN2/
+i3IECb4yq4Q6/k7aR880soiY8dn/iVu5R3nR/SMGM9a1TnC6KVFzHprBfz6aV7QkvV4eWqi3kz+
Y4X8t/S+DKX5BpKJ/wW+SXwbLTnUlxFbMYDjoetpXExNS6YgvoL2Nh1So98xNPP0gQTCYy3LAerd
KWK/PkUfMBvmL2ziD7eNffRxrtPzfaT4uQodvCBreX4OBZfgwLZy5gylT8HJyl99zu0eP6Qf+uCN
kBuaK67LDBUJ7EJmwDAGbWXbaKh8blwcQOT2CkIY56Vfzd0OUAHwRyjXcT06MeQz0/RONFiGd2n8
jaA7gUqOSIbvQGc7yvfzJK5VPkv37G1sUCHymn6n4DNiEE+5skfmObKORglNPtOlmZ1lAJHOflVT
CkQZjuP2OD6GP6+qzDCnzJnTlLsMLmQi6AF+PRoezmvfh158KcAiV/bisVI6DTRef3ecqRtfjPh1
zOBl2bsU7zLZC9nagEeMRtXVUZv1L8n81+Q4Xs/Koy/WVBUTfPDs1Xb0+fJlgDztMvNkgpg9IwUp
eZtSbuFrVSSE4OKAVIn+/pvjOtJPMmhXrS9GGPP3h2lkVWBs04NV8Rpm9HMHzTUINQnTnnCu9LUm
yVMXNnKN49+j8NVdTL2c3TaEDvUmDf58ah23xaOYFwt0BhOEjCUQp6S5+ulgbxkYuURH7RKD3J+k
DL9ZGz38Hl1ioHaZXAvVh9G8Eec06k9kX54F84FLvAqrzjbcWcvFWYt+CHoRv8Vb58P+NBHkOCQd
hMier8FHczZyrZL2TS08DtvRQ5YqzEGop9v6c47sgzTtwDZtcrOZL6md9SU9DnIcjJT/bIXdh3pO
pSkzx/GYnYIxvH5eRR4Q2v85XFQw+vXeoutCxWFQH5Oj2bWikrNhKNaLgIQYGnruzZUWDTS7bl7k
vUumxR2lIoodMhDazn3SJVAzFFFhfP+lCw+OMbjJ2RA+/pDsaGLnfYZpr2wCTtO0TO6moKbkvGlv
QhwE9ua8yhNykzZ1jYrYy9XhzzWVBNHpebKJxpey+BWY6ajTGT9HTctlUAn0r8PU9EGntdEzhtth
3aCnJaP7ir6gqzyFUdK4UCCzR+PwK3JQYoA2F7zJRfvsrIcsXJCH253jZwhxFo4KhHGzcEgfFQw7
0MwxtB+JOoa2NfPaFgkL/UYSHPi+py2G261IweLrT0YhsaYj25MvHIoJAHWo16e95j0+VMiJHz/H
4qvpwyVnH08S61UKBi1Nb3o8Wo/GNygw1+RQ8eUp9mnMCuJARWusQUdo4FQutZJzV3VPG9EzVd5W
soZA73FLgCHBLn18wF8e2+Q1MY6HAynoi3BJeGlQEgGPZisadLkqeEZci4uqkfu7Swro+piyow/6
fqFnTgGbngEsnPnL/PqhYC0ogvFlJSKzJAa3OFbe/JuQSMUksPNMC5Jem5z5uLJwBOVVNuIt8lzs
ZXUWYyEP5zzFWlnTaPw6mmw4f7JwQ13FWpUpfEl8fc1BESdoZXAECcKsJNNc5G4w54rsJ2gf/PPf
SLoZAKkwDXDteV0N4Hyacauz4bx7HsA56n8rI5PnyfvsInNsA6DU2jv3ctms5JWRFH3BThsM+8Fw
FcIOqENTLACCiE7qr/pbxQ5QFZwBmq9rHfdsx+LVUjmLmATl3A+r5DD6HwKqt7KlYwzoODYzxi+A
i3zM0FdvzHerC4hKP2CHpRhW7yE7jIlAcg+oAdxPa/QaszZTuSng5Bkmp2FZKRg0XuLmY1TS7e5+
E0ec9uRkd0gZ5F6F1ivisWWPSYDd2HWi/IpJvr4uATRPHLQCOHYbKI9qaSx/Os8woPaVlmTsgit2
KxXqA5gEMU4sqehIq+j844igUiJT17iITQ6DUPOlp/moSi3IUb/p4lvckEXrsKJ+EuPiXsMCVIGx
jjkT1haFaK+TIFHpM7e73RdNLZcMPGgdbPVRMXwYRcA+//iDpFiT3gRbCMQ1xYkW01tdpG36rkzC
eIIKBFZxd5dN9g4EDD7+6bHZko7W7nic8OJrlibUDyG6fr+lJW9DgFivEsFNAqqoQcMdj+cc6QoE
IoERDAybA8154Ke/1UAfwy3OUbc1+e7YeOdFrsWFhXOm2X2N+cV1cyo9VSJwDv3vnAorBAzpgpyY
WpEj7CRT9HeOIHVpvJoQuzrd/wwprGbFvkgbVoPxKyAe/dFJcQngyoq5fELz4jQtN4x6YKLJK5Zr
FlRUKhp1O3ABnOB+k3D5DYgaA/1ZEDUSa0gfAaWfOKfrTQwM8UawtGOoJGJ10mimI+zb1EhMdSyH
lE314BOExjfCs6Et5fQ2+HY9NRT9ci4p35vI/WlOU5vHvVnJHtUU1tVJEfjfovQlOO1kylsEuNEI
PExLGwvbo+a0ZT3dGlePthpB23m4yBHevQZ+Zei0lv5QAfLXe/CMST7vXEa5iIdfWckexPRqW/rr
VP+u41VprXI/RObuZ3PumNMhsaKL+PckDj72RsmrN1tVhoMGLzajWVKKKPZzznXUlzgKS3MrQ0Yv
uTw32u3quSWnRiuRdbnah+/dBSlUfgjUv987ftUPYQr7OSCIYPJluesxXEYdTggTgBL7nitwZv7V
aHtbqZ3APoFirXcwT6+hfLLLHJmzeNHnQhn0pOmfz8bMesOZYP29R3CaDIIfWzQQeVemq8zgW2qB
TKo+7tURVcabmX7bjIeUaEVgUK7devdf/a/JyzXCZbgu1uzCGmXG2bqQ0JThx8wOczvU+D75KhuI
6pVTJStAYy7FFj7J8pHwh9cR7DwHBVQuPtZS3DU69Jl7I4x2djpY0LdHJGUv70HY2PegttqQhj7A
OcWTShbT+amer/7WphnkaajT4qeGpe+/Ixfig8x98eQqTZwCM/U2+7ny/3WQl/Jn6N+RZxDSLycB
X8wCqfRBAfWB5hub36q5RxFOcLefwhCkQoE+TxIoacG+tQ1GGlbFKNjhW1XhtLKEKKH5iEA5HyoH
Z4ud88lQ5EnUwGmTYmuz1epm6V77+uDJq+nMdmrobjU0IjhXMILuIUBumMnGf7wBMXLOiwwlu1dC
+EWv7dzPpSsEpY7aVcxSRvybzLp+Rjqq0UfcH9j0QEGLUdUu3syaGL8Jy1E7JjEZMuXOGanOMlDf
RvVZHQy7p8obEj4s4YPOZn6bvuSEhoQC6slo2p2F6YGBlaNaqi3Nx4VvyjQ0h5MLWGa87ITh4dva
VCDKnE5PzZLSRtproGY64JODl/axbYlgATzoEWS44UVdLNzGkAetJD5lSjTTalmJu8lEJo0LbU+Z
I30L3q7k0w0ebmdME4MUBg3VVsXZBaE8GlnKSl+Pc3XJEFGgNCYQms9WzaluSqtL1iLeeXqyh0Xh
wc0DnBlcqZxmBIIW8GAkCCNRVRoDFkidSUZVw+j11FVpsnNQFae7GRvX8WdymJaULp1GXBiIFUpy
fPMyJDF1LBvBvL8MWTbOSoiF//WUGyTBJ82JTz/jDRiR7oAlZyevZ6eb+PVBoCoTD4EzA7j1NOhn
180CVNXnjEe8RTSruzNP/W25dzaTNtBSQxqY3QOv/fKE41+cYJagAwDhEnpfRbbrjd5zYO1FD9mO
blahtf6mmE8hNvnFbIGvXibVGMSNZ0ty8gUPzJvMa7wSVmhsmM0k07o7VMbPNvvdK9Q+b9VUnDi6
75clvN3B74fNM3Kgq8oGT+wZ1EfSgflzXJBofX6BIY3ZLomsQnyfPZhJNWqGtaloq2LZ/KeSp/KW
4TltPWx5QR/E5ochYiXdKaRYTxGuUXWdmTdYOm41+rmn7EDTCSUmFOJGcG7e1mgeYyhTmly17JeH
FT+PHg4iBQVINaUy9ZMVP1TTGJru5aE0FLthLr1JQBzeerXq1Bk/O+kRFDGiF376IaC3+y5MHjP1
N+rOMVFURPBwWvZ+8HfLX3IrMncQXTTTkhwDZSGoKcFFi0O4bAXOzHq1zv1QpEG62M+ppgj44Cel
AYDFaRpYYd029D9Uo7Dc9n7chOf9U8Ev/oBf7lja+a8fFRbSL8nGkGpG59ipDm7FMbASlsy0Sq28
Jf9jKByVUajRPAoXaqqRSMIu2jvCFL84CIEjTCyxmbJhbdVF2B18opx8Wd6SHnTTx90YIU5uVKjF
F8wr5J9uU4N8ZEx1ZNfAJUjYc84fcQpWdGIXf4tRrc1SqSGVocjDX2JdWG+xj6JRpnTSwcgQdtIl
Yy1zRlk21EktUNU8wf2Nc4C7kWi2i4YYOOBLaaXNl4U4DEecHVKwhuDoDWrxfMaf9xQFn0931ErV
Vi6R7beO9jbuTXwKH4E1vyduT+eibEfV3+CCGmIKHxwGKeEJwHdtBxrhitbqf/dJ15uu86WJTpBE
S88Kz/vNA0nSEDqOIJHm6PdAdVc+v1AEDINCXghxJxfZmSxuYR7qCapWzaPN2j5z8fhRHZEA7aar
XTXUukLvY/26gUbj3u58b8YWYepQLVcXL6EW6Ji0hD0BRFwXREuogdBisqYSIwuRcunlpcoLffPp
c7mQH9LYKOCaovMMbx2Xl7KtFlnlEfDnj+zBV6MANUyTKvWewJ/lAMeprjupxX+ov+TvR0eq/sS1
MGrXqRpRXDzjhF/6izm777SMswoyPTpJZm76aacDt/6NnqC2W9nZ+KqBCaUfpz5NIlx3J3qoUrT/
iOf40C0IkQHmTlb+v8dBdAqr8gHIGmdXWfRqmzW1uGWOVZTwkizdx9wgsbuBghkPK2wVthD3wBi4
EsYX6wS6aqV/ELt3kOFOhya53MrB76dyBaRXK+MzxOlTqJUQr1CNTSWUBm0gjpL9HW29LkB0MDO8
080E374luPEgt42IHUglS6mL9YJew6jJqM/ke/OstIVkdJXV3qKJ6y8nfd1ro0G4r9S8lMLDeqdd
IHScGOOT2RRL4JxbgyD+95r5cv2aho8K1XnMWgdV7dKXn7jKadK24kfCaHoUp6d91AfGny8quhxp
s2xbcKzDphRxWDilHw2PpqjOn6w7jUo0+sx2J0MsqJAT8BmZz8HY60Srw9ylIj1NoHkXi/ip9Ps3
D7GynLJnyEZeeJfhljPtlo98tcfqXFlomMlDeNirPgpdzxpKwzBAXNOpvVse+zkXTHzJmefqc88F
Jn55W74TOy4RI8iBa5pC9/uVSQ4QKBfDuC2HcvP9hG4rspphy3I9XRBngbNiUPAYStqZrinYyaZ0
pI3JOwEykkU3hZtNVOIL2fp5HX3cA37yGQ55+M1uD0jpLKFFDaGxK+GtFwr6gpjvaWQR6E/Q4eDi
Q8eVmUouVhCJ0WvIIzHSm3m5sDxwcW7dY08F7Cb1pfvrdZm8BPYmDPltzXDRJVWtdlCEScaCgvf9
ehcLscEiN1YIdKksbmtDhtPJb+r9pQE7iQ/9WSFKdLAYRW0LZ8um0uUAOtZBVAtgafSVrE1q6UNA
aOFwDtFlPuF+WJRU1VKvGolrWMNZ7vJfnz/0oXvCELAPGY2VMoZHprC3uHyVvKCILX+MdF3hJ8RB
xy1tjVElmzIA7XnIOdu5iBDiYS11As870n7DPg7MopMwrho7hLfw+sPfoARJWpyPRKfmiJNXS2oG
2WgVOmwfYm1qa4LfxiQZ2ZV40cLzRi0Qs2TuBBaFZWnS9yLunlx7eyLpfnYTWED3Ehbj+qp5X9RO
vgmZq8jRs4vLvqcyURAZt5Luc/jdYDaxMjJJF18pq5uoM/Tgb/N/ozoHakLwEZBf8qn+PfSNiEAW
m1YoDi0gAfh54p2+3qMjctF1ZkFjr6LE+IGks2TFnqjtf7Evjz/uvdldidc4TNBC0z6y7T/tQpBo
NWn42/xRktEeUgKM1Gxy01Lfr9+bEGoNc855/TOaWhhtaf+2rNuxTSFX+7xBOigDHLZjBX2RvRqN
g+XsmgT17HvzWn/cm2GwW0WWNaYixN4PcMiYxC6+Go8zyViZUeLL4XqecfGjSj8QoW2P7UAyeu4O
l0l7C1ByGM9dYW83bd/OYKnFDzQpf/p6A92Xjiz5nyGjTi7/3kr+71LDoS5StnySfFmJrlK9FPdV
jBZk0ruyzLUrVlJmh5z3kWlpmZid/gs2SiwnDOpbfXMcXyo6mHXvo0nxYZllcf+rML8/S7zKo1rf
eLiAbQh6e5JHlbyt5uArmH9AF93bEj4991s2432j0/Mp/3YNNbeH9nk1qBjNcPWqF8Q5MYJndr7O
2c9Wu+JhCsMGdkv3rxQ/JUaXS+cfFiKzaSkPIeu8PethceR/JhgWc6uA0MZh2yoLLxM9qOf4lAw0
6zErR3TWKQymh4/aKn5jCzc2qfNT3/qc42sNic1vWDDaMu2Oe2iNgNbLaOtBP7gePApG2y/G9I0F
bjd5GnEgwqfSFjl4vl2GkeX7R/Ph8fpRpng7r150gPS2kUbskLTdGt2Sc/6gf1N5uKD/GMiAe/SA
uFO4UngMt5OFDz+x8mJkcX39p9MEHtZjebVFmUy4JO11d8h4ISt0wYNzaPp2OhwbIazkpa4VllCv
LZ3d6nMTBJHVz3VfgN4ITera0Al/KSJsUSxjnPG3cp8Ne8abQeupdn4GN4YNblxwGEwulAyZEfuO
D6qYCdz/MjJ7w3xi+BgNEAYKMfd9fjKj8VLBf57FlbG/LuZpwdS3+CTqGcCppTOLKZwoHFcJYMAB
ahgH8u9ZqDDFiU4fiTOe44GinvFeBAgkrWCCZgdQcO9TS9/L6ouTFyzccPKq0pWkQaRdvNzYNRKH
BqSHJuc2MWbaac5dISoQaiy3mGwmaNAgfcm42xlmv0j73vqU8kJp9EnWCz9ihi0xpshFh6CAZTDt
+ogRsVXjC/Bpp41x6TgenS9n6PBPl2Gr3SFKRncSTcZ3QM1nt45UjvvTq2nRDW67MMGsm/IMh6tZ
C+EadIz/guE6E6m9rIyUbsrOZx0gW1rPdE5jDuNUM8/3W3+bs0KJmr6sKgM4XpQFkyc27EYDKjKo
5hZP0m82a1ffLAKDu5LUQEJ6kQYD4Jml0zyReFKwCMx+cO29CssYhYcozgWNgmsNGJqSDJBlf6dz
8p2VhIHtzc3h30Zd+/N+PQTzboBtKtR6y6fdwmmuwMLEM6ktgs/lVwma9f5/3YDTRMcPtR61CnuM
Z3PHU6TGHREpWQy2gbWWXF/s67zyhGww22skK4KIx73ofbJ28bV5IWtKiobfF/G7ri53UEzZo7PD
UZLItq/GmPNH9iQXbRDiOD1SlOviwo28g8mHxFxWloY50sZx9fXq3EsllCwPKI7u4GHOcJyqtFSB
HsK6dXGP5XlbBpvCrI4oGzI5POC5U/GIbe9W4iLlD6SG/BanCLfHP91Bk3oz89/mAS1iLLbd/w8d
XTfyYDwrkmstbqigm7/lj0S2Z/zrEwQKGLJNU8cw30E7xrolv74T9tGBaRskFw8lN4uifoLJP+yM
wigmfICnYCn012BUnxEd+joJovN1RajJs1TWE4uJr+eVxFg/bRoiJA4U+s7kSi/9ORh81mKcFcVo
mty0zD0xnFWPrQ5+tGW6UxnRDfzAjzLN4Y5h/5aecY2bJ1j5IpMiJjTPB9tgAiRDdyAGg0v0na59
Sqc5qlnXELV8IsPqJjvqYYe4dDAJtSJtbv/uNgXo4+I/c8KNYu2YWhEYor7jJXzMKWSFCnbclHv0
NAH64qnX27sqXoFQ9tLEQSAjl6nJURjmDgM9yX3POfeDaNkoZIC+UKisVbVsKGDdcijDJPjQgS7q
sOZna6O87F61g4NPwmTt4vV+Yf3lAZirugjKmK/zLSpfqFivpymD1f/HAQrsXVwP8rPErLoLzEys
kKiinq4Hpa5Y1gBgL1eU9hc2RwezVlT6xxIwZMm8m1XMScgTtxuvAsQFMn3PO65ClWR1+C13wSQi
9o7pqpqjEBxnplOWCWuZySNZ6YHM7aWT2FA8EjrvNncv5psuaU/KMsCHjVoas7LI8NvYEdBnv9Ce
I/eMxRMwb4q0UWjxgo40Uf7vqXj0g1vH7f3lpjFb1Rrsz7CFJIdDIe6vdP5Sh6JqjtultK2VLzH9
4McgXnP3Wpc1/6Eui8U8mp8z9M2fuN/ouebvGN7yWFzxr6TkaKhjNhwSRWROU/JK5S4n7xD/SNsU
lUgJ6Yz300Cs++wNW1W3irDTjO36gvliY6yRs1QGD6HhC+mKEXF83T0Xu/Da2DzvdOu4hC77TDJY
gl9+px7aPNpR1Nx2q1cAWaDLjce4TFNf8nVdbczhpTrxlu8/SqiotKNuutRaw6AEHCDeqdHJ65nn
KxP2yM/ml1dZBv3xqPwsz1XU1/yRMHKVCZDgv/TPH2pZEF1CXAh3FkFAtZJ1wNVmGYPg+OS9a16L
LFJZ3sL5AEe6vUAJCmf5NU3LTSZEH6o4ZCGM7kuux8BIcvvuCLO67iy1xYCB2aNbudpKtJh7jNhc
L1aMxzmCWiQ4x9SYCvwj9xgLJTeFl0Ha7YhDmgEONpiqsQUGX5pZNu9St/8+aihnUTMJYwa+JLIW
gSxCj3Or80acuItL5EFmeWIj6rCNsD6fTtACZsvY7m2W5I4Y7vb0bwfwzoWSj+AQ5rF7rpd0MN4e
/Udk1FWjfvV6Z6vRuOM3Q6U0xQlJoslEPIMDKkoPZw+gtZXLFo3LIxt/7ZjMr43iXGLDJ9H77U7D
WSEiq6aaYZWCbhGFABSGIo3MZC28/e41BdmhPRx8/HCkY9DYgXj5fD3CPQDgaH/+v5G1HLEnIZfL
KQF5/9hergNdNVbtK1HaiSIoKKNf0KbD226EA8qtghu4I3Lh68GnGCebJL6RbSCcfIcB0lmhR6EL
7pByJA8nFfDbBmPbsGmZsLt3V7saG6jLW5qFd/rAA1i5hpRs8HMVteFnGT+KfkWw8Q1tU5ud8aWt
A3cVVKm7te5zTYpUQcC8vHj+r/hfw0YPqMSwAdba57/QtoOGnkoEwqUKj0iBHhzheY6REwWsCGjl
IpGbyo1K5FPz5VBUP8MBCPbP5kv1T9IMsjG3fTK1Tq0OLB/NuvNTfwTB/RLDg5SEDyUMJP6SUZrx
Tfws03KC5wlphbHZTVW9K/G2o9YMNT5Pkrp+cGVyYuulOWvGp1tChvzELYQq7qeQpVEpvehS5/c6
6SZ6h725F+8NGkunRlBFS7/WVOWfoW5GoiAiAaGZKnSgd5u4HZui5OItm0vJmiZIvMIgN+2+3We8
JAZrRsZgY70THrXPmXpkdzv+4geAfF81zbcrne4OJsUZsPagGqF2Mv3haa0dkUFfgZvsscruA2Lw
hi14bfma0uQ4DlZDSrHuvvuvyxnDIgUg7FJv0QjZEc76XXzenil+jC4a5LViIOSusS/bE0yACNvo
bvjJoSLPozd/NFNydj2SvsCp0Y9RC7ulUNpIVlB6tUygtA8k5/Fdw4S1epF6WK2f3lwmXRu8rZUH
GLZmcwPq0tiVPlV1FOFUv9/VxYA594btXX+i+3hp1eTzl06MTeBBRQbbnWJ/at4ORuN387MouR+A
4c9jiOq81VDsKHGq0EItSt8RsHymNYVRIEWGBkFp7/GJCukbVTpSRz+i5p+hv4tlJFEp3Lfbi9+e
eq10hga3MXbVXV/gqZvWUe7CJqdPyLiquOIxwUoWd4bFUQ2dctvvbsoWaUWJLcinG/SfbEBRPVh7
M7M+am+xsxtt7E9QN6xvNrXXhdcKIbEfe+eXpPwZMnywATu67DrSIC9d52WfrWENPctcy0Z1b1xc
dPRhJ8XFFNre/YE6rq+UMKu3iBD5BHaWEtRswBPpoEMAusJugHyNlhlEOhUBXQAQbOO9+J+WHR2s
N2fqVFt0ZFLJAxTVPQDe3A2G4ztlrcG2m/39cXI5bcS1g0d81VPPLz0TOgkLGv4tpQX47RgQGVRh
UD9hmgc+cu9IVuLwHbi/DH/OWd1V6jDtFBVpkiTkAyTYBQpbRYEX+ChB3kZ233LJLgxOWza7+Xvk
y9rlsb7QXACLPtIkZ/So3uBHKyNLduqgpn/1SWp9RBQVhWR6q18X2iPlYWIKCVtnLZLke+cEtTfj
kBM2Df3Ea2yZ5AxPw1NHn3x90+iJLQJpT3LX0V7R644qXHFC+KJqYqmExEbxJqUHyBH4QiRjmtV1
OL8GKF9iMa17oqCsF4MgbaXKlV64tHjdiL3Fyvubg8Dzn3ufSanvar6AH79geHbidk4//2Ar/0qc
EGP4YoSJ7JF//m6vmmAMdZMCRbfWHImTp7JQQutR2QJgDQU3rMsMKsG0w2O4JfNSte5NPr26iJ98
iqiYtjweDNj+ogXQ/9xW8UPamjLmVx7caE8Ua6MV6CgXAjVBDFEdFPZ23WFgqYWgTBkIIyQyOTmT
/I35Hg9wZap7+OrRKNRdnSbfIWucP8I4KYwXealtFUsIWGUwPogVUkOUvlbkKo/M6RnnxiZBRslc
SsB0/KFqdqoa28ZbfsEP5XrhwtFUDiuWH+AUpWoWdwgwLFhQXdMJq1L28R2jbXsXI89AlZ5u4zZr
cVCDnjzoB9xjUpEVH/xWZiiY1waEQ8Jr3qN8983m5q268BHi+W96UhaujvrTJgaYyy94BKBw+wTx
MopxajPSMpkucnVQ10Rz+UWJdaIFwJ/PUkJ5g7I/2DLp2GIfxSQr43HBIetWzPDd+MAgHMfOot3L
v8TOW0do1NRVJJBBwjbtypuQWhRm2opcG1YTkJUs50U+o76CgGMhNKDdIVaTsXLW1TcyqdFkVTF0
5f66y+Zw2PhdYxwGa71rgXSl6S6IEV/S6XrwP+dqhUpv0rq6YzHODKIrkd1PXPbnLTWyGaN8adwa
ha/3yfM56P36p2agwJQY3Lz3y/GC7VVlPDVlhdXaBtuy0KJnltv+3GmrXHy9mTiZR9tmsf4+JHik
Xd6l0ClhTU+K0Ht7zdgrzwMHfHZvE6FPAsbuMDM53ieT/AMzr5xeV+zm3fPdmSn6xBFPlFyoFxuH
Nr0xyiNP4LBDRDg7CkYjlDIJI6KchlKFAcxav2GgLjb23fqdUk0wt/E9hJG80viDP7fmXcoJAohR
fhTggMpTxmwnHh4HANxFXEi4bRH5o84ZDdqaAIjxLGBt7XATlr8rGc8yEGVNkxQHyuqrtZkkPJmC
nXSXNzEbyd6qEzgz0W/B8l/tpXIbh6xbXZ6S7YG3ktapM+yjB2I9Q+4oQu2B4+EEM0sAQWqCQH2J
/raRsXvo5I0MClO4vFMFVSRrt+C0CYBdVVdmmS7rXziYlhQ7txYzdm3JJXO95wct9YlfkOPJO6K+
MiY33C+soWuieQtXd+pPkMofZxGs45G3YT0R4IYA1pteuWdgQ3KsPvrr8catfJZ2Yy9U9/U3Jg9G
HjQ9k1zbUA0RDeWsv3hhvJw1klyrYtBLQasSYZtd686f/qUPJ3BcMPGpD1TkxgVjPhY9sRGyGmyr
Zyi/wty4QhsMvKBwDNJwswZkYveCi6RnPhVEjooanqBFO0I2cfBrbKi0z+BGGoajML1VRz/8maMd
muB7eT0U3J6wifpJybJ4xyjhtZp3gutImm7GvNTB2Psd8P8WZqkhOekPmpnpiuJAPL8wXbLqt/Ku
f7KqhANC0EoEpZo6zZilKR2YHcGvCm+I4d1IJ0/Fx49KtdIo95V8w/CWuDoC1X2o95ev88ozIrJn
fZnpTxjwHxnaHiNSJZ4yvI4+sB7Tvydq+dwUpBF2I2As2fpDEzteMhWZMdnL8GeRzQ/RNm5p0Fuc
teqKs8FeBk7mLseSoi9aMWqQJ4S0p9Tw6fJh5PdipEV/iV2DrfQem6YnLGyOhYuou5vmF8OJjw0U
VF6vwcZHqXeMJ/Z9YH+DsYL5WsGIE1WFYeWfP1wzOhak6s6OQPGdvT99rrUFbAtwD2XN4a4unRD0
zZEFtd986c2D0G/FE1preC7xy5IKRer5K+tnBRk+fKPYavif15HC6X1Vp/ISJAKAy+2Qk1eQkjsx
0Eu8i0+DO1sC8u5zn/5MVQ7pcaDlb0+FTA6WQgZwiZh/2Fyb0WuU6Wi7mK2nULCOOvdBrarP5gBY
pUP3ZIhKHfM9voobCrtAUkPwgzPBKE05NRFpKdb/BVlJJX+oby6OoRx0nH6sdkQxjpndfVQgyuWP
HRZrQp47HVPzUSnlJBroCR4Ti7FDiEK490hJhkma0OmAGMleN2WsHz42e7RSHngYlu2x0RWsKNey
gp1r+FoTpK1a7RjEtJdUAztOLZ6EIcEPFQ1mxFIzUbc+n5WK71BLcoFSBWLfPKEGUyq2mVUSx5oX
3XxKTfAOUf8aRDMSS8n6r4RjGHUz1h5B5x//8t2B+2Yyu0Yg9GyHr/yJzmxp8Cdb4kWUEQj72uRE
XLFYV7QoT+zA8x8B5PjZE4eEQtidYk3RlDum8J9CToZKFTUVms19mX7Hhr7ceaZNxz9H1opVK7Kj
T3qQhhED/sNfubvboYWpVfo/pcTEA3HAdPytTnpbZrgeKF7Lu2OXjhP2QBknoGplv8m45lqLZQrq
bdj2adjOvWFVMCEtw1ifzWDq8yQncqwzW3S/ja4lIExdwvnN0hTyFlF6pBeYJ6s7ddOJ74/JgkG8
nEJ1wjFqjw2LK7ESIp+0xsJpO/jA8ZvNGjCb8za3QqGOWQeYSFHFvQhOmwsaHSHwJTvzZIwZyjMM
HtHqWVcGM+/OunHdhyyhh4QZ6wIqJvOaC54dWsYq5IEu2sFjuQ4ZEv8/+2HOPGPhbmMOewMl85Hk
ZuOPAczw3QSrkiXjltl1CEcRfYEz2GRtjsLx0pOeQ23vYr7vVBgZWbVSvvtBHwXP9ZQzwoTTh/6G
8wuQxU2TjggkXArjK0L47RcpxS4CbCuJg3LCJwRYv0tFy3qeSJAHhILJg0kM0W4DM70dg4NiOQps
yVspck9H1l+3WKLCRAt9AzWga1e11A2BMgXsCZcMqoLc8/4XjOy5gJgj7mo6RtRrYy9/LHL1Xxj4
5WTEOifcd4Tw0xMRd1X8HEYB2AzuxjtiQozRQmx/oiQtZ7NdyHT1VDg1EpDTi2Xtkjoxn/D/mGaV
bYVKGqAS0eKmOYuyXQCRDnG75a1nGCvdP/g2naXkdBdJo1cSAgB+ukTWF/8D0GeesxJYrvx+6Vn4
aZAdFmTN6vLvOna/dYy1TSw9+RLeeOt7GAFfd0lvlS4VkiF55jyEUAlaWtf93eNuKvMCNqP5g2Eg
oRyW1uoL7VoW9mxU+thyPAGN0+OvHFJhTVnAcHYBnSAWtjzz4gTPyZ13xh3HJeWgWKWZqFBip80O
0V4xONiMHTsX/vlgPbpdc/Z1SwEWaQLg5VKi/adQLdUQMZA4swhsowhOHR6kVJz1+XdyQxw8smMD
chNwX266AMniiIk2k+RLuj3kcidZv2JZmwRPLO6/wpdFgWWdqirru0Bo/eL+YmRV8lJZK54Xu08X
rrfYolpkiMM2DJySSHeDmUB5orZUpesbZBP6wCm5AjLcvAXqV+GuPkw4/G7EVqvIvHUeza6Gbg65
yn9zg7tPTjls/2Bb6pbeGpkqkkWqf8iWgHWKEKrWzO6ec8elqn6r3Keq2UV+H6Uf1On7LWZR3o+n
2B1n5+LUAEcGP4/d5bBBT9L/U2k/ozJ/LXNha7t93kVKCxgMszW1wl6g4KPsgRQhL2HBgQXtut2C
1jq5JubNHyjxqfGs9kD2zldsLe7ZKjpzTMfPeXYzLHLpZKBhZluS6epmoWgg8HQA9Vbtgauv3tvj
RYcuthf+F0v/ojL5yx9IO7qGSVreuWDAsJe4QL7Hmo3Tay6+k1+QMmX2UEs1BTzRYQgJaojBbLPc
0fWMf4ALMvo5qNkVkTGOreebi93MGHEjZO8ebNBk0IEtS0LgYspNGCg0HC/mSiR2RLgT13zpVS5h
I3rhXaGLrfhRC64gfLNu9nx19BBA2YfmuKcrnzN5XaSelqTtt5LvDreJ1FmMZmLykTd63Jos/H2E
k54uXM6Eg8cFR092wGYfAmgXYCzZLXpVmM59zXMwxCJ2HvR3kXSdtycpWB576EPjODh5cDj9FgMZ
vvyZI8XsjhaTOtRTjqQfd2khjFs/eopiGYai/ylF6kp9Lh/h7E0dxdXV9zkevTE8B09zZ19Y+l/h
CGFhY5dJ/77nW88WHa4ErtSF9GxDaiCQUA0kC1j+9oruGczfyCfGdUaDYGDvt56DRqIdLeKOM4ae
4IELvrYeFs5WYRIT1fHynow62AjTsmZv57h6lt425HoSmd8mKdOw5f3b/XClPe3ZqK3GpxnCEyR/
abMNeeRiwW1SNvhFz8cjAwNMaDWT5T4ThNeMHgSI9sUbwbGhSCMXT4NsdakXweQp9IgmBifVs8st
Omk9Khw532C3/WAaZGYbhko/P2kEQkvDYUf8O53J7f1p2lSC3PBVC92JIg9BCj68Pl+qOoygPKUP
uhinLVbo4rtb+YyJS7ZjqzS40BIIeJUV2qIzKYSr2+eNYW4jhKq3yERZREAC6Cz820xYYC3uWAqw
tHI5Soit69vbOzaVNrtnjZm/oEaOTulRtG7ckqZkLQ9aLJvV1C6SZ38w7YTbvzsOqSt84fdC1L10
i9dZtTPIkJ0fuBInOmObSGQLnOtb1579xlQQEFjKkhIDOO5VqreC00yzk7z/LDtl1Mf4DKxR//T+
pgh/F0eB3j4EbJJh/6V18R67ASuGWjGvVsVZvD/tckNlM4gJQUJkZ+BQK28L9nmHqefUe29vT13B
mkYbiYLWnPxDLsqUiraysGlXX16s7AumdpvNf9fvYTbiVt4YReYWV9OyltiPEf71QW5r3C6LzHfR
agRqC8EH8p9sOSGfIF44vyfUbo0iSZmYHE//kp3qVOClmgQREk6rNEkqxpmbMQVbzAJ7gwHGxLJj
cW8fate16kkScaZQ4aThDl4kf9vPsPLJscVA1gIcQKKXwEvgoPXcEHppiHGn5rtOC0n6UL7qLTGa
T/r7hNBJbS10CoaY8ShizvUebuDZ6HgNP4GC4WfloKsTgVwu2krl+0eu+qoyXbDf4qy+ZA2PcaEp
JBt+h22r7I84zzm56ZeF8liKDbCzvOLrawFA67xf/fbDE5oNtA/+Paf2nPwSTzv3bEKFLtv6de0t
HIWBQwOvpD9RPKBuKXVuJTFHhEnkd/bg+dqRUS5RXfLyL9Z10qW0eDbPYMlIRwIIPoQIjHTIck8q
DSzrAZ2+AUHDa1KJxCZG8XZPOIo4ZvBaKuVh0Hir+YJY0TMNl/MfFXKw0RNrM8Cp9H+zwiSUYFVk
ir6gVIVNnhydCekQG1hW+U/Cs/htGxPNMhhy3MUKu6S/oj8c5A2WVH5BOlmVVzv6vFWo5I9hzZ9M
cJV8AEf0IxWHVAYf5FyXeXymhEhUTeAcg/w9Kdxicsszax/CxHy3BHFruka6hj9TbP/ca0BCKyvp
A+CyhHmpiEz3V+VyY0xDgIOkmN/uQWUsWPBvFLAkfYZhCuDY/oypA9pW/nTGnvgJ4yCvnoisc7Nb
nzCpV+UUJ99jdy7Wawh2X7zHII3OdFL2UklFUu27r60j16EvpyeYy0I0V4f382QLD4ZlZCdVlzWP
z1kh18jo+8VCMlB6+mQdDffq5TcFbHA4LCh+CYrau9ASfyyjWfb7zk+ELaOG8uIxlZ8I6H6m9ko8
8M+LSfI8rUysBtUd+2A4m5TtTof/VLASOXXNJ6QaWnWV1uSg/P+4l+XLj4rtgGN7jlDxOFvhenIm
HkCu1zGkExnTJdpI+ESqs1qye1wj2l6fXuYY6KaXuMN7rafTATnk9xLhC3+I9U+Q8chXDn6SSLHm
73xC1mD20d3C8xfnIgtAwS8Xa4zwXBpp1tK9uXHCAmYknGBZ7wk2V2hVYoEN1rJoJTl16jej7vSj
bxz89uFfEZPtSKSMjKZmeGXOJu8lar8mRHPUd99Yv0ERA0K2sZW0wOa9TEaHZOsoyEv0s7Y75Xvs
5h2mJJr3HA6wLZMFMjuErnAYr96KJ/dXAlge3fvBakNqkoh0erN0W7FuphQVFARrFtEHxIZ8exyZ
EdC/6/0jsGEVz3mnP933qwXKAcmbTCoWG2RHzAUuArdlzyvFgqrgP9zTfK8bHVgWfV3bOy5npY7L
hF4i+Zthkcq7by6ntkyq6y5CKFJpkI/FXKP9P+qC8W0ODvNjBi6I5lVZT0fml0UWUeunDnRBm0/d
PdLDYgTcY3IIe6seCZnyY/cb8TXYGYwmoVNdCgVXlnC9oInf1f9ixmgIDHrdfeRHeJCjZeQ/xExW
hzle6Fd/k90dCG4xNsruNscCfcVtSG6I1bsENnU7mJgY5Q/O6kIet39G7QE1iIicD/gTfZP37S+T
KDSIFakZGUEJJIBWqJ3bb4pwY5P4y8rPtg/CJbnzq9r0DWvwTkH1l5M7pzOa9Jn35cPzDXvMalaA
TsJV3YMs8Vwpm5lSQSBrv7gOPh8vJovhfyRB9bRxcyCcVtmA3eMIQm6JYJgf+bhiSoNc0PNIw9iN
kvLq98o8b8Pymr81yM5AVPLaqRXqvl5pDPhY0bT+nTKMXb3Rb0FOy/l8XoToSDPUcY6oc7VVOTIw
2/9pJt9yhvqWnv6aynkUl7PQpxs0zxfwS7l1BKhpv5CphkDDN1mu0Ok47IuLbtmj5MlRYDWKrjd2
BQ4wjTrcAnk0GUxxWKax8knRmVgi/QaZqnB2IjTw54BLWX4BZXZ03C+bUp9o1BEWhWfsm3Irzt6m
hD7Qrqs/7CfcADpycPhR7t6ZjiabONRc8TYNhTNDSr11OJ08hP7XJw/MEpFTTDbasm9HaZz7YM5B
io4yPHiib2oT2AmIFQcCDFvwN+y8mZk0wfMT5S/lQ1FVdyg6AIYSA/xHyFiTrXUUNJCCB4dTwiA3
AJ5QXlIcQJufZWvvZGT5k8Yi+siZgPh0JxKFS+qEJd6m4Vhwfv8neXZZoQB1XRz1WXxbece2d55X
zlEgzTe2uE8xOqhtIxJI4HNHiEX568CCJCehVlgx3EOWbH88DhZ8UF03vE1zVA8n2IR16UlLffeh
GhYfJpf3EFgwZXi+iNbc5Kg/3bcu4uSi1guXHw/jG+KmFArfmVHodufz4MBzQ3x/JnBMYODrREE/
gq82Mdyjtl5ahT3ZTmNMvuJ0U8Au7Dx8ePuQnCfzszaHPfyOjoSiqV9rwR556/Wg46tuWK4gIjmV
UJ6e6K2XjTkX21GdhuisFbFRpA8mU3+TMDSe6c195fYVJzeTtIsHa+FfMzLYXsmOw7vqo8Fg/0te
C2dqLvKnJm2/6Ex1n0aKTm7lpQaLQKmeRLv2DbpbnkIdNS2khy0tVV+c63kgw/iOPh0wZL2Z8+KY
EsqlBOlQZtc5OwzidTpTdeqUf5eF22cUPrrHsB62k94sHrv/pDmsVEiWbaAogB2ZCNOGbBrQeV0x
AZY4nsriB+RBnaYFPIGwtEd6lOJNPDdOWoxRR0w3ldn8wOwD+dZi9pQdLJ8FDDmZnvvdgmt8ZD45
t9x+BY6JBjymppOq3hPuZeI7EUJjDm0kzyNeCYFbvbjmJ2F7IG9f3xEJp/d4tNYJe/FCHjnZ1M5/
CQoDASIab+c5M21BTsSe5VJVYoQJgZorXf/wWxJRc5gPLZiZ3WumGnqmCNA+4EYGktrZUze5Q9pX
/FZlBCf6XaAeVGmer+4OWNjq+m+Br/4sTPAYIfX/dJU8/SzVNGpQQfe1pLJrt0M+PyxbCYF3THG2
cd1hcPisZ8Lev9YNlCQcjuEjd+2e2kyT73yy1fPq4gk2/7IjETpBjDpjCcC1yaXYdGJNLFRnv2fx
B1WjEYTJgs3W44bRUyB/E+WgcdlBEXj96c+VHH9q1O59nkxBXNu3bt/Le1a5qEdrCxkOkPrWz4O8
6RCjsI9IVAD3k176sRDWhgL4jgyEtW8y30aUyb24AqmKHsBxhOgWJ5Q8TsEJb1H4TzDquEqIJDxC
CRypNc2DRYSv5OJlYVfJK4YrYmdUQXCEBVF9UlJ3F6w1OrfhWONlA+HH0jVniYxbFVHoDFx3Lumw
PZgTgCUthdvqONQeyH9pC25sIQFIJnP1uCw28Rue1lBtvf+mjHdDCF+4htDQUnt+IBAZarSA7sw3
I51NJ89osTficSiALudfpVwpa/OLN+OYnc/3v3m62AylmFRvbPmTO3uA7DHYIuReomC6wSPBhNtM
wWyVqzboBLqqvz6EmMPXvGhRiZqjaQ3GBsdEqvXo8r1Z7BvDRtHfm4asNp1eNAooyi0AjAD+vTZZ
JmcynbnWYp2MkWzng6CVGXi3PMKlBUzU6VYYbfBHDM+3Oxpc1eIcBHz5pHfo0XvZ/7l4GRGrW0wA
Sy7nTL0RglPsGD3ijDXb5K94c4SLJJAL2gbbsKWIajYsXkqBzL1KF1WWX1Tupv6YtnAlM+dj3MKk
sKibONWF8icYwWgNGwM8eQhPe3TRcPk0EfKvn1/De/o+uKLLsHnwDTp1MpKPgz+d4744zfS0r5vD
Xt5UvXc7F+ncdhBhjkaCvUlxg2jN/rJK0oGoIrY+ypyyEEi5BoGQ5Xz28wgqxNnjY0NkXlHD6YMe
TcAk/kas7dffZLTAh4dnRa5dys9Bhs+5ufOHUADmZels806TEdWoOQqa9kUaP5ITuWmQACM9uQyJ
kJiv25K8jgY4cJ2GQtIdx/4+KyiIzlVPsBOvReFu3mzygIfph6nlbzpxuhijazXQU8f5eC9dcono
hE2GKWkR2LmTBu2ono63Ix6DslzOXcd7Z1lpknYSyRKR/JWyJugxFDETfYlmdfCmrowrKNBVD3Hx
yBQABwXvzgAxkVSNp/GKHl2+7ImMyPrtBHikdSxcCQkdVPjwysYzGkwApJIXmtMY7JQax2q217AI
evdqAecotUmIfYaw2Bl/oEkix0vxUw+FbPJz8b0BTIjL251cqyNo4kgXGJ417hD4cCLv71eXNWXN
jU81si4lx4qf6zURo138IKJO4Ck1xd2heQX17TQHuQ6uPf0x/vatex46B0KtwGA51ccDjz8hRZGv
h9cdN1M5s0JzdrlFRCiYTtRNQHEW2ISW9WlzWXOCNtqWotgVYVnSaJDG7Rx5aKoR5QaBFEbizrj/
itVX6FsLt6EJWDM1dRyGkVMFglJz6KVDP0ymXRaSU/u8Jqw0w4oVEBw7NYoM3DFH/r6/dVFbYSJG
XsXr6eKDFu/o0nag64IT29kSuJAvzgeDwl4hzgkcKxy3PJxW8rzR3kXQGEKsUdWLlRGw2G/5BZYP
CjsmdJzqyZo5AxJtrogH5uSVnJBMXW9dMNGr8TPpx/n3BfCcw0nGfLhcpZAugF5oY1/AOgqi+blA
BATegEFTY1XVy9uO1DKNVvILd3IA1CxM1AD3LuwZS45NTtMR5O7mA607q76jK2tg48gk2xJm+pKo
F/Y9vf5fRXt+fA2h22Hxya6gFtMphZZxPculsdOi9GZPTSqOaoGawqANOuYBJNZuEogZ8p/xPM8s
xu43H9OhNbIuJNkk8QBFI1iA192Vp2p81oVCCLhhw4z6ZyPNDoo0gOWiziU4H8lKZKiaq9tCa8bx
j/bn9c+YHNLAx2rgTQuv4HIK1OcfFP0VkNsSszDk/h+K5x6Qg4tdY1hFqudvMH3L5nUF3HPNZC8J
6NyUfzYHn/4wbEx905elyOlXlNrpvWLv7G20tAbBh5nwc1tVF/ljvYFNxEChemgDfGe6mwnMKGzl
+DJlUrwYKn53mJvMLrdtSD1JJbdZIlRvVrWe3EtsHA6N7McZwrpPQgYjfGqyydvuoX7QTFPyOOcv
Cf7mCFJ6o5QOTggMfU0/xx7Y25rsVxR38kyrXRNeDpTYu4VkR3fT8q1Zw1h+BvJaQGhQVPz5kqTf
zva/UxNuJnnkt5x8sQ7c1hAguct8CBByrxFxfyQ67Ba6YrGodDH1mvKIQBj3eutlFMHhP//gVrfg
NgkamLGJbz1QxsN8DF+5GP81b5MpoNd9sagmNcoyWBRfH42ISkD7Z+rD3bvz2wZgOfN5z3guk6Tp
cKeuYiGrlBSPhWpxiMe7uBLQzoTGjomscO4Ls0JjCiPszfgHUUz9fYNCSSZNZSmXW3gOBRcNHmBP
lB1pPGGTEo9QVxbGovwtSmaJ7s4GsQGDC7lMwl7ATu8zsRNSC65c3h2v0CVI8oZQ8wUi0N6tgBdJ
v+uJ4DZYIPer/PfqkkieelGJ5qOlfneJo1jrW7VGcEHRaHo2WCOp9rYYxPmDtx6KGi0Elfjc08sE
rRoyC9u9IZzwcpi6aeAuksAh6QOJQV2/2Zpormsu3qsL+uC9HYMlRn4hREGEGR645q1flkEuRmLi
rE9Rs6meebfgBywyILJj10H2FleHQmLoSfGMwocLJWe0eygqVnuMAMGhkB6xgfWInMVLFny0WWAQ
1N+/yg/ASe0+bW9hJl5IWfIBZ2Kg2Juma/wpKxvsyIz5i5uAD4uaStC2fIbgKXW6I7yRTz11UJAe
quZmfnmMdzTDJi4Uj5fAYpR63ae1L9yDeULp59uHxjyI67DTSVzKOnnEWRigIpSb+28CNNc63qVL
cLzX3DE2bH+DNqZnY9bHH8Y/johzgn5Hi9t+a476cB95ATEQIlz0IsbhtLc9lxT6ygawS9DggiuG
Y9PVlLaXYBQYjZ0bnWxFgoL/FNoJaTtHGHkCegRF3uvarypfhmmRLPN4pH2bXIacLSownYx44EYd
scXqxnycXrRFPFSrkMUdvS/HJ9KFdcPNd5dZw9HeEkvD1f8rqwSHzLuXPX5fuTv365VTr7yxhZln
SOXq7SPSlFOJopVAMp0Oz9NYMjFEV4JP6cDNtTwpShErsb5dnRX2rhkcdmC3oQ8VcCwRmMhKByan
QWQ1NWbnOVHWW+TAug/gd06bBhPoOFztEfpq/+pEi5JoC7VZ+k3TTW4zHWQ1dJgQDMdB18JNwrZi
N5nsrGh/KtITbHR+AVq8IcoZcSSpL1sz75g0qWfmxOcadD9RPeGVVAiUgNzPd+58H1mSDkseYlux
XabaJgrwsAivtOp23h6HRCVFSZ9Z8UhgHlL/wjUT40GBZeL7KatVRRrSQqrRoYMxvAkXd26eiAYz
wUIXogQe5hcxjJnq0v41UlnGc2flzLhmCpxCS29k6DmeF0i5zYrSxujBHuRFfoQQVvE6xQcNJ3/N
3Glw+uKBDYtAvsVzYXrcLWFpXquLlLWgWKXA/JmbthAuI4c68yg9x3h/845nt9km50bADB/4jvJF
GLICiLV/sIoPhWIsn7IEBY/WbfZPKpvt32sYF62pH8eLdoB/ZVn8NGEgwgVujPdleaog89v7l2W3
IrP6BtfTAj+Xn50adX9BrN/Vc6lxC2iiUriL6G1cvuzpbXC/245kAQjZq1kw8tOxrlnWr/Jj1wpu
3yVEBqmQ2qiXu9jtrDK5Rj2TaaITM3478x+F1tWKNd8yrmoJtB90Ue63/jssiZF7D+PRsBOBb9J4
zuKY6qFuTYgTKlnQ+QyOMIIzveZQVAId86H5xa8goz0VXe+KZXpNQvrDJ5/0WmQagv8z1yTnKXt/
5bhj3QFrJ349NURdE/8qfh2Q9XiOeJKu7iCygNRAEokGHr5UGu9S+PIIEFjbHMLh10cqwDnv8xKQ
XaCg5Qy98HTLIgvviW740r7A7FyaLFYKfMArpo/+39v8X6aUkXFLNybhE70KYmc8MOrm7TCAkh0b
2EEz14sJPQ8eIEDGPSn4di9LxNjF51STSKjXgZdadT6/DJ5aGF86iIphFNjJ3lZaK0+TzSA8kDFl
FMrPpEudbYLZLw6epeJ2DLoHwOp+gVYDwVK8ErC3LNlkhcdP8j+0biAvoaiq/Oej/PV0umfTDykU
bVRZ9MIO2/o1DHoXBzpaKd0qCMiC1bERkspq0OEkGQbhEl5u1qbnTyJJzf5Yc9ECIJCbgTtZW8h7
4Br+cSJ08HFgg3+IWYn3cH65dTZX+WZ8eSk/GHjhdMEiLveXSPxVCZObsoNXQIlrod6r8TrweDPJ
v2YZcQY0ZSlPTECMa9z5KxCPtl4biINp2xYjIe5FsSYu5QoLb7/MVcRzihEj/oN/nonuu0Ha4ZWb
DsliCBOsiRunI5uHuaRxwtF2d0eyXg7LdEZ3L48Wkq9AcPugoMAdeDgdF1cUqhe3p2WPgdgUq3vP
YVgIwskH5FdpVRGT0yo9uCaNOHr7jKHviGWkxbp/zQSbUu6HeYq9kEIt8TldqA6O1QzOvzZs0Jh2
8GhYYmt79EVpYiRMuby4NV4LAgFBwwIQqbY9u1YjxWiJiSgV1vtC0s2OBWE+3KzZbTDpdfsnTcNR
1BeJuxe1lSMn+fI4uVx+eaZmsex2QtnL5a2/BKyR20NKPQYDpVHVV4ky7Pax1OpM+5031RljAVZC
oG+9Jd1+s/Ed+2vm8BrRJSc+6j2bwn0Fc9T2WgQKCmFfDtpPVy8MviLgs0S8/mKh+hOq8Cflvplx
xRjl2XjDTY0/c8dxlj104Te/7vu59L+6G/D710letmtotuVLeCje4wY8cGxJix8AB4jJ+TX2jjSq
mLUv9uBgxhrpemF6rOy1kxZP/7sZoCS9rKeo8eUr0Rj6LtBZQqrOXiiUn06HZDRdkUjCD4YD77Xd
FeWs4zeTS5HIrqFevGvKYCZGRIE/WgVegQKVfGI2lhnteJjq7PBg0P0UZrlmEBmHqR4db1Cnd322
gYRykwWlZTB/cVEruMQb7iweFgCVgYumM+8grU/XSUzCJ82dj5B8zmi6zCPtZymGu6cmV+VywVWS
0cwieEyGAPPLHbFTrfyl+WUHsZc1bbwotKwiU8lGZeeWr3t0S8a4rpuxWPRMuTJ5o4w2dVSPEtg0
AipTeXy6D3bzM+kY19D0Y7LbjLdCfUvLllywdPMBgD7veIjQEz2bZGOTEnn+0IvUDOkAkvgLbQyi
+i2kAN3zVcgxJ5DcCi+VXALd+OBu7RFOipEoqMEua7fEprFEHQ7tEgNWAt3EJrOzPYMiHzlOSd0S
oF7B4QbjDxqDsopxql58vtuueNcMdhTd3NoNqiXHqH/Jrfa+t2iUif7y275BWnKcqJGUuogQ7W4X
BLFlP/7gL+34uZt0bkHIp2wtg/QnGiblWmtXvxQD1qq2OAdD+LvIlDQ8OAMkUajWPDFe4Yjl/pz8
tA8mh9aIT6v6PMl4dueqqRg3ylYL0J8oUE0/iVBD57UZcDq0ANF5vqCv451SzRfJg2ZIoCP91emI
6xEByaIixRgQMUM197GWV4ZHZY13pCDY1lIQsjN1H1Wduo10qSHaqrFX1RqsxF2k6JXY0D56SqDo
+Z/8zgFmuxGfvZhqUeU2j+lH57zKMnNCVhBlnyBzqTCUBUP+JDb36zZN2RuJCZequNf/C7NbWD2u
n0t7JNnIJebP0ve7RjHYLn/bwBpEUAl0yAW7u5gGdoA4OgwrpTWBMsYRv0CPfm3JWmksnwvIQHwJ
KMK6/QA7N91rWJcEp0rbWAodMfCQvZTXtWUtvetUu7LXENAxzLFfjSt65YZ72r54fRLjrLRBbvHr
3nICG3G3N+k7nafK8qHpTxM7I8/S9fpp+uBZETX3uzAM7ZKy5U1R+4ndLYFl0kcN4N5tFb7J97y+
blv5maKxp/Hu1bYxYzkHM6fxlG56BVPX+cjwwfrfUjD8MzEyQGkb8sq9sGl63kD6aOKbiz4J7+Km
TMOyyBaoBRcC71l4kYj6+p49ap/A2Owzp0NkTf/Fjfsczo7uOkVkfBNIXAnTvwjoZZxKaIYTX2zS
+5NzSdqFc0XF68ubMAifVW0apbFPyUDgOnA2+CsIZRTghODgjdSV0JCZuM8nV2zS/1+xUxgVROBw
EeHKD12MmRIGc0bdGU4Dyb6jW8CAI9aKD5KLLAfN1KR3sZLF+VoURNyAWMYJzBJnj/fy+xUXySVc
iw86pmcfhxWANRjmx8bnM/Zx+emsYLjwfr8AWMpbG39XDSSPlZbt3A7hAJB4FxcndRnAYcrcy3/+
/jNZNBEwdsULbZJEIMyiNNbvDMbchOu41B1lIz4JPDEgYMQgUAyn42Pxk/HMGG9MjYKq+pu2Yx0g
MEgAfomrheEet/xFcSxaOuuVFO1lKY4NvVN1+rtmI1czvau6ssXZ1rE4/CJs0En0LhSxt1d978Dd
atOfP06P/eCAwXJhQpqfXs0S2QqJr03Ws/mm0of8WfKdBGytGM2gFGbVxENhEGVmDJe5+mNJoTxw
u9gntsHyZHbe4hyBwTIXfzb9pzTY87tcj3/PR97Ps+kTAnI4TfQgsDxrcYqdFbMwdXRjZ042MOJq
TJRLVH+DUixybCoTGWj5skRttBO7Qp0EbQ6Xk/ofew/eZqiQ7l4jEfHClQqqG0FTPq7TYIo5w+MC
UY4BwNwgQ669SuxdMk8ukiC93LJFH/IumeFiX42OchManExbcQTMukI83xgYirs8pWCqHPAIcIPR
7SgVR9Pjys6gWdFcbbZbUuJqzo6GbmSpbw+YpwU7ZPqEFFcIb7vGE/62Buyqbm7L/d8aY8vCb8As
oxtlhOxqu9zE5TEX5uRRw/SI06Xn7UkbBUM/tGq8JSfXgQyVNELomXqZ8j/mIzrV7PVsWDnN0w4y
DXBWRDFFjkp71Yb/G4aRBhhDqQ/+QV4mGPGqRcP4muTOm61duFV5l8J3PKAgF4VxJU+I9jPJXYM9
1DSZJo1hojd2k/5bsMr4NXi25wLp1KZsqVTci0LnVuHQlkHoE/2X8vWfpKBbYIdvpTer+EThpY0U
EDD/QdTRJ8s8kh3pSUlFe50GcVB1LXsOiaPjf1BXRsDGIoOqLYjT0HfAnJqe1+yEfaWyLiOwONt7
5wuArLZJF/Giu+SaQybQzaNhJQ88Lu8DTktbfbK6Va/KKPY8RY6aoHHmFLtT+GPcIsJm8m0xMXGk
JiIXzp0y52XaW7eGDAtZjd1wiZnqdn8Rb3I+2DmAEx1+fVWdU0oLkEYgtkgmK/DYoF1+ZL3/nB0D
SYDc7XWxU31hfgmCK99wxnGUPnzMoVp5rtTZm1YDFsRVkDaJ5giTmBxX7dmBQYn47gk193JvPmAG
2xyfH9N6jXoaClYWOsbaWnsxtFhpZgbPP5oei5hZwFdnJiR/25oE+kMiGVeI9sKYQmR1WmKnRJ29
LSK1Wvh+lHYpmvMT+pbhbnzALW187Ihtg5sbJ96Sal612suPsR1ZBQq6wSoMd4eCcdP335K3Yicb
rbFEPUXvmkhfKnuxlnU5bp4quAZpqZuCirk6M0+JBQ+SxoJzag1iYyzyH03c6BGJWujgmRNq2LnB
gyeOazOn4vtDLqtt+8Hm20yw0eNKn4TRgOfdwbqeoqZZ405WNeJgad3Jb1IJfkmFu/8xQmsNAXQs
1ZSO0pfdWNfEF88JsXNm15xpzkENUbGgNtPaYjsHDytZUIv4Ex/4KJ1amkv/XUNfCiy82MNQ0Dzi
pTZsIpan8pUaU/4L5LltRoXgi+BEEirL3P25/AYVbdsOAGhtHNBd+okdBCQmO0X9OwfkGHSI5JAV
F2SgoSMPAe2JQSbpiDypFaZUWuvu3KS8QwQPbTGWlCre5IB9d9UfuQILHi46P//5VyaI+lgcq2PB
N7L6YgGhlmNf6CrojetXZCSvbKOZk4X8N5W1hnUoluT0nlvVUbWnnXDiP/opYjDTk57tkIbaCwv5
aK41l3WTSolM7ES1XT8W3bjsQnqCy759MjojqgO6cxOmun10Yfc+CxXCmj4O1TyeUlQOPec2W0T3
noUYlPgYb5bh37R50hLPgPLyZE0xlrV7h2dpyRPXojf1gp03T3u+KdDp46hjSy4MPQCQHpjqwxMA
YmehA0n8dVE9yvxqmKEYyRYzYKav8OaymrrleRJN4RodR6HNqXNEsXPxOnyB4ZsqDGCw4SArnYmJ
Mj5oHeDz+6e2Wr24hzrzzkfYgAQYGq0X3q+73ixyNlQu6GopQe8v4a9n5U9mSmO7jhGlG7W5JLXO
JdK0zlxlvHk1vRgqVlMLpM3zfhrsv2dTvTm0aKH9AtvGxwoFPyvCf3EHMQSH6pqosJ4vjy08wR08
RcXTl/Lovnot+xN5cy93+vs2kpT4uSiVihzmMw7O7VjyaGuqtTqxCYgz1fOKAuKLoBEzWj1ubjyd
VrEL/4O2w0teTMx3KtgVO9kZbsgUsGkpSUDkfGLOQrovihU7KUA+yJjwhUokg0I5SWisLYpy/7L3
QWi1Rk31sNdeM9gcnwzmT/Eps0UcPyrIyZETGjE9+xnxhKp9QdsO9HurKLJhapcl/sqvlHAjdV/m
/pXeuSME9noO0a/wzq9WG+Rlv5AwZ4xyoF+m0WvDQSgdLnJgCCL9hf9Y30hV85EUkKkYw3/wcUIT
cE5T1VgdiOdNpt7fc/1F/hz6SscX106ngLjo0qxlPtEtvsdPHgdsswXcF5BYzgCXj4n8CnH3Ct9V
jEDhckKR9w70/VDe9m86pflvBGXmUQ8F9z2bwW/A67IMbiiVL4LS36eAuxZodEyv0IVU1rnuLAmt
1RAhsZMX52ajrJNygfBhwm2gnWNnqh32nKga1vD1SyPBueabGqqAoOWrFRTuqISrxHnnKZChiZh9
Q0mXV1t8dbTnvMgc5gwjGvQLbVus4h9eVkOm64IxWW3nOIQxqfLsKDcASJvKNg2vq81EfjQPJufB
XcehJXCBjG1WzBjWTfyVIQymzswUGJRhl5xZ1sE5pe/QYjDzJIcaxpDkjSPoyVrvq1oSSsvh4Lgh
oroV3MIZ4XpCW8odwix1ra1X7X36GR049pzeJuGMAUwb17FKinuY9n1EQphqL35rddfRUMvfnQDO
mUbB6nc3L3JRnlCtYlM3F3mRqEiDeeXUb7wt4NjDE5i/gIecTSy2XGlifNGWERxeSVLhNag0hYAp
XEOV7qxVcm9QRNoWa6IQlFYxvxrDfxFIn5FWErZqdvTh8gEN+1g4ZZ1cTrgAfZNCAV5XupC4zmWI
RgovGvtZxesVn0M7OkFZnFsUogLmUp9IcS3E8cjpZtkqCXP6kEYGitWgns8bBGQN2Vh4eq4OGMLW
Nbf1Suw9uD98NvviOuiMl7nLeEB+VGQdR61uw1LH3jIXildvrSFxpf/gmNC3c8ue9YQSwqChjSCO
V5AHYswo6JLC4vqcFhU65asYtzDC73CZ8b2Kp5vLG/FNLkBO77XhgzdFWG/qYrnjSaLSxcbRwoaa
MjOkn6Zbnd5a+vLtDeln2b2CxPUrpaFp5Wm25G7jp8lfOvRturC49otjYO81JMrVyjxLgGYQvv9p
W94XMMbTekLai4+GDCykQkq3/ULFXJ9ZwT+sXOTQSIZGFjYRNoGg6YiKPjl+H6vT1BpdayqJG/xs
f4T0plTq/r2M1NSzr8WjqkZLPTlhCQPJM7VpmBxgtFVlMLSuEoTUFdJt/N73KYL8ofuY1jNCu6g7
qF3jwnzjXh5YI5dlYcVPovSMiNCKEZ0KUXswa64PDtnJZTVkryc1VWEA5qr3kzI8TbpdGR+Q5zKa
sQkZ0eFr/Yy8/+ykGG2jLpiUp3+8RKU13TzpNgYXvsNYFQ1P3YroSdD4lANWzubkWiJvY2UAdpWr
JtKxCMh3qx4nhcxGYAVMkqI/GXtqqzqGd3tesH9ybzIjLmvBSAb4PlMC9fYOpsTA57SczMh+KA7F
BPlGKoIne8wgavFCKRlJqvkxWIme1Vt4jMaMAYmUIO/NLroC0N8F8CmQrUFXjdNorprp1FWKXIfZ
2nDNAQQkvtQXxbbd+sBAgtiplEKZouDhg95K8UcaNRK6lFFq/+CGFx4/2t7F2rinOeEyAJv7rrv2
xaD3BTwkcmlVNsdOqIVIiMiocI0zpZHmKu7CPnvf2jl5d23DSvbMgG1ffGnaTTKoS+lbBT9G+6W8
8WuN9lb9ETRpQw3pXcBhBTMJSzdT81jhpG02zMH+aNgU4lXaTp287fZwfcH10+is5gZOravanXSy
0zqmRBw1Njtw0Jc9TAj3bOPgW+bWhLa6tY5nHyIBcfb3hLcLYnOyoZz0lFSM4haxOJE3lS3y2iHP
6fGeFBOUEqTeSHFAgliCuZweFEnWgDizVOrezgrIMFm+N9MeWJDF6NrxMzewpciJWUHqL9ECIKTM
2DvvZ4pQYz5LjBLRDX3n+Xv7HbJQzFCCVWegM2f5P8yolPbaRfqV++tnYYWf+ccZEK3mkXQgv4rF
URj4Cs47lWUb27JaXbDTy0BScN9lRbvOUsjRohXR//k1thspSzY6edCt0dOv4hEX6gCx7xdottAF
O/t0NNzGwK2VnYEV5V2UgE5ZkQq8o4bOFOqJZfeyCejJNHErPBeyn6pOVR/Rq6r39EHkb9UpyPl4
VOp6EiNHy5cURqAzHDa06VgePVOCnxmvbq4cpRnIvURhgsK2mqrLXidPlmgP4TgqIMgfjs9quJ4r
iCF69bxrlUT7TMj2enDzNY1yUKcBowZjVO3zJ44GJv6P78YzJmcQyfPr4Xfbt+WcA0EC17fhJf0P
URFoOZzNH2YK7bqEjdGoioKjSO15D8Eg62pCHBa6tk3N2B+bDw2SEwEH4FXWrSSLf92bUmrQGpbU
Rt4PEPH0ZaJhsmHfUuoR3S/A0swjloZE5m2mB4WV+NVuSYoRtNaItTcRHlcYnXbE+xu+CKrKpT3N
c3CyIcAwWRfsCDbBrN91tUG6CdqmVGiKu8U8Hzl5yVJDi8KGp2U4s3gWx5i0qOW4kj0MDCO9IF1J
ee4LA81a54Z6dcqTvowk0QXijW61vY22m39cAO7PDjIqhH7LdK6jyPBSXXxQIHYGlvQte3n4iv9N
0cvh7f0vs/JHIU9Qfgu81H55AiHG4R/JVskHoBFtFCgOnlavAsLQLJx4ZDbIFE6vxomepOVvTNlS
2a6JgLFv+aLGavWMkYPhTdmLrZVlPmpgjqMltVP2uwJhfNLkmQq7c5YXD3KCXzIwkFQOWVLjZXH5
rtamDQR0wL8zeb7TsUeMdB7bWjXtRwdNLs1LGJqiaSXE68tqdGi0MFXEQYjXr6te/OyDtgk/21vd
ttDf6/PP89sVVDSj/rqu20728iF1Jl5TgqUqZ04/MQ4wVTUztcoY32PxzspUnK//O9Pa25X3U4f3
bPxjJt6fFup9kPGo7LbDt4NAabigH7B6yYg5V8hce7X61CTsSOW8ilV+BGc+U69Ciy2c4+EIEBBW
XGktj6Z4gmCr63MVBsTscncg/dNHhXENvEHWfc5E051og2ygb1IBMohNhHdvD9uPd0mzaZvGg3tP
H7CP+lM1L6bKZJn62rZA1tP+ebJNoRTa3eLY8UHHQqxQAbSh1a9XWPehudbsonJY8sn9s3sXjnCA
ZU/qZDfhtHaGIou7SzJpHBIC3Io7cBLjaFXGyw0RKYclr0TY6zmoAG6xlviMzkM9LKbC80qyFqT3
WgAtSuHgFjuKTN8IDvS5IegN6JVQnsxU86qY6W4U/c1kFEOr+O7eJLH42wlFSaW/LB9K++azCyCC
lQX5sEefaERM/IZIVqo4aBek2wjxU/49ZwzkwUbD0O82EqceQllj2IKEkBE+m9m8JUalW1fDzZCo
5PL+/jyDDgu0qH1l7QfYTIE5crVl+YSXBTQ4HzHumWtRme62x8i0SQsyAcgrnv62b7rKeVon0LNn
znr93VuM5DfQdDheze9zw25n/oJ+2zHhIby/i8MG7088/0p7HClN4WNpjMefclj1UOtGIS+7p8ab
Nfe3qDYZE0dsUc33BFSvQMaMBNz3yK3Hhjnl/RYLZjobDKJcXo5S5W02l433sXEdLib2BmfD8mmX
pjkQxNiYc/vH5IBLm9DrgYAkP+BtHLATOLB2P/kWy4fE1BleJ9XNlcyYe9aY0octlEDmdIkrfUeo
rMmqmKUPm/NLTb3uTYlLRlMgXgYmHa4ZiH0TRGWkOyn0yamoI6fTi59Ym4Pjd1GuDELVBBS6fNnc
bWiNmpSt/5mFsVo8I0fwJijzRSL2QYe1uD5DO3cu9oV3WWupmzkteqsTasH2wmBTvqXjL5FIVvfP
qju3k0N3xwNUvzXn/UZqI9jxAKEYWSUph4b9L7/DIJowZdQXFvzYQhexv1hDmpLQKv41nLAE8yZ+
4dG2X+/YwOLHqQ13JsP301MpgqMHv9kp0aLYMsLyd2xPVy71HUONrRM+huKv8XDiOfOXS+UmSL/6
6apaRXGdVyqv1f4rUlalgVUJ1tZcDVunV1bs/XokFn7mKbNRhSZ7jo/h4eQXR69y+tp6S6/tiYA2
fmV+HR5TVaPnwp99jUrnWEwhvU35huM8b4VkF0Ut6OA9MlDdOaU3VaIeh+Xd8RvNFn1wY7a/WZMq
TjZ+1DMZIZ/Yr6MJaoaAb4o7BXtWQXp/LQmb5bW8RzrrZcG5DYcMBzfaLOMOk57Kol6KRG34WOSr
Z1JuCNndHWlWp262o9Hubuvs+J/ECil11cPIThsFbgwXPXi/ACcfxL5cOrWMZDiM6suvmPaOBEDV
g8n9lNOENToMSMyWBVZkZR2AwG27alAjZUVzQftOTgyXdI+7ZTa8XQcvw95TLjqO05DSsfYYCBeB
IzLh2LdZQtciuiZXy3cOm02e0puUeiQgmYbN3+aoz/Nbn4Pujt0stA/Vj10Rn7hFosTZaeSsFRAV
9Agmi8RgF1JkfE10lmljRGBjHe7aYA5T46BBbuyVqyYJdmw/QNwV6CvyMyZJGnyUZ1ws2HtZktdV
WtSd3/87KbFV/6Unuq7beA9tIC0uceJ47TRRWq/FiTxtCuYDHUS45Bpj5nWeJHQ7duLtqnZAYUIe
hNEdqsuuOh7oEAC/lWsdpFFxnrawXsiH/wDCnfrVY5OOmWC+rCIzWW/u/NRGZsPoZTacVjl/eg5Z
OweHbwvZv4x9zc4OvC4F7z4TDDZxkaz3TAutI2+pmWGeeeZwm8dxRE0eXkAH0lu9bLsIF/2/8sMt
Q7C5zY3Edp3107KCo4E2fcArhZrgSdIlsM3KRowV6u0B2EPPlGhSCB73obe8UXbQCnvWs1ZfsoGY
WfnxwAjXVTbzxkgSl0C8QSOFuuDfc7a/IMFsmSRuVzNQ5c5imSN6Cs2Zks7ns/fATf97MkYdqzt/
xDE3vz7XUb7A98yesW4yeyCQ9wyqoHR1nPgHbuPK8AkJCutOv1DZZ6dszGzIExWgxVFk/hB9EVmP
Gc0RX6Q8LIoW7ckcJuelCeSdkQCol2vTlCiUJikOvmBlxRzPzNXV+7/U35gbPm4Wh/LrVLZOADKr
dxUeFF6hQbCAQipXQTXEZ2hkUlwyDajmvEQXgbPhiKexWAAbCkJl7W08BPNfvBq0QtklFJLKtGjj
Ndb+2VQZcDBM96Tzue/fuspkh6HCpr+XBABDxp8rdHYwJsE4ChKzhM0yFI7XEnLmKBTaoHvGHhvy
SDdvET0rT1wJ6Kb6y4fq8xV54oIRH0v1QbXPtKrEAcqmvh8Q1BHyaADJFkr+x+Pmbv0WzNZe1+wT
VXbmzk8NPjKxp6GR6/nO7pnZ630edEcyNBSRtNIBE6tSKEiMfkQ085dXa36pcPsGvpson6OBTktJ
JTO/oBsg0nAIUe6TSvFcMSchaR8SmJVoo5GEIMqm4G0UlJNsijvsMVesltCpWM98cmwWRUg+NGmE
Qp8k/9oHG3gutWx6lKiv0rm8HValJT5Aa0UHiuMcQfiKw9TSWOUe/NQDVgXFSfFZ5PZyKphjijAr
rWPL6ilwB+CWfEbHGYq7mlbauA0NJm1l259hY6UpjxCG395+Xdx3yxCIMAOYsAsz2lmDHd+ibMxI
LIexvij4NsDlCKan0e4/fQECYldA5OaSCpm1/v0HQ3061G4ULsJUd7734M9VmET5h7ufyUXwgITq
rdADPmpXaRemZwF89vKRyRH+8ZQlYw9SBRMiIgYGwLoKbngNzkx98krV7lMBUhaeW6zwCb7pAOtj
pJSm0lBKPdTnlpSiS+ZDancgwUTPdgbNAR5xaace9xbWOS33hOaDT2HCSqSts89xwiWFtf31LCqR
GW/VzC9/cadlz5JSjFDaM1Cq6C/80NrvKCZokhUkUUHBaBepcmM4SNr//gG8li5QzKWpHoA23v82
qfK+CirdVukleR0aCjSJY/6XTaN+bcQw+Ojt0/gM81ajv5enfMqF55GrWn3bbb6kkjDR3Ts9c613
oxH59SRrE7mvzR1aKOxaCeQHOsP36qXP2k7ggCrzfFEz1+kjWJIjIW1un6ehJuU9p+3gABLOeSBm
s9a2byrb/YQ9bktoaNZrxRQsEhAeJKXzghy2gU/dSd/keMiKroA7wflW8ewmHQac7Ci4H9USjWH4
XEuX5LHFEuukXy/PAUnhineFo7Rr6s/p2iTI/Yy0gwygtv9EPdQDW5OLkE8hSaX+eYzyK9+4YaXY
wBcR/QUYoIU+Vs++Af/pMRlCjnjrfR4dr3R0XKfeZSSP+rCUOkDU9SyF/BmSLtI/z3GzsJ1tFVwq
tfyH+n/IzQDTTQC5owNwvuou0BPCMwbwDG+DxJtx4BleXthqw2BQMpHV1WjAmW2Im/BNrkovEQTf
V8/+TWncbEgvHiF1ax6Lg8Fz6aajaA/NBEjFidTIfkh73POXpDLNgtuZLJC7G6eXNgzPNPJitosQ
C9tDMPdgr+Yb8ldEpEHCrGt0TZY0nmff/LlWg6qGI0p1Oolef4q1Z9qmFEperTQL3oUnb2BsQPnz
X7smEJnt3RxZ2VTEfstTtT6pmdiO2ZbJ5TDAE//ztvc8+YqCj5HFXjfYzLSYEYF4bJFM9ZlRTqTX
amDx4BnbuD6l5EtP99SGDHRRp/RpK/5woq6d5lBoLBYc8jw3hXlq9zHTUKrtVe3UaN5E1HmdsxYc
DLqA57LGe6h7+E80vUo99Vix7ggPo9HQtGmEMerlWnKmPlBwzFwhls/h4NWYOyknpkw8YUThWQwd
PRqdzxBuinUKwGwY8Fv1846uiRwPltDzF6MceG2vG138Ltg7leV8jvmtXltGTmvspIKgNN4iUFy5
PBArfBzNOxT9Fch6AeyL+w18VRA690ptio5sD8ZaGONJAhTa07XAdXMkRqIsEOeIDqPL8VQLHlNp
aaxwHRYCS3+dSIjxSOPG9hGtoxEXIN81HBX0Sy9YI3neBE8ZapL14DejfvTMSM22cDdPEnd1/KCA
dphKxGYWzzCAhE2j9p9XEWp1Sj3EN8kq0KqlLa7/SWDFBOvP0o/LMT1lxWuSFej0YY1bcWh0DNsm
6FI4iKsP9NNfp9jWOLUbBgQTin/QyUOpGkm26+6+EW/kmNHQusG3Wmwh/7VOn5IONe7MNbM3jsY3
EDnleyAwIXU7otV6WTpq2G3PzSRDTCpMmN2mzQ0WWMKITFpkvg4BDg+HOEc3GsCsLj3+hr6pU9We
pZRnvkaG7u7zIWPaUopq/7LixFcP16bw4BeSPhAsSKShHNUAqVnqsb5aB/ubNVHgbj/pscGDS1I+
VF5qzZddZKvvansLoccS4l4RXWRBG+5UC1rAljremAPMT9Eykyq9EayWAQ7M5a4zuhQG65Va7Yi0
RSS7WQDaU5Svp3spOQRs7wEMF4/1+o3fU3c+uXMpOZFN7QNvqFscw5enL/cX+PKXm+ovTGSGJKhl
1ELnN5E7BIwtDWZ1ZdGxwMN14ovuz4UeWxc7ku4qbDoYOOeUmR1rAXCwI4iMYcAN+bbbxK6CrZPf
B4DsDV7eNFZNNiqSx3aDe7DccZG4GbrewEs9+LBoig/TGc2JdFGn3tWYC0IQ6q6agpchhCECMvio
s2seZcke7WWg1x5h0SybwakDqrp+PkH1BqftduOq/U9rS+TvAVH7XmPIDjE2TTZo2OZtFQozPTpE
JN/eF0YnIhzJSuL1/6HJvOmqSPXqv1B8KMmiEocLfnKVPN7wkCY7L/SNfnQb+6EWDeBHc4UbO6X9
XYq7DBq3VoW9O5cwYIUrmoJZDTOAo+A8hVGsM0Ng4mX5NvenT5yKPj11KCQ0P2Q5yZPfV0PU4fjJ
/7tSxa+dUtnNhSeKr/V8Y2PPpGealEIJfAdAsdpyBtxkvBN0QBftOcIqBoVLWgXWG5MvryxvInlR
kDSrh2IiK1B5m/pDG4EnZlNPFqcoWJBpInQzTEXXZtL1t5k4sdTiQu0CYOIozBdc5kabTkpypfka
X80hVPnjhNWovXfSMlZSoDCvpqbqe/CYro+lZjQW8w4+1A2QmgiULuuwo95D0vh1R90gMiyEO4VR
D8V1Yk4SPi2ZiqLd2dKcKZbWdPFlqs7RqyAECAe2d0Sj2pBq7tLIlTapXYDUa5D0Z/UHMiyPVLZ+
dMa9y3nJbODS9Rd9GEFQRamAVJruWfPuphvKGn5wbRZ0rnSVsqC8WZLKOuKHNGrhl6MLTK/TsLnJ
HBIJQ/R/A8GZS0mfUslMaw5mdAJfqmqoC+83v8l/CJE0oJoUWyy0wQ7clZSVNNKg5tAHpg7nYTpm
Q28J8RwUvVJj0+McQGzIw4hRi+sp4ne1Yqkob/vinAWHWVMGiFzqpcYqskF0H/HQIF9d0H/8Tc6t
Lufm0xHIcK+bIyCUjcd0nYW88FSvmf0QIB0FyIvtbjaYG1IMi5r3LnKb90ycAPrkBZ61pkWYUHeo
0+cLuziCSfxGcCgEvI/TIeO+SFqOfky+nVGa47FEsYmEZrRVaOtBPJ27CtD0XH1sdZ7/xbl2/Tfg
iVzfXhbsrtzHMivlVY3WGuh96ql4FjwCvu7LROMM0wQwXxc7aqo6DW3qxqAIHuLy1DAA/lg4jIiO
rXTHZbyyBgN0IUHA3xXvlre3OP5to+d3Y5lXEfc2XseLIbIh0H0S5icZxQ8eOK3NuWDus/bW1cM6
vFrViu/8zWA48CMVPwbSObdeERZPMot0AFOSNFYjFujXTZ3r9RZ79o8mKXHs900rIjBrk3jZPptV
lMq/a7VCIgQa8HxcLxEK8yIjoJC59kPPNApn8/RSwlr1iKxiN4qUrNzsu143Ov37IQJv2JPE6lLc
EfbtZfbPlRrV0HidcRsNUf8BUgRmQk4ekHQFz6aMZ/k4IvdgQQ3W0IlQMeSraAHekuxGqvCZYk3L
JREUpnEv33873uYAXA+Lvk+0Fa0Y9ysy5km9GAmHgqAOTsMw2HSD3XF04ACxrImfKrRFivN/j1MA
0BiZl5tGpnMX7dGI+jwYUEZKKwdIenVhuv+ua9804atDeiREE/YWvn0ExrRIepCHZ7LfFW3r2Czu
MBBY+1p3FIqVb36/aIPbX+U2E1sXdirlsZAiFqszTB22eLaD587L9S5pI8dJC9GfPZShXjyTHqC7
yFbU27eeDPp7ZrKlVHkE4ZklXbl9T2Bkn7CpQxkMgDkSPgnHj3+fY/asW1r+JX2ZD7RZMBwnXhIn
RPQUkd+eN57AOJLUWWqS4sCqKIjWU6CxzzyC5VUY4pH8KFx1/+TjXFbgwBn+FA6EV6ptsQAkJSTM
YXGCq4orb4AHbvEea0viJ/Vr7IS0RI71pvgcWPy1ptkESdkMYvJW3dpQLN9M1kO6elqnmgzUafvw
Bqf7AAVRCCd+zhJPOk5iMA/8lJDuue8HZFnghD0j5oTrj9BvfW84l8WFeD7RwJdv9Ub6Ap5usR8C
Yhdnuo514z1tsve0/kIjBDbZi0a015tawHtNnFH3cU/wiZSj7i0fW+nf6UYCzQ9Z99x+Rts8Uoi6
9rjnPs4Vt6DV9piml4+cKDmBCHjYFYhQnrFcBUHaj5N+hMn3m9IHWxz0CpjqjqpgukAd89m4f1j8
mqEiJ5QoA68t4ZYAIifpEXzHia5xJoNAulwyNhvpaOWHbi+7pf+07YuFmFyZP/vEIrDVXP9qCpNF
6JZc0OmdjRfwlPn5tFkcJY7pkekHiwmzL/pAA1VKhj/HQOrjGuF36heZIRQvM/IEbphNk0XNxj8E
OtFIPNYu27Bp96NJ5+BQe+/P/rbIGlmUvhAN+mAv7EHttvmEQt6ZJz3Gvu0ln+U+7i2n4fOPkjvl
+GGmBlaGarWGcTrVMQhi8nWFKBIw5gUL3WhOLagKOn4rwhRkcYUfpZmH+RccCEY3ZfCS/B4cOaDR
WEHHNtK4xt77E7+IomErWhzkDE8mW5h8uW/fj+brtGVm6XvQNuoYoTIruQf2Eztr3XaU9NnSzD0w
dJ95q/8waP6u4dmulmzg6Rvb9iqKzn2oXYUBjE5sJwfu3AcHIaHSMrk4SN9nMzM1j1STwm2pzDua
AWXaLfZstSCC5yfyD1yXoH8EJ66ehKe4KtS67TW4sHUkAnb8uuCj2Om3mILh7Ks9t9e0LO9YNU9k
+elLGDafW8KJVEGfAFHg2hqZ87h63nubfLbmAaweHN1sMqXtxYu+fkPQd9SLJ9rGzqI2cDp2o+59
HSGulRqedOJK4CLcN272z3eqaODi/iDXVbTEj2xUQGITmLm5mawYkyD8yHIUlLCrzzkSLBJ4t45Y
dxWY4hoIGt5TZ86lh8wmPp9fgHJQY1I27DpaTZgK6ZP5U3auF+00AaQCNNnp/U9Or9zaIn2lKYoq
6i2N5MGT0v3CTDk8gghQfLYFXqtcrD2IChDUSEFuUmnzV7OxWcHtlzr82jKuboHt0MGu8y9pThUa
TID4KqcE5E45U5kbo4iPijc6AjnJRy19J2E7vokS71lpnjxH3RMfplugj9V9JOTfOWEED/sHIbj8
uX6oYz3bir/jIOqYWlU88QddlVVg5QU+mjECk4Mp8Iy1N2cdBGom6cZuSzhSKZ29sjJbPbiRvN+E
z+Pwk1ZeDQ2e9y8DWNYZzWyBuywUAq+uKNfHn84TKcFMmWtDk20yZS186Og8dUx3E+Vhfms4U4GF
NH0j+0GNrKMUUKZ4NdG0hBUBpjuTB+9tkvQJz1TnBOOrtMUsCUD35mpBj6zOKxWlZPYwsPjMZ3og
ptdcpsCFaegVELOPYWZBwIvjmDRTjWtj5tx/DEOECRFnbQXEcPj3IjXimGxpqWuIcgPNxOmYftvj
jNkfHJoXdi5mWRAQZEIW43zk4y+gwT/lKOmL+AigC2TLT4nRQX4Ms07emCJyJPnmoFcn6S9M3tgF
HNrZWAtKuum+Xq7ei+vmGrb+42oA076kBf5bIbuRYnZLs+s09EHMQERZ8Pczf1gNM8qmNRiyG/oH
shW4n32Fn+sJnn7V5Lb1ig6QSv/tpzevNOgyGlBWq2u6R3k8JN5WtKWvBAzGv2DopH8kQmpJ9eJJ
X08Aor7K5LoZxe98LzZKxuYYPMSBEft9n7tKSehEAW5qOzRHTaC7mml9Q842QGiekpBhzfFBQ8sn
MdyPfGhn4lvyqCNNI+dJAx9ZrcNlpSC8f0o2OKmvOd0eBCpaiIdUSF7cIbtqJUqYl9hrcn/WJ4kx
tMlsfWiTpXvVi/jigOlegDLKbzRSUmi0hB+6jbzFuU+bALbRUL6wql/tK3SeAdLRHXzFU0n2+VRy
wo+xlpq700T0orEPmG0a8TfIXgR5P5t3/trsU4/F0hGM8ruJM+YUdllQTUsgVQCp1v9X3xWDvAzS
MutBtnC71HzJGIKUfEoeLkGLvogi9JBEIqKOV0DbjsfVxH5oKLftHRuorb2QWMshkfcKhYxT5v+4
h4qHAElVyBWnKFLWccBxslNOtDmw0X7He7qWyrLe9CR8QQxtp9Je3sfNsKxKcJQL6dQkMf4hKCsV
JMMOd2efhXtbkl3+iu6CcU7YcJhP8fw51szUzjb/p4SAAF+uLvyeACCyDp/kp3asyjrAnPzkk8Uc
rl9Hp2Dfo4Ba3M+5Blx58ySFh4zVKbSOMSoPzITOCpM+TOn/GMhB3BukadWQoZF+PYwphibWG3M5
LtDy3ywawlLLHqqER67Phqphs8iWZdv8JZmod+X56UXrS5csYu1BAwS7vXf429hUfUe50pPe0X3C
I61jtDMvbraZOGxIM0+EwtXYEuq5A90hH4yceQahLP/VZrZ5o7qSHeNmJFWGitVEBkt1h6BVhnos
GyuNQC90DNR5JRos6DrhkBh7rgS1E1OCKtV578UByYJOVenjh44R737+30P4sSf6xpIviz6Cze+9
1F5WZNYHOK38D1pH2aCY0sOcQLOuVG5Y8YW7jA/il2KViSUio6hbDbAl22TKbC8ZCxfL9HZ722WN
Pj4JskR46po86nXuOYHqg14hCzDzQRH1obXSCIN7XO1P8HafHwgRx4ZmSXVu0Sj7GefLQCjn6Kmy
NJiFKK9gWj6Y6CERPRC4eCTzwOL4vu/2tyLp3x5dttme3u2WAfG/D5BdI7ErT3VUfSbT5CnD4H0a
/KAZceiC0Sx2Ek7CBPSI6+BlaJV/+t8awXMs+yG28/876TdlWvDXV2sIbE3h/J13yX59xLOK2MZC
OQhYA51zdcJQwhJCzJX+s03NENQwulF4pgVEV7f1zPCBQ9+XnuMxswJJC1fvwt4bsSIaCaU0roSZ
e03VdjRiKkW0/7lsHQOe3TXiAbl2gVObTL8w0kWKmBOrLf4piPYpK0AnGwYZzi/YEdr15t2YoLnO
25NULMhyN9kFp7v1xlwNfSGxZPoO6Toi1SqMBuLa6dokWTz4IWt2l6kp5jfZLGKtNwJ/M5AIHgu+
Dih6wsuOZbkGO4t6+uE3h9ug5AKNOeQQAb+FNu80b45eBzb/ejtPFKKOJ9ojutw7E5djEZghvU1g
UsLwldryFrNp+WRcRwSk26mra2BjUfuTI7FUEVTDspXvPcQTpolblJRJ3hM182629pjlLahG996y
M5l4RV9xWD01+ZX1u0vAU5+ekf8wfrdYHfkePIAb7JSXv48FkzihBSrerHCfxpJdPPqbhn99Uruc
x5MzZJyoKr2BGYyS9tEB7pjaJJNNyz5VLixN+T5O3ZFvjy1CUVR0KOB9wg0QPBdGMWi95dtZVq9Z
UQ8NF8hacS0lZfvdL3oXvoWEFqo2VkowVppa57CkJqW6Su9x1SHNeDuhXE67/cYyuHpYcvoUKa4r
UG7X04hhPvMPM6E8rERwThruvHRNa1tWX/EKoUB/oKhgpXFRbgc8+KJT7q3ONwuYgPhaA+w/EH+S
eSQgWJvWfJrBA415g3pLOulWuXm0oWd+pXbBsve4nfmIxue/sppcDEMmZaPQb4Wdy96GBTPb11GY
ZoZYiZsRNWLrjPTUSoP18SxonjjWJu4+8QrmTFKPWFeaCo/3e+W+veuU9ZMunnviOejzOqYn6PT/
2d1z8lA2/XCkLaiodjzf8py7USc75JyRRwIcglAlUgnN1/QIF9SrrdH1PEapEu6gYsjTVW9VkPHH
Bf/5cRCRIwtSOR8nq2aRfSUUZl6yngfkGrX3lBI8godyImBdagDE5L8RipK+nVbahAerVcPMLYFR
pnauEGrnThrQFEso4vqYy7BewXd7/NSNA5xsu6lCHnDgpTcQJrkn0WIbZfSNcH3ufJXI3qodLU5s
e5a6qkfxwhImkA0DhmMXt0ffRzHjrUPc7cMarMA9VhFSwT8PN34l0C9syQx+HkCb4tzakI7R7VtE
SzcC+tvqOGs0W3C9ZN/a8FPP0M26QPhevySCQI1J5mkErO+0OpyDD8SbEyctIgoZPW4ebLHO5ZvR
BYeeeW6UmNgTnlLtXIwlmVQx3pe/h1qAUTKmwimYjO59RWYQRsuSCD2H58EbsYpyMr3oPeAjOPBI
A/+dTaGAxYSTDZkbxcU1p47w5TF7Iy8fNoOzr2JUss02Gb3vM/+xxSz+fKEhqXnv41liowpgH7qc
doGbNxKZwS4tW9rAUZlMv3aLL+zRs8LkfembTg0tZnWQq0luTvRjYM4oz01JDDzg33rCKdoOktwM
KgowkE1cRtnd54b2/qb1hBa9Vjsex6KqY4Y/gm5O9v8ipK6hoI4SnIW2ZF9QFD39Oq3wTGANEIm+
fkgCSVHGnmhw9JYknivfvABrAUKvn0rgjqj8QpaXjJKOkN1haVmxyI90+iMMis7CAPahiM3eY+Ec
pp42jPZJDnk1muGiYqbdIG7R3iSY77MohD4ZFFeWDjMvLaBrwzMn8b/X6yeDTKGq/Wi67EVeGrRq
qeQWCfyf1d/0zUhkjSFSpog3rtCj8LgWCIjuxaCdZ1UuF3toYaMVf3AsRmXg8nDMZrm43mKiLd8H
PIkbm2zKbi/ENyHW1wU59wW1KLq3lbcydA6llP0sFo1SJgMRtRwQWPyQt+jhNQolKAtlaKIasy91
YGtSebqkMWR6XG2omNVq28zFeEJzPdbMpWr3MTbiDQpAG9m4HHboyJeo/tE72NrV0Bq7uRBdKvJF
05G+jKTCGTGFt3m751du1u4I/Wxw01/LjmlfbZ9AsXyRHEJwZeAiBzPs1mCk8aAPbKks0QexIZbu
KN6p+DW1ksWxoG8H54LvZO0Wkqhihfwc0qFpoSiSCLl78XvyPzUmnNVMoGD+Rs3a5ZI5cEDCzP9T
C26RMfRJ4d9haeegKPZRMshbSKsHcAlbkaGcPNS5SX8OipcCWVt05h2ugIZG+8dTi1ifH7I/RiXB
URX4+RIuBzS2XU82zKUiWIARwFbVyjSOw+hCAlIZh7/BnEsqU5pYedcmuD0wgFyBghl4+NVFt67e
u3oAFGwnjiIei21whjForTtuG0gFoyEiDn1xd9gt+fxWkqQlew0rCcpxgMxjYMZNAw89jGa9vW65
1mjzYIp1AbuLLxV/OaGr5MuXSUgIRYNwGpoBtfyOI7L0Ssj/bz9N/rTt9rp8Id3c7XAv1EvUlTmP
XT9EPUPq9Oansd9iW+vGbO4B6I8XYAKBHVsHKhh71GVpcMJB6/RxofYqSIYSuHTioq0xL1lTkX4Z
E29tbc5fZUH7gw8faGG0UxeJ3sQT8cLxt3XftF2XQZWrMdAWeAvikocMeLm4oiERYFozn3Xrte2H
gSGhjiIOMzo+n1lgRWpy5XbkOqPejnK7mD2bLQ18TLluUTboNJjwxS5Q2jk1CJ5tCDkZcKGWGN/X
njTdB0nVUCxxqmGyME49WtQRN1d672HsQ/+qdQy7eR1koOzzQlPq0Of/pxeMlmSgvNYNTOeSRBMT
PhbIUKYlyC4xRRkqTLsdmL3c2ZIFaoVVv4rf5mXE/VpZ0KFGJg7W3m1xSLWJS+StR5S0p4Al5XO7
z3Gl7DkgsFUr87mrAmsDSEk7DIVf+7J+1RKg45ZhM6Up5X8NM6xtWNOIDGYVvvmLDgAPCebu8D9B
ciGvYLgaFf01wofdDZQyY52svoBRTGh3Bb2v0g7g27cAR+xaKPsP0vTS54BlTckDUGGSceL2/uKe
TvYzwOqk1Ndsrf23p8FpTJpXJMy9e+YMBU2eSwt81y8Zc2k9OtZsACq9/VkLolRlqMo8cSJpI+iH
+EClJBPxMD0wmJAXPcLvP5fGMVfAAFpBs82iO0M5o5eQHbttrLUWo1VQF+asjT6pseJO7rgWpEUH
lqA2ewtVFlOMmVMzkfeS0EHb1IljwBgUY3aJtBeph3ZhCKMXrEIXRvaGcTu169AoKE+H7USKFDJA
XQUkAe137hclhe6WJfH+tzYq468LQrktZ2afFKDqkiYpiptfiRlwzU8aMtifGmqBUwIxiBox0tl8
DLp5PWHObOgU//R0Hlnw+p4Zn9vAA9rGEaCnSYjTDlpGziD1IvprXJnMgjiukHmp7sJIcPEyTa9T
nj56r8zKtmIRP2c1gttcwo0IoJSPk2dcicxM9wsRZ1LJ7FyM8pnnpKTaU6BmgZlHxTsM/pC2IFvs
V0J5xWMzP1saX/TdDlD4c/eRpCJRTVsi40Ol4G9gwjmQgEkVtFbggMjVg/gneAlYfqTtuZoeYSTa
5Eoq9n2UNuFms00PAvtTz7Qd/1nkymBAeO6UQPYa8vbLSSkrD5+bQl2kTq2aq9ZWXGLmDUEX9xqT
k1HB1Qd1gMHnLeRW8FNKI9ndnDG6Xspm2bMYn6lZjqgt2JtHse2IU85AgPZFoe4sKvNVw7p7boNb
8wZrsSxILwlpPU5Lhmo+CO69PirlOH9IPl48bszhQNmOcYeJGCxh1c5DEJHYlRo9jfdC7RRUCB1z
JriJ0rakcTPaqWVLDXnQKC25gjp3gZXq4llaNrH7k2m42eFC6uBRy430YcrYqxSBSm+0OFdv4WuO
8qBWPOlOUznojGTOFje59VwGQshn7moTGrEPS8oG6XIhY1xQtBCxhBEE/nBKExFOFhHJ5nNBVnz9
SGixxyT3IAHqYnQw2WeQn0jj0W5V/sWSMjkWogDIpInWi10qRS4jx7WkOaUVDCEn76emiu9iY2s+
24ccbAScfPysTtDGKMvQfQpHbvF/jw4MEvspTOXPYU9nma+/GdzwGTKknrz2sVfzcSoI3DNZzsAw
CqNEgz5g0jjapI3GXjbpNAJc6b/M5t73/gkxPi2XG1bKSGdAhHrM7qOsvOsMkpm17L7buDnWCxNB
kL7OM6mI2Z73jGpPH4XGj/G/tMHjwZEkbsmv52relBybYvVOWoCRi1XJB8/YU5ISDrvvXdE/QKl/
pvUyNZ8P08pKTZTj2VIlOoiHeBGMweMV0K5kZCRngGZ0uCN98Lfo4W++RSNed/ymrXrsZQ45GZ8q
B11yUawev56cJXuU2NS5jdyXor9QJsgauSzzOLcW8U3chP4fVY6JB1MeS82U0BdMgbOBIYXCWaJ6
P8Qp1mYbGLIJMUHATS7hjlT69+Hx0ea8OzePt9sduNOLefvIn6f5JF+ytscBEPrVUFHLRcqkQWlM
VABOaawzqvprpheLnpqeonKnIk31cIQyFGxue6XfMjKlLftJ4KvKq4AaOxbJ5rKEVoZL7a1Xbyef
a0h6KDVtCpEgo0+9X1sRkTtIERc8kFoROvyM+IHBFV00sJN3nBANGtGrLlzt7wVjW8p1EHmb9pnD
8+h6jkzCzCo9EBq/Kcah0PmBBnBftA9NGYvyCz6cIx0nYrJke5Tu15yA9dRm2PGIib+kJdvvyeJX
G+68eEqAfD+IYaKWoWdJ5sPfL7GxnX7XMDPP9zdXymupgW+RTvb2rY6Qv2foKcbSIeby2VClD4wR
eubBQgoyYBKR6I1iiUWRGY4kQ/N7/vl3cKc1tP7VrZwOb/NxNE1+A7cbFUCmEmzK0mwaeLqBV4wV
SMhUS36lU/t5pVX3iAMYHPQdkpCX/KkcHS6V6dQNBN2oN2po/j7a0/VpbUmgMarxsa61ac7W91JJ
Xf5QmhFjvj+j0to9aB0th0WhqFJt6uGLC+WZpr1tOVsgs+GDGu68SWVx4tod7Pf56fJPEgH4eGaX
innWBYW+5Y66xNDn8fKmclsUpEf9mCPc8PYjnhIm7rEfHUv/OB0mjY1lvjkn31mcj7g9K7bVH5Zq
2cTi5WD8p5RL7Q9my/wcUD841n+938NOw0rns/pturoJmCzka4MeqAGFFjkGc1Eb7sL3tBOxIt0C
t8kuKzthBGnr/TklG4L7tmHUj/ZZYF9ZnrcuI2znIZk5SS+LRIj0Cmv953rcZzR+RddJh0HiLA1K
9Z7enkhKGXOrXLZelNJ1i4Ft9+MO19zqagwW++iMlOYE9HXtRUiG83IQvGmRkkRQ+WbjpuUbL1ms
nushNdYt+XN49ohHMmaV26WnSa52XCxIWRqq1a0sh2gmyfLh2utGGkwGVM/mNtTxB/wiI0n5NoUA
lVAaJ/m2lHlw26hpCgktTxAJ04uwBbd65sephuOLsFhSuWVTVY0F6Hwvo5k/adOm4vvaQaXa3Gm0
2SigdsZmz2xK1/NAioC/Re4aswGwEQdLACUjVMbonkMJc5BhkldUUVc4PiL5gwVxdW4ET+E3CZob
nLPqQG5xOV9q2YKG0+3VsCqQQ7IGvwqx98UJzLm/b+0ltxsNhstM3EdjFgqtPmUuHruOYNqJAh4f
FYrsd5BfDv4ZYw0vz96GFCDE9iWJl+ZxLVImTi8hfkjRc6fUi3mz3CFb4EX9VWqMuDdp7WfRijNF
Od1gl0sq5gePUiGlBY8JtIMulx2thaAK3gLWiOdo897ibYTDCllwVADtaLsZMbobAMPQVE0bNwMz
Q/HnSqzMJ/XNzKO+S+tzUJMl+DXlNClcFRK4A7dx+ivXF9nAz3s90RLTeJfwap6hr2f4Ht5UZgC2
0uHckR3wSA7+LfS7bo6dL6RfJKPqKgemjWMkVZhjQsQwX1zCnPATHPiIO4Bd5prsOTT9fuzrDs/V
2x3MstypOKWy9khX30Y9tzdYeo/qBAgHCodEdComrOEY8eiysW0CvHloJiQefDxe+EB6ylDy9hyD
OVRLKHI4Vy07WN06o/59A7znrEGrpKRk/fkfj8Q44/LZ24/NdDo8oIFCfXPjmEgH+tH/U8Y1x92V
b+kRe6kKc7UZh5gdhXzlCwitmA5iqP2nmQBmmt07NjZbOl5VI6+ZGWtugGPKjcwnDkLl2xAHhB9n
6fPS0WzIYRmDCuZf7sJcyAp1H3geIaTxFUe1F5ZP9OdHrTjBkoxgPg4dA6ph7DMYxlwXgB3BDrp8
OxFLkgygL46EN+fHCDkbpkrYoydW268XHx9UF95o1naj6L9+sBCo6rWzo+PafHt13bkCEij9cM95
I22iFiloImhCgCVQ1ml3iYLrlP0fTMj3hSRf+79pXAD7C+fh6oKIyMqWc9jxePEHvOOv/l8arlfB
5vS8+m9Niy4tt9tiGnivHfOa9yGKGb1RWTEGMgfHXXHqVy0wfa89dqIEn4rW/9G81E9FwPS8WxQ9
4HCbmLe5LA5v7KKyJoIl2SfL28Y+BpgDjJkoWsRvJjSHO0qEXqYmdQCTo5N3PbwoAg9+9gEVuhKj
zg0o4eW+pf0zHTLoI3LltJfo2o78gwvHS7Gwz7jIKkLUCq4r7esV6Nm9MQy3ZLnJH+wdLfmCNOzk
lmixppEVxk1WLiyaedYhgGV73MKerYEmUarIruVTNakzvma3Tir4uNhA2Kt6gleONYcd9Ezo0a5O
8aDKifkHWrCJLMMIwCo+UcLPQ/mDTkBqsLj4Z8f5ZGZqLURlQnKl5lV7UeH9akJxSVrUdIcaaRYV
+sxLcU/EO9n6WwL/HOMWRM3VKLzSp7FvLMvytHgFUeC3GFhilD2IUmdJdXdnj71ubqPzdO43+I/8
FocarcBQrkG2o0GB4rPdFY/xoyQL4mzYQdTA/bnvqJzEvUVMBFjMubGgH0cR2EdH3XRBMzmTkrpV
tnu3eKRMQNCRfbsiORz3+MBGDTNnrox82PK3oW9v6WEu8eb/TejHwHdtKI4+fjUgWrpyibg+XknI
T0KWMvsm62JJXbluz1PjBeZZkrqD/4f61A+nzo0LO4AVl+CmeM/UWzbNrip0Xm7lzM724tLWG820
lw/3qii39h5qiyn/rbzJeUuHOE0xgFvETKjk7Y7SXAQjs69KtnFQRj0USUMkt0MxCKKnXxgjWguN
ZRfmJN6UMcqpTbKHgnoZ3p8eMVUb2UsY5KFb3VUoTlOHM8ziA6a3i08DqPJrxwSa/7XHcdZrcg+D
mvzUiYNGsnYtvzH03tlT2qCdIIz4+rG5K8ZFeqoWJgIjaoF4T+s26xduKn9K2D9jDhIX2ZkOu3Fx
ZBjlXuXC9NFup7pYCfTW79xPOF86hceq9QLpuKRfTx0L6XiGIJSoGiPDkqch1/pSiekFgdUljtMP
tn5EsWpB/zJeTzm5XmUfgYotJajQBB3Kz158hDvjMHdMPAZdJTPb/wk7Gj7UEsOtSjpjnPjqZCjF
PrFHCisFkOqD+Wy0QWWUgXygkbi9omeJMWOZcCDuQ4fKg2ghgzRiMA9Rh6rwM8ssq1hKdkpCU6x8
MeqnaHu1BNiHV8YCNv0/YgpeIGu1IzIAmQVuBVQVEf5aRUu71Ll+WPnSw6Fb53f/K4f+Tg3xuChB
fSgjvKnaKcNph7DERAM6ML2j+E/ghbjxPdppvEjPV6kMCAQN6ZvUA+/OHdYIxGNdFqzSNraii+iz
A9KujYEe9lLUGTn3Zk6/kXECvIDwv+bkIqtrxffp5CLX4kyJyka5aXagVqmSaIZcrG8nUw6xqSnY
PrEPm3kR1Bvz1n/a+LH2xktJ7SSTIKfaOD4TaDmAYXOrwZde1r+0wdDg0P0TSqydddnXRTipikSS
mLy87oxyMQJ51w/LBxz1K9zJYKuRu476eKJFboTU2lQCpEx3I/1VS7yMDmCookpxoWxVYEpxpyoh
nsmbs4QgiOEz1GYJ+HQBYigtn5ttesIphTPN9MJoTDwOyiA1sCvdOohAXMpI1xeIL45eCCKcpee2
fs+f/FZsKlRHrQbQzO5yfe8xSNP5epkqRiSsDcDxPgfOGKWz1XLv16QeI/n7nW7DQOW294X24fh0
z6Pe0S6DhrEPwKDkyYkctf6ZBaH221Zn7m2EqB2vN3LItnLmkDfwbpg4g+faxWoPAqKPdEEI9yHS
LAWs1A6JIyrLCkhpoz9+02synqu3NOtCQP8DU91UfrJGOmaN56Go7htBUQW7IYKvsASBdUavW+hv
igliSIPYotAwKeS5mgbGglW5hDQTEzhnw2gnjwuqBHakPz8TdLtL3Txu48DevhZuOFg1JAGJxNf8
+XuZUQrd7sD9wmK4+yCgk+A3nDGIg6N4dyUqN11NFh+ezmt8z7ASfdTorUAAvCYGddO3QpX7RKvx
4oB0XFJWspXxJFwtcHPtpr3oargfUmimEhIPtZQBBybbLc/WL3EpdxM3nCA3zlxt2sZfyOtqh9Cv
UIxnd/HjqeX4FIiJgX/mdw5u5rWV3TJAQI9mPOEU4ZGDzpjC7dUPtMAmGuY3Ud0nxWr/JRS0IQ0H
8CwToG1f886bh0mywcQLrkex1ogctDnofZ3100V0zN6roalk0+sLC9D8siJXQcYros56et9XH3Z8
ZVudO2dF30V52WdPAYJSyD1tw86iS3Fs+X8n+8hggVX9kJYnvEjlMAmBGe9Ia5dyhqf9gkUzDuMM
W6mWHZHZOB410xBLjHqj6qRj8qVd9TOlj+KaOJ4ckuS5oE0S3Xuh2YbuoKXnf+u3imq5O5gS23Wf
6oIlt6rbt+Iude2Q7dWM5p/Q+Hv0H1vfzjYQxm57IOXwd7DQMbEFh4FaaQnX9gZA9XBguzuotubh
wwQJGiM0JsPKy3hLzGKgCpjcGsh7wHoMpqc2JAvNoMMneLify1IOrmZT3WZIepq0kwXHt5PlpS0a
xvJhEHAS4aBzb8cqTPX0I8r1nOQE9rDEWJwRlkQEXaY4J3Bjg21An1WSj0JGLQkWSJzM+eNKpS4R
CUl+W6XywK9u3JeGq+AJkBV5lE7KcO4Xgfq9X6JHlSSkBuGs407sHLYi0cHLAtxY+C5PVD7SfDlt
32GXWhC0kfzNBQeO1vhv8lBGX3uk2+e6l90R+XqkSoouJUXwq4fvHgjvzMTQHM/DZ+bEzEL+g+us
3WPNTQoCEi4zHQkub8Mk8xscE+SFbM2jXcr7aD0SyXw+UtPFRO5zAbv2IyDagp4ZSKXIqMi+cWKY
M8yjBGh2XenuYuS8B8+Tz3Hz5S0nwpsiBSSnYNfGlWWNeh+W8t79oO2InAhwKhlD+kVp7oAoWBk3
Kwx63DrN057xYuW3aUITz/03k+QYsZ9ICXifXy3y4AlHLgM6iYWMhgwwomK7AFIfyYiB0wNTvK6l
F//i6v00CcADpskFEXpWoTHqkT9mdudjlxJVrDgr7nXEVw1nuIyOdSoIAOOjpALb/gIlurhW8Daz
/AievgiiQN98rzD/qu5B4Kdx3cNYo85Uv9THL+dxpubhKT9RRGnOHhlcFwXbHlGX4BRryn7aJjaJ
Nduxhqs47BfaGCo8cU7wsmDABKGAX9HZSG3d3Dy2/UkegJR+o5JKLCOelVa77Q01bRvWAVuiiIiq
w0owKkTmjs8L+lj5D8DHIFNfmXl/QXGiANpoZx0dYp62c+9xyV8JlLDfJItmkOZWz376QR9xbI36
G9JRMElp2zey9M9Ps8YiiHQybUf2FZgHuGyKNPm1PHvj1X4/SE2dNVgLAt9wLN763H4dBE2DDp5U
/tidGGJ8OIdnFF4uqrM+Z2F3zj8iQhGsYDdOl5vRu9U/k/zmgjZuW9Kev9OFUIUj1z46u8HZfq02
kv/gX5omcucoUW2vPuVaQ9mOxS5Vc7lh5wrhxms+Xml34IrtV8rDZoUnkPR6bX8h8GSvTPcRGWHD
hL3QEFBFVafLGWY4deIo+NeZd9TL9CQ01htvGl59U6SFMge1zuFJiZlgSdfOF4gT0WH43SqYwy6M
RaTdaamQoLh8FWvbw3+EefQEUf+CQfQEBaKjQJa9R7rbPVC2OdSW4J8ZzsIQdqzHa1G7PHTyl0Vz
8QZD0z8ITMDDuIbc3om93pwB5lsiJvFVnAbArIzEJKqG+BGxb++LQpDl77b26uTq94mHGRyReOLM
uKkCyFlDK1AvAy4McpxX8gK1dP5//coEfF8OaOv4/Fza52kqUNME9UPGGUf4nf4GvQufzMO4Dx6e
6MJh4ztRXtPQpiaIXvekZkfyQ9WcetzQPXKJ5dlmQu7PMmmLrCecUZP/669FWWq87DjJ/SxtNDyT
ATKo30XgLEWEPof2IQpSk4ilNQWeit4PrO49QcIWJjsZOF7xhXZwDd5oEYcj3XksPdgubkcHa/h8
UzvNc21K6vNpbPtD21QQ3eGBVWyt7ydxMbhQlmwEOegE8xwvlb40TRBIvy1Ooctk0RI0Xmfno2p9
QtdLtTPkHsmx2NzBLhL0YHSJjT7hhYYF/gJHr1Xi342CFa9c65gb3eFGze6Cip/Swn/YGuoVxPBq
BYUSNNGqEdJzbOzPxJ0rUUEJdoS5yB43QyIfXLSzUfSZg9IQRauWgBYuHC8wEnY7J3LptDX5YEvY
5Z0h2Cvy1u2LhJNGZyjboN0dno6QUv6JUd5i7kJ2OOWLNrG0mvkF5w28klRpgZajzGKOFZNOa6VV
FLKBXKmbfrNsnSIkN5xWxzd2/D5so9XHE10UfxIic4E1s5fCLkuG0cY0eNgwUNJ7nx63chPpz3SE
T9IV6nUWKWbDiPwGXlRMr1hoKzexfCGqUSzzy+D0M3GarGFSfySujnpQsNddUv8R/TSI0VHGIZd8
2X8gKJ5XeIGisOHm7xiufV4HGge/5x65JcpHuip6eRnHcb3eP1cr+D80YJqrXj764ABwdPXX/c7h
iUvueW+yo1D9lmbUV2sEcUMg+4gW7BS8vKU4xhzuhFE0FSVb/UsD7s/JBhAOpIy7q39mjTchcaHd
hF6Mgak6CqRpJC22XXZxPKwk9d3+JkG7M9DWeMNdLkPYQAuhbvrsk6GnHr/O9C8ZnRw3WYADfinh
E/BK9KSchPqU4+uve+W6atekgF4xDjFX824AiVXycvXiSuz7P8ue6fkD6aP1KQVRaeLCSnr6dcre
lqfQDZ099MstPAb0fSrRO7E58dQVRESg8u4AEJv7F6nREC5gFSsRxRBt8n3DKBa5PqEdqHtFNX+m
l8/0aTHp00YVwCCFaVkPlx2dxXMUIqdqznpDZfb+3yJCKbP7XsfZGqR0Y1N6fifv8CN15za31mlF
7RIXfMT1Y0AZix8p9MLsyc/UfJ+WzD3KNFKZZKL6uN6EDiW/b5AXhth1CR5nUGLkgCpXiIcAFJvc
TTIUYTRZpP05vwLnCp7Q3905gjkQyIEQwv5bxkWiscjzrCydHqm/VxUz5832JR68bLWAFa9LC3d7
b1n5vbtKo2+dQnWeR+nGUoZJTuMXaqJRofpwuoQo6Kg+uDkZNtKJ8MXpGJFlG7oq7T3l3clO/jx8
uqNpGnWdyXrp3GmmIG0C7sWtjn7hBd20s8Ur7rxnohx4CZ95PPgvnfRzr/8hFbTDGJFPJ0K8MK1X
JUeCNjzz63FcXV1S8YPPbAsri5HDpK2WOYfjpqMC/Ye9YlDN7jCbZ7kW/Z1ASWh/8xWVfwj8PNgy
Fk9DggTeAnu4uAh9boAM+v2mrzwYeKUnqSIJvFGpUwDQ7Ol8R+zxhW0czh7eTRmcMaRM10R0Hn+/
4w+R6kqNMBz3gwmSRzx2FYCA3SkwiWu7sVAm+bw0jB1doxclOz1oLVjIioHWqhMOirKio8Nh/+mN
/1NuEBwsJSQ36XmwExxLdhoPGIKIGaVPXrVgFOfc3VmOoeTDNfHVYqToq+2uaXW0CHtyLRLy3SvI
qYPFsjybLGQM7MSBUDMJHw8T/rCEAMy718rr1M+efnSuplED1R8GtxDT5U4Yw22bmJ/TGBGH4pMN
XGLaScmRC9fCe0csOC2kx+u1ptEzdwTLip60fPtnnpPuTzffhhOtVO7GvFkGHSKhhDT/JoEw1P0w
oItuup3TMKTFAV/TOVx2xdI6JGZOM8EWf2nu+RDuKnm0JXi/ysVBQF1wrrgsJITU36+bMBZ21R6h
aK4wCTNb05FT5XNQYhSLUGYo+Wr0SI0FYUAtOhSSdNvRurRObmyBS8/FZ2zv4Em8ea5fqUlBXo6k
fPzPO7/dg9ToxqQ5MUOtG/Dp7Buk9GbbJqBmRbyQXZZtr3ayBT5czCsVZeN6JXHUtv1AzO0rYVth
S8I0eaUYry0jNj8MfRN9ymMTgI/uE+UkCu2AqISs/m1GaAtq5yqBmGK3bDv1HsHN5NoJOnOkT6Qm
EyD85JYMbI8kRioorBIyPvrjpFcFt7s2N3AmNklkyk4WI4OtTJkkxoNqD8MXp2QudKVDkDroxPVT
Kh0uer+jEHRXDUpvv/J579a2oibC4uiClBW7ChM3tNkXlvhmXi0N3SiQufBqeLLDmkRovkE4KCNo
HU2iCXYHz2qZQdqddgKH0mG2DNVhHkZYrTOBB+QOD+tGlx7oL9fXSBP/zdBzl5pTUWrpjZ6VgEs4
3uC50AVPPPnqrvKnRuzyTknqjxIVfm2ebfimFBbqGz0JT96XmsrCLl6qrFyFwKbYxIj1/K3oUsXQ
Vr5GK2ZzJhCaNz3jjLsSzmFJ5bVziFZWkVy1O4mkWlCFmmzEBmCEXlp9X98+cCHikl+Y6q0oUqog
qN3nCATYaOEEG1+/8soyHXHqb5vx0ApirpzjZe7hTRqVvH4KVbejrrL6AB9je88WgT/RBbnkCM17
b+ZSMZOci7yR7W3vO8ZbU+3bpxmySflMLCD0q5/CeTZKF7Ott5X0rh9pSJDXuv9OLyAbAbtXKeok
XzLFeG1Ix7YDvTzvw3R91ixSLoLwf4dUmvyNbYFcIlbNfMaGpKOG1e1aAj5r0kVkXE+6nUucm2Y5
6PeBxDoyp53fSfMULBBuvCU9D5XlXTZgYPhfU6oeiKz7JrqgyYApWg4EywSZqULXK+2fQlOMgiKg
Wz8/e+SmEHTMvF3ReSUyg8R/1p55mKLxRB0kRRBHzO/KVCoCJ2Anm/VyCtQLJ/K1nnBorMcizZWf
lB26+xe+6lgKFSek5Wz3h/z/kCvSPZJu1Hk2K9YvmW0IwNdrnWDLd0WTUp166qq9ZJEQfZptShX3
76PKqknqiUg3tfeBEvSobhB32YDihiwqiCujk2ABINbZPRmGvrRoK7Xt5ccSHJg+5Y98Dg6jUZrb
ANsnHvmvevREQzro6xm1e6eq80erxZj2YNIBN7atG44Orr2JJBcu4RLOlSOyB4NCOjepbM/hUKQR
gYnAcouF1vFXeSR1rJSmfzk5ExIAukx4Y7cp41LUa3T/IyKnJlGgpHuoeBsioTUzCG1fbnhvkTUM
oQJytRrT4dhhRgx9LMl9b4sZ5VzDKIw3L5KIxXSOZuylUGs/CZSJj24i8Qgmd48hDNLT/hZTfzb9
rp1sd8/wP+lzkwsWzyh1m5pVy0nphG4tJrhZ6+XQcSVDkqln61Xa/Dl6Ez8ZFJOll01xuIS/y4xl
whexWT1xVUJBW9p+XZunnY9dVX5GrD/s1iXsmpD9KVb45q5DN31gk4raa7qINh8bjjelINPmjJhf
fKGvgAOoMV6hqVr9AG1FpataeKqzg5tx0HxEVzensS1QImX0LnnKr0jXeQEZ8Btek0h9dIze1iad
FCPPxYNEQ6PDMLksFZd2peg6LHN+VyUU05S5sSS7UCl4g7+hUE5kelGzj8lFEhpGtdUhZOJiE/gB
jQ0oZdD0Zo5sHylZWxkKpE69+ez+QJ1DussbMwMOL5TRsgjTsaS7b4VRbxxpe6r+JiqdNofd+t47
kDWaxzW6RTKX/W36UMgxnq9hCSICLbhqpm14xkNJJlpPzbnPAKg+CS8kD71NPu6KugvGx1IBuUZr
s7cm1h3Qk395wi73t7bGq/jZ0Afybstspxll3k2XOfZaxrhnHBG/wphFdM43uur1lcPQZjjXGg2k
deGZe9C7eZelctBG4Dwy7ZV2HNhcDHt9j7FJMaTAjRCGSv2wWFlBwgRlIhy0D4vGzuhnUSgfq0cf
obBcCPuN1qI7aU7bSgrjH1Pb8ztk/9Ly3RSNhIRrzYRb1SlRIwEqweYTR/HB5mxq0dBJV1/tr926
Z5VMRAaPLWC3SQGVuMiRmLfXnSxCbH37JrlGpWP4Re212Eh0N5bgaXEWbvrV+ZRQTD9ws9+NbDTH
1I3HPXOtznSFnSmNwkzlJzP2EB7WpFHS51obnMK8rt89M/5FR1Ix21P+xiYa2GBXTMxjqAgh76Mn
aXycXOvzQRMo/gXH7igRL6clyyGPVLL1KHUO2aG/79QjcMrO+3NbdMKJYhMa4dnapLyipWsHo0TV
PPZ/FDZqEjHpropN3FXoSzEnqCHSU+FZC7K9lmUfghEjw7wPMTDVBV+rkXfdPelnmTOc+w4gYOG+
lvB84BpQaM9TaAyf5B2/ZkfdRjN6wN2DGoyEkTfFfrNVPjmjx/HQ1BBD6jYXD5p8vsOFKjJEQWBQ
V2YvwK5jv+XgrF7QRj1WkZeFEfsaTOVowKIvpCDUYPfdxaQIiGSWOrWmgRfgSYL4AYUdOh2dzwsN
Nc2JqwFwXou59c21BcZm2amkblA7kkkculium9dC9evAN37ti6nxIWUZBYGamrB1kxkwoU+MytUp
ZRijecEUnIK09qcCyW+EzputMG/efWbRf+mKAqO8A0kdU1dTS0TBfl2E8ayA14KsXqkkjHstGf3E
oBpIxOMw9IpAP5iuUFJMiopBuykUmn4sBZkbeJVcpiNkXo3HmKv/eBNjNrH/77BH3PHuyYDYkVdf
0/bw/J5MN4wEWBXsBXjPwxYdFMjrcNigRO2PI3zzh4IPF935A7CCKmVe69yjS64ofo6UVBjcnFTk
H1zRHAA/5qlFjev+0AKZk/vZf7nVR1ffiUwTnBDIhZqmnL2lVbOcyfSYfZmlFqrTbLbTmoK1bSoz
ovWVWA1k50Gd9d/uFEcA7Oannz3JDCj3Oe2GtUB87zuZa4cHpw3/I1VtykItet0p+hMk9Hzd9613
xAfigG6jCVn2Ec4/txEUJnKE9xmV6LpzuvzGWpFt3ppdAawFi9zXn8Rbs7a+ay40EMFTi5vI5KFd
eH+D1WfR84q+vedaktMVPCAa5tb4dBGqOD7jGFwqfmkh3SfHil/kT1AiMOBABvfJc3sWhLLBjtFg
fmy4kUsUvGCw4Q3j+XkQhlJ3kOXhME/VcR277VZ6k9XeoN/wqbXFgwS9YoyQHbUV4Uwi4fnFF4XO
XH/vlsZ4XpBGdPE2CMJtINvgfzI0YcMcFpOVGn14v/E7Kg4cOgjMhxLYzlZNCCpXOqX9/sxfyrCw
7YKaQJU612JCtmvKvkaprSGUNgIgKxMTmPjP32U9nhSpxddAKFUPvim/JAj+g7fcrOH09zlRgtBj
AhoaQ0iBplkAN59jst9MkTVlYBmrJl3YxIKWFnpc5ibl9QDIgcKqCSINv2H3koN0mC/W3Y+me1tQ
Q3LojE1nGKCIf2hcPJ8hQbPigGDFSaPLPQzCWdkg+mj/QwvBkOaKxlzVWWu8CWdI5pmd6aOQjS/Q
bW0kKiCOJpzzbhEEAb/IASNlYTv++qGW0QS9ut9BjOEe2pHHzx8Pd7mtwT+hRqgCaVMJVjBRwnwL
b4U1F7beNyYnTT8JpU6Sfh+edx1W1APP9n/8fw4U0hqb7SYabvI7jDcKKaPQOKZngA+XQ7+g0KLD
OMkTI7N0d/a0uz2ywnGOHkGv5jGoh3a//YTPl+PetNHljHnTFrHMQFNj1dsvUHEu1Fn/UIlGTDMW
Um82kb+qbQUfN77fi9jVO4imEgf4jOU6BAfvgmAba/CdcHxnhvxeP7RwzhwLRYyQ66Lf/OzvsmSX
GIUbLf5m1zICrrPlae7eMtakkEHt2orsY7xaVFSj1ILmjFub+Y63mJ1tFUWvioZYtuRiwuCIknuY
LQkp/QBB3ymz6fwW4EE/I/vIaMjve9eP0SQn9hmGz+mStDkSBDXgpuGkVowswOUwXEwqeZhrpPHT
MFk9zIcJWIRTZXVfMoPLLSsya3EFJODofRUNECBT61k7R32A3HnEkgfD/u60RNRzQ4ShCfVplRBb
5AYYgo0v5mSDDGICiR5Kma1xxDs+focReIw/HRbmpin+b9ovhdNmLHkeDtROtQ84higIEddaPul4
DXu8nIFNjbsQ0Fx5nOnVjeHkpcekFFM04/KtpTqYFpMHINr9Rzna0cI1xnYBsrxJu1mCapn73IXo
bSs7oWBhxsxVFT6MpElMvxc1PxQTvwdmHgE1mRwA3vCUAafHCSpzuurOr8Re8Cwa/Z+wlmlxakZZ
P98jNnG8ivkhtamU4Ee7aMC3eQcftBolOnKEVS1pIBFjCwITp4kmYaHCns85Ik9X0bvarljx3/Ip
hktot99zvFRrmz5CEWbzVqYnUYTN8CJ05oKDtR96VqKZyB+w6K6cmUCU1e492or8ZlZy/Jgk5tqO
+w03sYXvd3XGj3leSapadcHs9KYNBNxIzCKFSvyF5DLw1R4IEj70x3q//zNyPKk5unH1XqT0rcrq
+iqtQWMCnZOHgrmow9DyIOHbPMjPnBCJxiCQpM3XRWuNcyDBLoOAzC20ZBYH4hAxqY9Akqc4Al0G
gZk3N3omTqW0IvOJCQOrcpiesBKzIbme231EtEtlmzYMB0uwq51JB7fBhj17GAyIMICgqBo2USV9
5GG6S0xFYlcJRK9D9v8ABL2X7m5xtivC/CujtB/SwyiMPpLTuKuxyJ8pVKURvrDW8kIqYhv3ZVbA
MuSxA7jqP5Tv3mQciSe5FMBbAoq/5Htcm3inMBXWljd1hXQASSCiXYybb4efGq5q0he6qq9854Lq
pQmDAezZCxpkOHK1H8juesOp3nXf5yymRDbKRaIACZzGSeio6/FwAkq4eaVXKW2mz8Izi//RdMmp
CEBCmaEZDDc8YjWH9TWKZ6Wys91deGK/W0MTOx6yJZAEfYdVeooT++rSk/yQlDXiLe+fVBiaPkZr
3JodgLpnLsjIUdcCJEqjwqn70LW4Yc3Lhen3qSQ779/CWYCw/3RxNJkR/aR3ZUPWC1mOwVbbEq22
C/X4Qe9jNAsIXnbBmBT9uNLjEseKZn4dGvQdykWdNUFu4ahXc/1kJWpIkTnJfbxCPlOYNXrchW+Q
bRA1vb07pteYwOJyd66L1RA96SXh5CDxyZ//j1YyANy3OBDIvoeS4CdSHjNE8PtJJ9nLTWVCIgjg
2B9/+nh/Y8HdiDhvREyCEQK2U1jwpGkJNv17PhX3+J/G4FFrim+j6aL1QkF48rBK1P24DHHPrOQp
pEt27QDvIpShe53jneLq4ZUwNv1DjlAr3enhR5YnVT7PWGSURfNm4jHE88sJ55gxyj5PeLPrwK7n
WdEZpcJSaJRLif0ZE4CImxcD8Sjs+/RE7FNEpsMnCMchOGgdfqzVAZOYLYQfUMbRMJyD/br6zSp5
BCjqtFMubFi5mc8v3gWJRo5xueYXb5pWxAiE3t7NGiDx7s+2Thgfert0Qqhn66lNWWZPONTD1V2r
I4H0HhGGumd2DT38Wd9I0wQGWZ2QHnx6V/R4T2OGLl5QvBA13BV/5hSNBK/60GY8d531t1HSlqff
z61KE2oyJDPpj+p8TDLJb9rC4rRPBHMoUsNFd5YAqPH29SKBW3MaNaZ1I1fhW0kTxi+kTuqOS1RD
phZzGGAoZZ3octRtN+anA16kmPdhYtJDA58qi1KMd8TdyM8wwv/Ea2na/YK6ykJs/B30ajXvxi6U
pVQWulJIW2VUGBl8HtjGiXgn79C3dtyMBFNQsdAMjti09ZQpbz61o5fmDygKXSJX3DyVXPXRCSYV
d5JjZdDSGwSJ2+WYLWssH31YZD76Kv9plNcDF0HJUhGw99D/tA/0NYKWT2cufLBeWFcLpbB3/l/H
iNv6aGMsBairaamhubwn+thGQ2XglsEe6EUHw3KSJcvJRZIa/yh7WCZ630sqgvlnk/QKKcAzfAmj
tofL/slzloTBF4bk/7kYhYBzqVf1PzsWP41UdX6UM73aykhifAn6oiM4fAgovcYfJ70QsOnaQ6Vx
YM4QoFQ+Lw093Z97gqIYDEzABs4dy2+V4pP0Mj8gq47u0k/idqLzxt9pCMKiNS3JdFYsWAj0ZTZs
qPhd4RyoFcQ+1sgnNU4iil0H31b+4IUb25IcXmhpW1p1fm5uP8SeHQpbLJS1k79EmbIhDuRjJ1k1
SJ/aoencUzV4+Papv/ajhhqPsYp1D6OyoW+IDMSvwi4I/jpW1H9dRvnZLlOWijpjsttEOjJpbXtB
ZDOJLT78Wfdwp2Xryd025K0H0HEdGOGmSzonWj7etwSh0mSF7MKMVy23UjhJb+lQzIwKuTpKUd/A
dAgycADZNtb77ej7QytIY7yIDe9/CHuL/ggOWSQ69mcmvW4bgXQCfMjIkIgtn/2peufPNO2r7+sB
y0n2FFXLc8VHuOWnXb6UAYUGbAisFERKU7ugnT9yGx0R0Bmpn6/xp4BLnm457QG7hRM0UmV9i8is
RkPwGVQC3spKmm88Kz2QaKOsdCDrtBltDNW3VRwTuAlkTj+v9IXgXCrGEvrNqtJqFnWEzsiCQeQd
Uw7PaewDXthqu17l50YMqOMGSqk37cW1GcRGZqVwhrjNvUd0hPkp54LIpx66qJq9vijdd7MfrzWO
zCGIbwn9IJcxc4/qnF3Vyjuv5dg7GNE8qo7M/BOwLCRx47+atEVCEbCfE7YVb13ciZLCJWK++CoW
8LU6OYZeg8CRTBVTNBVyGAbqj5i2CT3hrNytZa6Kp2Uuk7MKhj8lGNIaj0JeoG9+/YecTsXx+wJK
JhiriwRWvv6suzhveIb7/ehUUHgVDPx8o+N3oX12xdUVBsK8C+5YVL0tiywfyntxxgjp3xvFMmrh
wsuXSKgu1JH9ROJ/paGfCysxinHGUb8tYRF4vgoBTGuv1SeKsseYeQrF1D1nhci5TgVDPHtbMrbT
Z65cjDxMUpuJ1FKew7s09QTpwL23VOvkZqGdZoqiWpEmvIBBHyteDaieJoFt/vDl8y7S1pLi4vfA
NSciX0ziI1EP5wHUKKLT/bTfRtptTN3q4IMX+BRp9YIGwhMregwn6o8YM2CxpIBuclJS9hIee4q/
4/yroGCVvciNKBhKa/IKCULZv/L5qvXHOE54f81uovwfSbA+HxmhjNpTZs3p6ow5NDCYcp9QgBgh
14Nnlbtn9R9gjOmo7ooZ56hkW/6SAYHhJC2dtVZ0SH9yWvPcWx7y5LUFL0a7/f5cHTM4HiUQjm1L
7F8CvDzkFiDLEsIqf4B5K/kAt6wPZSQMaN7Fd/JwUf7raQfHKWqnPp6FWydw6pFqyS74Hi1c15XK
LaDIiroG4DQzjHN+VYj+jozG9e0fEnSLrzcmvjgEzD9FeNGdoIpEDOpjmkZpbOj6L0r3IXGtbdKw
TLR/e21fyIJQjHm57Db7TelmM3xdYjVdYHIlLBgkoynV+rIfRHfMIaBTfNOowuFGM3rnax7/ri8j
Fe+547xSmd+iEtLxhbezcZZZc5NU+QJk+BAbo5xLJz0ozcA4FlHMrS4Tu+9Aqy2v7bdMXOvZLjS8
6v0J04t9FNmHsqFMBCNp0rKJgY3Ng52YSG/v0Fmm+EemJmKzpeP0vcyD0tQDwQr62DpuRRF3yf4N
4heC/uMsX5AxFgs8LHrM7OVWxbpLMuAhQigd4pdWzO7aizu1rRf8nAgPnRXGwW4niO2WV2tpDKZZ
x4BwmDKH5nounhrUuEI0x17H4uQH0UPtr6WTb4/ZvWiWXtzxvWfH1d3m8Qwdb2rDP5n2YkXHbTt/
IKX07q0W16ub03jtTANJZHevE3KObHOrPfSz+b5GyOJiHnhOO//UjqulasPemjcHQzJfinAkumOx
ohh0EwwYVpUO0zDD+8Q6M5Txwb3z+O2Azf1Y7Sf3VCIPKxDhK2PieQi9axw/1opgA3c2sMuVxyv/
hfuSov8Il4KsCIgLaRtUL1uiGz4QIrFLZ0M2HNBXI4iz1AUa1NIaLpHiPzGAFzwtIRgXYU0SRG8y
m05ucGBVUonQjTs6aEqK9cOlZmTwhtlYO/GcFc63pWMNKkXdFDILPge3vGy9Wb5uJXll7rNeybTf
/Hle7UNEZeOe88s5dQypjH/5qEVYMG53+sWJdiwLnxJ7NJpGSmfOIDczulEIG8qPYP+RIpj1AmyP
cxU1KL7wTCzWOF9yJpkeOB1+YdwfVNRmB1edofZHF7YVeHv0t9XoXDCg++WPWT7A51DZpogiJd29
yjkSrsC9a4lNNTJzLhKkF8wE4yUo3pDNklLKzhfUwgcEENgx1z9czxMbFS2Xe289U3Pn8qQzz+X8
9XMqounEeTqMSTrz1UI880NtrVmk7XXSJ6xAJ1yyG5LXqf+7R7/XG4AJZJfeW0t6Bq+X/cXx7iJ0
/NsReG9zVM7OwbjC7OPni+4nqnYA1b0bNeXmisRKRzMcoKQrnlkxImm0FsnnicnQki8TaC/QxnOT
Lh010Wj22f0X2A08+R7bz6n13LCPXC/+RoUYas1Vx10t8Z3cy6noE4PO7XOOdcMB+rwxa4RopSzO
2qcf/lDPHd8HIJXIGc1UzF5Y2nKrX36+bI1JpnGBNOtUYKn05RB6t+WuT1A1HafQNE5qiQxG4pU3
8hcouVX7tjFEYamxScxKgp2jmXoh24Mn9om5wZVLF48OFpC880J9hv1m1V6IO7EBJgnG6XpxR2mA
T3Ve4gjdh0QFU1fY+V8fWxCrmy9uNghy7rHfDLM1+H91E+AbNJSiecMYKulzt4VmXCAAUHHqecZk
0wiD5OirnftUsWs3M5WfDazE5lXBvfikvdNpcDrOO1CePUTEC4gusbWeRqTvequxclpyPfOreDdT
yG4xtW+mnO22JfS6CIlRwXBOIw1POlT1d6BtTi2R4zcAmSmzA+fDcYADTIOBJIw2ut/JtcROoSXj
FH0CZx2kh0EYBsdKzcsmOgzBVC11/I1UPBC+h+dIlIxG7+7YrcPeUwwAfmpKHTIp0TGEnBCfH9EX
NoRvV5Ezcw+bSny8ASETLgiFRTib2NIUNpvr9QVD9sPRxUGtOzHt6fgy0/gwgwZlnL/muFoU1cG+
IujrK/bNbMDVW0wwr/zrJN6hasR30x0cQjqR95O5XzL+0K9udl/TCy7oKc/mNJk9su4TAgOtWIDQ
LditxapoXuX/6rgKiY05XD1qounKXhmL3FuHtVblKF1bYW1AXj35i89zs+7x8RTVuSgaeF/J/7pL
Zv49fJkilRRKEwE3XRFrGnvWq+x3HoLNtPgOqCkimgwh8CUoBiV9yhjhW/Z3MTXBIH5OmrlGTEc/
dnj5+NQxCf6VNuxzTmz5lKkZoBtSEf+qJrya9kjfE51f930ZGp6f3e2RCep0tgUDyFGnt4K+JSM7
1HN7V01kD3dbB3IsGlb/Cg+eRzcSXxl4qUrFxhwhyl6SeRaC0oh6DaOeyehHrBRZjv49N71MycXY
9hwadM6vsnAOVXykSHxWdZ071VghJd0DWG0FCyvMexeODuAn4IYRVLgtXvKFUTz09Az6M8c2HYeV
WQyJLoPgx5t9qFq3SCKfj42k3MITZgmtftxhwWUXM4o391iG+NmOqrue91uh4kJnJflxl+IjE6M1
1+tT1izWY+MoZbJP6kpClsj2+OfJZD+svlBS6fqlPyw/z/zUW7oGphDt31YSGhRDKJaj414qmk/k
09TiXfzHxdHkWzYcvDO1Q9YGl2qrak55gxhm50XJ8PDPQ4KBZfZAE0SKMFc2VgYnAmPOopcJLVgQ
nRcI1NMoeaRj0/CYpU9PX7pihaLCMveQbzfX13zQ5wQ+MHfw9bx6KFeH+OWGLJQMjculcqvZ69nu
ifDNy3fxuKX4Dhn4lqDu9Y3AHcuUuaEYdWzCFALB2F0a+YExm/c2mF4Ds+Rm8rbZE8wPJTiPf2od
ycL0D908hqMYL5liyqXtuIUcx7giTwFPv+RPjuz62k4jBD5vbV0Z8DnqYJLo79TldfbMhx6+YvTY
tF/Gzu1NYKnZHNNTFtmwAaAec9hGGdibHQCMaZd39qFkqwpGR1Q7rdZqXgCzxrmOr//t5O3g+ti4
agFjW5cKivo6WhFQTXW39IAKS++bWEPDg0ApJlkAQTTB0R397phtY8ePydNCckhkTCCDya1oXWB5
4xG1C8uKPyZtxNsfu4+XW31cxnkR10lBH4l6jkWE8VkTY92g0TauthpsPGc4TeHcPLntAsLcEErt
gZMMrI7LiXqDLMpLFn6m0N+eRJDZchuzeT7rGb4DkJ94KoNyXkD5mMymZZnzbcho2gIW3K/2a8N0
NwOPzN70pvjbdU+3KOUL+rBlwHmoQiJYjeH0zz7qypn55ljguhwX0cOTKiSE59OukIf5b/rr/DUl
EfSq/TmBQqzEs2vc7Pwdlhs3UFD2LWt64L4FIbuLkinHusL5czHjgkLUueUeuTDWX7aSKpBs3JvV
VoSDp8Ym20jI2/BEAw+nkXNhKicjL/4gC8FuJamtcsIkJ1NLJ2NjiF3O+ECKKSfOWRoxmghnxLjo
Bpa47KQTFIPlQ+JGGPnQ7feSBiytctV83OEOG8HOZmAYgoH5FwutDSBhY7ZsIQV1gJUvrBKbO87K
btCi6s4hPTXHreqcqDh7urhIjkjzWDvrR24hm27rDHa2uBL6wA2G3R98CBwOAw93n0LEmxaWglSV
C6rggwKPJcHzixtdsEi3gW5TdPfFvMdnr5aMZULGCp1zPibKWWczRYGYREXgVz4Fz+eDuICRkeFs
GXrXsjnJVV4OV762Kj+afegWklRy7ox+wda3nlGkrftPTsXr6060BrNwl31eZqXxKkQc3euoqW4Q
cLvcokhuqNojk30dJgwRQskZRPa05nhxcAuXfHisAu/FqbB+xh7SmV5r5H8h/GhHn1YOE47g+fed
UJGTeZyrjWJka8UrZvZ6gSOMwyxW1147CBheY3qgNumHq69LMsTZdxUGfSA3KG0mFmFBH+fL+cy8
PeN+B3JqvYWntm6RJxpke9GTdpTmVOOZIP9XPLQOc/JjfLWIdsz0NrEt6GF2a2HC0kpJEmD8WTUz
F5fx5b8wFbBth7++6wyFx9AWBan6SMx/mF343up8JGDU+fJxwe89Nsj58frHtlX8oZ9ozfTJvrYU
32onfwjEc1Y9NemFkj+L83t708oXva1MNOKRzsvAVZS6LcW7cRH7tN8qwJ3hYKkjQfMkDbdGtjpw
PtNE8zqsnhuPaBngiquSo0Zpz8dj3kAG9WPA0P6Cgh1UBaeupI6HHDTjyHxdv29cZePVTyM9guKr
nWIOtc71svhW/LHd9BqOu4PF69vESfizhkiCpQqmoTooaT26dlhNKPFmW/gzKu78zpywTSnLEy6I
Hkr9ZfC/ub/FqB5FwHqBte0Mymn+LmlWt6NvUw9eDn3getuEnNumgNu6FhDnrC3xmjiHli8MWfM9
iLuL+3QDld6GcRTz1iwqcKHnjbh4vsUznypn6lyxcn61upJhZLRbeLvZNbrL0ptZPm3YBhmqcdLR
r31OFoPXyOnZWegWNO87KK9IADnkFbiAFPsTCcnDkYy/8ELa9LEv492/43vj2Ofe9jmpOkh0zbbT
iRWwrd6DmZmPhZlyHXW79YBYiNGlJUsaVBA8B14hrLLdKyVh3o1pCI7V4obonCi6l98sOOfaqrjf
uxlmePw0ow1vYfnKzBuBn4SfroBZSqEMRbbOf3t/ioLQvHuPMDKkNn4CZQ3cgvfVcGNiXdLU18Ri
d6LDLakcxDcMp/wje1Q+1cp0Y0Ngy6WTEu44B101mzaaON1HS+9xp09dOmJGO22dwqC5T4su7+0X
LfhBy+DuehnzNSnLbJ5HUFHkvPWQ4a7Xx9zfS4zXogJd+ygLF4qJm7l6wlwEr41SafDhlWl0dvZo
c46hwVograDoo+0HxAU4DEHLJMqdHOhYrykPT0SIJwE9U6I/7DaiCPbeN2VmosG88Ghn4TL+QMMx
akLvlzEFAnmyiMqwBe0zzSqwrzYEM6InjTpIDqV+l/dIA6/Y45ch28cWRIUm/9TnCASRSBxIJYc8
qcYtzl49/qzdqKMJq2YfWAELb3FlQV070v2EJB4L9v3dswlSJtzMxDGEByrWKM2nhoJP96k8dzOg
slztCWrlu5KSETpvlzEKKU0ut6F5W9CZ+MMSix2dUF6BJ0rSOi1LP/3i33TBX6Njsonxe1W6dgQX
ujRVBYVvPpMAvt+6IceOmj/bXJovCUcBPtS+VszM/1fUwpEDN4oCL8JIS+xsjNuzp1khjImQShbN
DxBvwIArD/+wiGBii3XaJ6ixAWvvdypU+4teWGX9v+f0T01ZUewOrm/+IcQClhTwpGifqO6Q+E+Y
AiSet7PlQG0+vTYilk/heWvNXuUi993aJA/ieoIfuZvMVcAqSSXS8J674YJtu0IQjb6junlg/H1B
XY8JDhey651Eem2EyO/yFDUBFa3HcXVXLanPrP7Q05+6DbdQ5XPLbwuqvsoVbUbkWkwLfo3Kt9Ut
sUyULvi4MaaXu4oQgLDaesWxLExoFhDKbmp88WWZqFzsmJWUT21UwoKfQwcqRpITLBMbr41V3poy
C6nmintZ/pM0KKn8nBJsKmo4MlfRFJqR0MaBz+8Z7Dd2NnngZNxCo1WvEq5m8gjH4eCH/70sG7gB
4GEDVMhJWHaOqwLy8+vhexCkbaeh1SuaoFkrtDq91avaUiK9JV+9oWlHFzxKFc1DAQbWsErZeIYh
NL+HcjsRyMi51iTuRad1YWHCsQbuBTpdEl4JdvQVbHwTbsc0x6ZGNFAtDy1g5Y3qPXFmGMM0FVh0
ZUaO/Roqy/ZfH+erH9A3X1f0DQXnCLUfelrN3peMlQyrOobyfJwOtEbDp2SohG8Em83gnS/a2DZY
dqRSjHlnfCSBAMOP9VjZrLaIE8rwd3oju/hvtp4Bu5XrqSTQJijRtsDIfhVdB4yUo18tDFiaQtEg
gorKpkSH7+BWAyZ2XDJtne3HGH1MCVyuVL4pNynhmZOYh4z8RcnglOQEYpusJIHXZYNQwvqIL7r7
nrI/YwPB8DsBiAwNBeu8B2SD4DyMXNaIfww/rEwJHrv++i5m1+0cCviPkXekAlF5JAlfS8Dqlfs6
2i1CTRTJjrzEq6unzR4QXH3SYQg/9KCE3jSowauTm8FazGLLprsvMYCLpzCzg+1+p9Locjg1ISpu
HZCYtSoOIKbxNM7sC5IOFSPOWiXTHJSvovjbmXSrtHZIIpisWwX5ofr812ZDZXIFLalSg8xyw90z
kugg00pFn/KSa05Uk5TX+Wvbb3jVbu1l49BJvj1p1WKE1hZCT0FmuOkZQsu3MUN7SV2lPiBEMo2A
k8lfbrLqA65M5KN6YLDOPGAWcZjjC8tFXCntZqCPJHv0RrfQLOqq/gw1VS1EiiE1WSDZQ7rlGkVb
QXCdicbqZtfF+J4fejxiQzxqobskoGywN/1/Tw0aDsymJBx1goFzbq24gAiY2LqbzrLe/J12JMtt
hTkb6BiJgkrtu9h0A4SEBlr78wk6KeE/yiwZVZPDNZ/qVCZPlkfb5kPtI6kUtrBZEe3EuVnDbrJa
JmKanbYYLJ8iuwDAKv0WUMJYEbzUaNEQZwwS2j7DBEjipcx5qL4N3tfWFS7awccgxqKsd8bPg8NW
p0OfEB+mBc+caXF3bDU0TJEvYseC9lJFnnrsQ40dDyKOg1kR+nHYsti0zVUnuh5mkrpDkgnlQcuu
neEpg+IIMSFiW8F/8Ui+vJ84rCE2mZ9xQGI1pFQ6eabIvNU/vfvkC/ZC5gtJn3jEIYpCdEzlt3UT
RQl0IUFCV6ZQydPZnoiL1JUCyApo40qLCAktYXVGz0XMhMfixZi94IFGPGWL0heH7rMDvDkgy/EL
iblLTSi+MRYSHZMYHPxF2GiA6tEuJi9o2YJmGPQlXYbWPbfIGO7N1NcDnd3O3pZaB/OhLV6WMs6x
qyd+XJzqxDiOEpb8k/QzWz4tKtP8xF/b7t/RxF/aSm4BjMaDTEm53WLqpMlVK53zOWm8odyryXBe
27U4iUdayt2Hkbaol5uE3h1O+OSgU/JPASqwHRiCqQYRfhKuHLVUREi9s4lizsRKGtjJd4Il7+Ki
p1kWjQ+ANl6r8aWoKSTELbqChZ+gjBq4aaRTqNsRlclVTHgiJJh7j68qz/mZV1TIE6iqyujyrrp9
QdnyxDYUWCEyOpaiLUC/ybMdML7ZSzhe8FHe2FY01N5Bo2vlZbfh/lwt7M6L+L2Z6OkK7dhnTKIB
ErWRYZgs0fJfOIvM6am0QzYNhW6JaQZKRkPCJ+9mRBRFrYPE13DBYv36WLOr02ijhARXnouULbWs
ROdON+S2rIHT5aDeIYkr0qv9zo8fmfrfXLPMp0Z6AyWkUG9K370hbxdqDX6HWzQRxWFAp0trjlov
P/OCcw1Vrw1MfWfcga/9WZu5p9YJwuJ5zQc4jUQI3Cp7hf7YeOG+xaqpur9QU4LU+T23B9CpLw2G
0eaZ1nrAwHm8Nv7Pnyr6aITUV4u7G2eoiCy1iQhKJLgn2jyrqMHVZZ3A7Lf5dLevaLTlkPBdfa6Q
zkj/b3K1Hyte5Bl3kxKsFD0mz0IQ2DLLxiiuiopsirEeVth4POPdfk37uzKFx9QUpOar4e0uM+rh
FD4Zuif+MzSIewXUZDYBsZgTQIcvsdLrHXlNVUDCGtSZ+F4G4U8kOslv0puPG1BBkrRSshS0vx8O
PACfclvMC64Y3KK5pCQzybKjYVSbSVYfMz+dtfPxE990EOwxgSGn7LBiixM8KD8wPfdJVE6CiUqZ
kOu1DsnAn9epkPSaxsevs8knoVkplzSVfmkIVFjYV91MXXG2knZZexZtzoe/0hmMxwleKUIlO4hf
cwdDVKJ4KPVBDqATdme3kGJfMFKz3Otj1tCPWJ15fPsI5qCHhEWeYteKsx46wIVZRJtLwWuLNSQo
/xszksu3vURLtW26CxzWb6YX4OvdJ7UnjPEPocg7Ci9OToVHwCN4zOLP3e8yTxaR8BarPWMe9V6Z
HdOlkk3NPNGDabbHdQGamKE9ya+zUYHcrWR4/B0XaIfkxudRsV4ybBugkR7KopyRV1YFLTkB6x+L
xQSa4haduguK78PcKPKkbQt61lZc3uZw4nyAqLTkeCNLnViHu0kucitF30gO+WJbU5a4Hab0LmOB
O93ruZdt1RDF0IqKEA1t8ekJHWMUGYTyYslK49zCKrXbLe3nPb9iooWt005ILRc71c+2u8TyfiK+
GTYLFnpoIOJHsv8vtXpDuTa5qVX50aBqub29Ri3qQGxLSHN3HA2sYJBQTQb58zetiUu7QZJRkxGZ
vclDPgi27J7cCnWV8ac3AacNsavZtAn2uMX9+zdr5RSWjn8bWT2A941gy4m4iZc0pQiDBKKwv/jG
yTqiLok5WSDgwuxtjxbDlpKE7ySoKs5BYGCmHL4yXhvKpPPu5+5TB+MzIpGFNnMsKg8MQj40SNXs
tW5AUYBqCppGLuWW2kHU3coKry3hvG5zPFFE+83ruq71RmXoTPhE6QHbvn8FwxQTYIC5UPDI7PTK
yZGSqmcEHfed/dAg5v/xbQ1h0U2q59KU7Mn7jJKJBwn3Dtls9HDeM7Sy5cJWt4YjRf+/FKcO1VNR
n63uTLg3znnaGPc6T6YlpxYSi2CCleqf4YnWwvo6h8IdlZpeCwheobiumXhYUetshBFC2hzQRPiY
YWzMvOUya9ZPSSzZtW7XehtxD8r0IYz72UkE/rxBwrNuY17f9fbiuRDMTpc3j+yLiaci2xqWl3aJ
KObysqLLQd4QvCFFuNw2N86hqcWdBkdwjVJB4mFWltU+U9W2Dur/CtXEFVQ03nUL/DWI/kUeBO8R
mJkth1H5ePgDI0hG4pP4e8pzfYh620g40vG40AameZQrvHVUI179OBYHpNBojtQtbkfMoYbca7LV
aOF0Ps7fVkGhd9gfESjOCrfcN86qhlkO7a30oIapY1uLVqocHhw0MmhmJmut18gq1DuPkWKx9gPx
7WE/oceG/Z/wCw9U34dIcFQAFduZMGPu9VO4ZjJvkEbqAuwvFRQqYkGmHf4HxPtQQ0IraNUjMghp
HLQ/uDkFnCaOciBtUKYTZmdb0S7SiupzESC98J/1soJQsarmokhnc1SS04c7NeXDbq+jMmSXDJJv
hZh7hlhe0MFVyJCoz3Hqkj7KH5/1QaqyfD6nYBvNh9bnwNlzhIlO2LdXqInVJx8C+LNkNJuUNQlQ
eUsuR0zJIBgzJ52e1KUumRAQnVlOGuWrgc7C8oPxvoPrtpT3UaPn07ii+1mMfJTccZ8A+9wS+z4O
1bh1RzqhsACll3XR9Ojq8VciSVxiXEmLKDELNkbYSPG1KqZ03yjhBBq4PGN7k0xfssflF+Zbfy8+
HBipUTlj6IOpjsttMNroOBf3o29xBNuJPOvtGwE3g3zRT0LURuC6iMT35N6P92BFWTcILeDFx7QJ
dhbW03ThAvs9crSOrTdOPY8p4A42U9CjnA6EyeIxCbNgnLy8U4cGMWbk87HigQcxzaLsF90Nxhlm
yCZ13wglvKwwMkOJnN4yW7ktrt3pBEsdllj8cUSYcVP/LXxAnwLsM8wlgF/AfhKczsyD6AQlWuN7
Cdo2DOlQCXv8y2R4uyGH0Nplbx9jHzeaOmUpUHL7dV0c1rkPi9sCjDMUw8z+AA3FrtaD9/8sGKdi
9f9Lkf3vOZjGTeGp3wPPNh3YA5pt1UF5opkuoxeW7KqXhTzYd9gxSRhhuFo44T7NlJ2t7T1tbzYC
y9zB0Zh5xqUoDDT9B5ZNa1h4f5sENVbXfaIqArOSbhpS5WszoeiSRz1/HGRRqrI1a6UogKcw4Gtv
NjeTuzxHky51i3kWZ4vqJeol2MwUyTW/eTl+e12c6eABhdhhmG/JCM91hxYeP4KCpthvh7EpLvRD
Bd0AyYyrXWyp7F7oauvfOCgv29y9O4Fuqkyc/Xt1DE/063TXv2S72OzOJUmerH+kAdkzQw7B/gRb
RFlKTHYGpfVloWBbV2aH39QBVp83QToFpACfiOb5RcT94WYXh2Lx77TRJtd1P3TYcWeUIOq5uynz
G6iHc16Zf2iZyHZYkK6mEuU1XQ8HaRu7SzG9w9y1AiQwA+O9+zxeBjyPnYq6M4tvBv8WHzC8BnZY
XBHkluiAHuasIvN4CcmMPhddwkxJ00uSxrPkBAjyboBYdbntsLF6BANS0jz5V6xZLCNRozLTOJ8v
iCwR2vZ6JVal/PRYwfLz56PhQp/MtO3TLvBmBeFk6fKK7AVxo0Fvzt5tIA5MLLdknoHj8Ueyfgmo
WQ155BzDdMgLnlEv1vDLEdZr3e/fp+E+AH3OAcXnJM9J9yV95rgBjoqPy6Qt1QbvfKPyTlypIC9A
V3JQVuRnbwQ6eZudOkKv0cfhMyyG46YDPGbnhkAbKsx+pabEzBNxBYnop3T68MrBygjQbRzUJKDO
Qms8LXI2SVeSbo6fF/XGt63ZZotvzHdJZCRuZ/bozEhZet7xDr8npXtME6F8XG9PhHnmjmuCD/UG
FmhRJQZQKv3stS3KXVp9H/RgXTIP8+/0T62Xaj+ygIUgk1rWFecfgQT7ZaMBPRg65m8JzRRSOQKb
bXSlVbW5Q96ckj5TD+ArwYdiS+KjwAye+klXY4FhDKeb1Aq/v8dM9Jzc1LEz9t+rN9bwlQX8qMLf
F9dfTTqaqmgcNfsGwTRTeEpkw8PMQzQDoSTGQEz6n9UGNCoSvbsOMUDABO3wlylggXRcgOQ6AMrQ
xoWtNyypKweZbf1wvNDMvNwmyGJoddxVjHXWiPJ0kbKuIno1F2vxRHNycw0IgCD6nMFQT4P2UdOE
1hEHlu8sHj8VuLKD+UpsVmNhKw7esrYomcXTyeM5QQru0Mm2rzxnEmwQ1ywQ3RK84XiJDgTke5im
ThfK9NnNUJ/iZQtVIfkkVL3S8aVWFXVxxvrfbEtCaM3n2lF89OKkBx7Tga6Kfs8IQt7rkbYwB4gb
vaZu9ybkOkwxTqod/lLdJo2+7r7NgNjHlHtgxqUvx1h2qgNdMpBLFLWbpWhtB2GxqyNOqNZs9Kfr
lRe4tmrU9r6aSW8LwrTQIAdL+7NnqMfM+NhP40i2oFW9xH3E1MfOqqYlW2FSXY3kcgw5LDIRbdI2
9d7IOjsr0sUNamcnOMqvzQ5hnmd+np755AKFGVHZqD2ZER7JSn0+2WZszF9a5xdfyfGAGnejr+1H
jvYOXCApZ/d/Uc/JoPq4uXuWSDQE1MoahnRKqqdVRn8tbA28VotnbLA10AolY61LjptKuTTeuACr
cqhrtI5YEJvq+BudC5IDdg5ZcGLFmL42pCiSRobT0sf4gcOdqw0luDIZOBVjbrLDeKpROYKHtz02
UVjZ9S2zHmZfAeo+vrf1ABA8m9k9avEh+c9NEJxHaITapdBpXFh+iaLyYIuSa4yyWuho8Hit7Seg
KJ88k55xKOsmV3w4Xk55XCsljwBupFybFjAhrLBtoF3ALp5fKqtUAQGgdYZzDYZ+TRhek9w9rGe4
YbMsBVv5EsEkDOiPyybUgrNiMittuaJi4RAMEbLkB1X+ooicrFfJqRIaskVqXkjniBTyJBYPN4B2
aGULXdtOjSxiL51lC/8PdaYT4cqV8OIba/oGgzH16nfUsPMF0VXrgz6PEdDYIAubB8Na9HJA+Tkw
f6gnrZxyPiCfNMauS/L5G7O8vksOVysH3WvDRWARzGgBzJppeLdZyTHGLrruD01xkg7UgSzo5IOQ
7hxv+G7OR+jp6wgOhBg5S/17mxyg/G8F6se6lsZwP3+lfbsc91ghQn2XvE0bDTmlWY9shpFHaiCJ
5Cku61C7Y8IKmBx6axMSV90L0V1jtrMno6ROguUq4yH6GNCEyQNfmFoNcrgX3eTYM2sTd97ZlhTk
izQSSLnCAayBzBc5lg8o2YILooAMhxMUc9YIiW5Vf5P5+FVU7EZgTnsjhQPaqTAmYgoynuSZoFSZ
TdoBvglE2vASqrzOiWIGW/9ihLLa7jBdHisJhqk31XRcwZ3Nu4Q1BlMjBSm3r6FfeoBCl5iw671q
jyo733TTSaGF7kqhs4dAmwk1kpiTGH0ydsS8j9arLSFg4a73uOoq6zlkZC6vP8/Lp2vdzdt/GwyE
A+gyxzYN/HEtmyLjmxK6Shmx1kldn1kcTXrreVmXA1h8Y9wJnggXgrextxaSq6EM7uV/hKgDPVcP
PCkOXIcRd4BWUMnLx+l/gS/drmKk0gHQEV1Cv9BZ2uDT1Nmfs7PvaeVtE5uz2DEbc5p2Ae2YJdZb
gIwxksbJkhW/TTq4pVj2Kb6EFs3uzlCnRLIQruh5xpLlrCtwY0qRsZqj/RjuNjhXAMmJnflTddUF
qKF5Arn0+aDUdpwiPOzca42iNIitiWnNdODNluFdqj+BkYz6lZVLLiM8Qjh/s3fby/WIlNiiGb+E
J8WtUGMxeWCgeiPwshoPkNNwPRSFKTB6atFN8F+yC+KFkVze0MF+EdONSlhGZdjavZaK0EMe1QtM
ZWCl37Eyy9/5c7jjm9PFkiBlQiDufFl8mdsmGzqkCB9OEGTahgibvhqiTr23G6Z+o0iZOKFUTuzJ
iklIfTd7Gu4WLQkRXgG3mhNfAOi5KYcs/M/4b3GSwvHyAVISGqelURD7IHWa43OHVtIg0NBT2jQz
jQwChrzZE+FxlbGzAZCme/FGWghGfr8x25mDoVOzB0Hn+k5NcueYQ2vkzRL83XocOy7ZH7B1BcWJ
pQVM5dKtYUhJJhs83EgWI6lCzuv7jb9EOmaTfMaL22QjNVjO1uGgwXBk5DYK2BXvbRG1DluQ/3B+
aoZ6j3w9vn00RDfbWL6iu/ypyS0DvRvETMCG6K6fWu3A6NDcY1yhB7aH96ZrlQ7TZmeUdDBeANvM
xjL0IXwpJHWv0kiiBQK3m3WeQ8U8FUOIl+LHpeWvrGH42RTzhaxEzNVBJoYZt0mFgCNG9GnVGDAY
Bip36NNUQfhj/qyrOOZx94vTGXn2A1RmQICHpYhUjvz61LESr7UjQWddjkg5MkJIAMJb+Bm4m1iw
mIh7eiQVgrRufHlO2/IxB844pC1C6Qs6eQa0/G7l+j8mqId1k+dckwfCN+FKTUz27IMcDWpszGWl
++J4curUFthLzMUzJEnTt+pbwLvRZY03SlAlmW1cyIiF9J0MV1tWLtwvoL+xdqXa4V4Gu/BBvl8h
sAjF3MGkZzeLzG2LHDkIrrYr9a2nN7HjaZg0fQYG1MaGuw4/gfl/XLd+3hXodTUfH37+uhE8ex5J
CWw9w+DCF+tsQ4PlN0ivfLeRG0DmaAqANiRNTcPBojf046Fa/WkGq8qZYAHd67kQiabYPINWurlO
YEUUgjjJD9LKKyqbKp5pp3Xph2lnsK4ITBa7b4xFByI6QY7qBM0ryXzjzeNS18Ryc/UAWr/2H5Jn
M3+1Ul5yhaaAxuDZAwQilKpePfzSPlOGJY+mZENeDX0IMHubzqN7OB0vyAcjAm/BvIYirowAvkVS
tNpb/uJoQzYoyGNQEXMav4bxTBFlDLxUSU3nlWodgxiLbC9aspYnwiLWo7U0yE3ymYrZcjEUdRh0
QKs5f5yd4J19otpPFrgM4Q9StXdwyBPUkO/x+QBqd2vF8f+b1ThyF034sBLvRNzJXO6qU9HbfEjr
0uEUaf0+y5qXKfTfoF5nWtgdPQOfOJ+e9lGz5MllknhpqfLNbXA7ijsSA/UupyQCmqQf+2QjcvRy
j8TaLijGr3DwwN47oU9qLuEseiOFAoRMbJzlca9r+S9vsnUJuMFNAGkGUHz2ELdP9TfbESjPujjW
JjRCfkjmScLyanCEMhYyOGV6jmpAeXJShUZHyfpjylVI5u7OXK/KleMoroSUJOGEmj4TojUm1Dzh
XXw22g9fES5VbvcsdMyMbSQE2cK0l2FuIilglti7kOeqbTZiqOXBcQWopfh7UtRJbQahbH4U8stY
CT/aV8J3x9U9Fv0h4LcZPLQtIsbnzBh1NzhN9m4Z0gtUn4T3iidoxl0abKhHDZ36x2dPHE0b2w96
YD41H6Iwy2uP3n34QriYk3O/XRVHZvMzFzTpYfq+6DTZx0o6mee67Cwm3dfY6esdG6KAH7/HHaDK
T0R3s2GOhn+GHWlmurpgTtPxpaLckJAbTiwB/Win8LsglYX113FhBz96i4zwa/th/ohgY+3Ffw8f
sP/jcpcmnSEkpp8dTsfpE+zJXbNdlVlAfZcC7m6Q/ECzzRjTft/G7arPLJuhbykV2MgTZo7gVvUt
rCmBJbpgjSyiZ455fi/JRx0symcS7BVU939btP8SS9EBJghCpvw6L82apdHvpAOyxonwTPlWQLtE
9PzCKtVsdhm/8Q7xE5Inxp+Iky5Xyih2VjbnXqitSc1qAjT1eu+DQpKg3wJDW6CpKaAycjjT9IyE
WeVmJt56s0JbvsXoI86WVdvXlQQ7KLQlYHwOMLnS/iE3s0YxkxWCS+2WDLaqB09scegwQmzplSny
PYJDMFMsG7/7kZ1nNpv9Sukda3rBAd9Z7eixu3PaWDv1iH4DMebcAkg3zCzVVYAUH4fTOUaVOq66
NHsWOxssiQnqq44IXwARXozYzrWOxyVnRLlrWs1Af6MbLMXIA46YKnSB6YgENycOk2RjFKymwNZQ
gS6coBnaUpcL3+usD9/GfzLos82dTCtf3GkR/1vmV82WWKTi3GuzG+05hnqCt+p3Vz/JhHXoUZOx
owQoBkPU9dEcoXB91dFBqV+pCGaCHn+fDJLmvsKzg9or3wGPJETibsLs6dXe0VETVHf/lv5dOwx7
5rD9nKiHXdrIkQL/of7xoAlmvEBaf9Tr+YBmMLx+vat2EOrTiHAP1/XzeR1lCejowGu6sLBvQXEC
C0Z4XoV2jUgzm/wfo38FIkJA2fybMru7hEzdqJDBLsqOy0XQHnnb8g8yGBRFGEjNLWS0O2o9ELP6
8Ul1KngR4BiKPb6bo8RswLV0ymmfj4iXaKjfgX+UeAGjP59j6mkgZRC4GXB5ZDySjrs8TbEuTGcz
Dc5pKjRs7INXkhgJUa3QiTGguURSHLUxssAXLckfEQngcHTvyp/BmcGx6Gx/bIseJ8LgEKuJVANN
tKh5uflu/Mjzq7+L6XqlmN5LLi1fJpG5kQ4Do4HPumkshCl0RdCtZ5wTCIwG18MlBOT19uaN5SpW
ibNgOuK7l6ypGHLG+WXvFGtlW+LqSbH3queZZ7TCHa4NipwJoDCjTUOqD81IO7365fCLkWmwN3FE
hlnuD61lCqScbVwBfKuroNZU/gdipVkh+thK9/3HCPruzFvP+BlDOC6KhdG/dGPM1oeqsPUcHrNa
vSj4stNHDBCPUnzQ0em7xl7ItVbL8+inxa02Lia6zoBeXY9nDFaYcfZP/i/2pfuprHUKYK+OnsrO
q3LjJNSHDhStGQjbRmzB69Jz8V3p+Vb3BtCbENeLfoS8VJPK4MmSYHHnF3PVcVbZw1F8VQexA1ua
eWIcIv4KAQXOQjNwiNWHQND0WbikRk9PsJUZ54tt90/Kw0tcT36PCpNJyOIq2qmyB1e8R0Dt1UZ5
qAK7qDT4qzV1PAt8vtUiOQW8F/wfWXXenJenisVjfLOwDuznPGNwMy2t9reBFW4kJB2s/o0NT9KD
Jf9O4CEOr7+SOXVTtGixeie/VAyrooJ7BWO4HLmLgyjLf40KlRSDm+RyFw6UBz7ztqwMHWppVbXA
cnsMYCMYmBBK5k8QGMwRTtzf1q2DKy/3GQW0frhRBtfjSm4D0aU8JRBPPLzAW+oH60VlWY1hQ+47
4gMu//np/o2MrGXaKFF3FT51xC2LADElKeI9TN1P+8scC3ktNFFQPxDVkK+pNtwrCdpN3W1IB74E
gE+vDWnDQZyF9z2YnPB3ZskhzHobHYklBNxPrnfE9Rrw+pNKJumPf0IKprSTVszcvJwTZAlNpFZF
vfrbkooxb8aXWAvsljZap1L9S7x/8SXUs9hGL/GRsLh0iTz/bYUMQ0wnMBihONvdxGvYJv/gAxp7
/FW/QgH/J1gITg1vugGvjpl8Fxx6YBg0//GySjh9DcvYWis7/ugZjqsAADzWLFM0pZmq8T7pBgSC
qNpdMyKZej8INX6siPj2N40WZKOE7cjrxsFAh6aSCBO0IGhlGhrnzQCvsIXSpmTgOHlrLaKI9B15
PmAJUEwNxwPYAOfQYegHjn+zXlr95zMSe4Q1BeF6FeeDWxkdg3U+7s0343GKthCiLaEKR0B7OGF7
6iArEXMWE6U4xGEiQItLA4qTwbeknkGT1NEaSRy/Pr5BW8SXwyFRAGb5om0yp03+Js8yGXlW9OJ8
fZ/6PZh+9CXJsM2DJF+buXVRm0dUiMCqDl4ffi+g35YFqT15TNEt4YkrrENfzvZaEvYPJlPX+Dui
EIhVRGiZBQ4JTDOXinsu728F7MFB3jG3cl40R1xOlublkqQY8u54qWw8QDSY7gPPf86kd5g+3WvV
m/L/Pf73w/8VP5ggdgomgRr8TFJRX2MWKGVK56yFjkQVPAfyQJyljBnnI59Uva92D8PZd2msGTzd
a5cIOeBLRAVFR3CY5rxlGH9P2pJj2OBA69X5q+bih0D6+jBvFwPh0qfT1SuYD0eVUlXQoWAfC0tU
qsN7rxjyE6nsEaJbsy/F2pWYZTbbT/llDU/ZLeG+cWflotsoCch9rSZFMHoKERipAjYxfL0cHADX
UP26KilYeEgU0k8muQ3g7Ix8TPu5u+NgpG53GGy/Bb7Uqu2zmrrUAhJa0ZuWFO3/t0LeI1kJfXOV
V6X177EnJ5IOSNucPD5HorZU+RDmX048VBj/OAiYl8r3Mj0x6BsrfCXabBmkdmBz31tEb+lfCiGf
9R/5cV5i/s3marFR5cskShNQC5b/pxbsjKgvsmtIAhAzEDMnQrepMghAlwkL5uPt+L3jOpmaAA4A
cDY00mJz7dBpXz6lLUOYs6oGro2wNG5PQ97EfCICYgyvnIcNYMjXp71MDU0VivzFu7/CnaGO3DfA
ckAcSH1ANkYQfa/TgpjzKPH65kgSm9eQ2wPchSS+FVDn4WxKlSCFItxGz3Q4qhwJErfMNCocMyLi
WsRdPN1fdNsl+kVS0wBpKYb3Myb0aN8svsFF0plh3hMhLKZWqU0ESJMNaKFZlQZubdDn2Y9c0O5j
BO3U+h6NMf7Cw5yMVLMorfBbBLTejruYneqgmKdTDweaCHGWqGuPIHxh3ov90X9VK1jXtd4SZ8aS
MvJYysDq3a7v+/NyHUwnhdKg0vGgFJFcyi0MBGdd/g9ibD1TEs0vmS4nHofjJW8MCz+0muQ9TJoo
XZ1BtHeUxckDgoF+ko+PKoFA4xOpNq6yRy5Vn2CfaCam0cYSTmDqcLCRSb350GFJxcFxlMF5wW0V
+mNlfi8aArtWP2IcFnTZJRKN8ATqdPhNFp03h6akWl7F15rJkvCM9bQKfIsg5O6FfgWQjI9Uw3qD
ZZ8Rwbf9J7DAbajf0LUtJF9CVoilt4iuJ/5QMKj7cm/1bDqvujdBrfQfr9uvUg1dfeE59RNgbICs
f0myeFh5LDL06p0FknrMJDDpis9Y4T3TpgWy5J8kyyLuuk3Lh+25YK4pO9/Buj0N7K27/4IeYHsi
041OEay0iroe8+wVxiVPz0aNIc8lnUS+UTpdjM0z3gCZZNi8z3Za05+IOtHFZMd+huRnmNNNk5ya
20lhenlE5RbgvAH6eb+KMnG7kUC5JvmZyDQ8uUFYxj8Kj0I/3BTbNRlQ6zwBQa+P/KDTwFN6gDAz
2Dli1HssGwFHJUSUnC/BG3fpRFv8A6YINmxEzKIIKhmHQ9TP/savglV2wtza1SNgX+CynzYjc7uM
QMGSfEn91fA7lFsZpn4cDtya7DBgPaAkTt4mKviFq/E44pdk0rsL8IqHuBeD3qSS6356737yDAy8
BjezwsY1JZCAuQ4joM0FXC/4MmvixL6Aiz+HDRWEeFyIbLJXd3ojha9zs5by+i7kf7mQo9mScBmn
2fyaIp2NaIvGRuT3ltyPhFjpmyFH4PqYz9m1iQiRdjm7WwtNZgovKk+R1I1BIzOfqbCku0oIg31F
rspwjw0lnRVHyuU+qmTvDFWdHGuCoDk9PhGobWhCTWW7PAZN0+FCveXALk6Hf5lwHZ3RPL0+ghMg
r+F8pFZ9GF3NURSTCm3i0ZVCyaVVQbcy0q9igmnCZk3YfOOT0vcC5zs6ufhHP8UfYCqqN9ZRjpDZ
5KMFuZKUXGAJwBv3Y7VXbJezbiVzDTbFjUSx3rUWPg1izVlWrJOx0vLdF1TweBSNK5MuWRolpmH4
C6x0y9ZtCy84ke8L0VzpicFV+i7cm82E1fmQym5EVN91yMXOPk2gGK8edbagxJQSMVCEpkAr15C4
NOvWDK4Hh7+vmb/9pLeRxl2BiBIQ+0GJWzrTrjhXbOseXpq3MaWc8GKSoe2DJv0+skLJl9KByYsB
h3R0vxAz+OiGBCd3CAfJZheKIoNuJ5/q9Gw9I+NXLcH+gWV5t4zjiC1BqU/r5eGTW4wRnR9j5zuw
ud0ZtUn4oMkztlB+0H/yILP4nuT0aX2SnfRyqUy1Q+Z0CWf1n6xX8PvVcguFpsPfbKXWGG3kusNe
ODCwEWW+imJWyyDwGkVPtKmxLi1V1Ls7hAyg2nGB+hEuFw5lJI+PPgs91XHNH42JuXuQ6AC4ENM+
RuUNu8TZ3+xTjPFcKYGjBm9koNEwr5VlhFTxAfU7GKR/CHYMIDIF07OcV0IhOnzb9UdX52Upn2A/
+FaxY9QTVZmtRHbnrBuWKMIRgnhA498HCe/AH+Gp2i2DAKS/k04sxaGPT0ncbSEQUrc/kz6xVkaB
ZWhefYPAxX5fCnThOD5C2XskQAt8ckttiU2UGK3Ishos7NActXuCZSlM/K2SyYfQmQXUE6IqTw9u
wEvbl2ygJIH6FOBQ0pxiohXr/J8DgKuKX16/wFa3bNgX8Wg2juxEaZKK7gvs0rqP6eWA3Q4LZseS
vL6SdSgTNIyDEFAiCPraVqCrX9XWbg2xfaBm2lDGj2hYyigoPLc350DnRxqW9mISzA7b0fiRDugh
YnKxxqa9w3HC20mz72lgcn20wTFyxmM7SCZmiTt2N9IpcUIjWVOtT76J56m4DT6GhHbwAu+4ZdLb
HckbnnLvpSAcuVauHBzRM+exlglsTRXa99ltRkLBwW2FmMdZVIZhK2MccCSWFe2C8sKg+HKn2PQp
pP2FR2uahzu0qvK2zgznLnV2TnIIsMGh4wxfJSN5n8oRPFr0D57jIo/vbo2ZABTo1JwUHGRWaByN
vHnmC6ZJWphD7p09UOENX9mhiMpXwSX1gSyr6RYb7Mlu6qVriXOZsGnqWOtAaPcbrLP+VSzki2AR
ZzgnPHkILX0wJYz3TRmYEi56/C+3Oy9AmwLXYvlCEG5zq0fPHPwn05pUm/y6Ew6J8mnx9FTvNnmb
RvzrrN4k5KZo3MDf6ozHkR+QcYgPiOnowsmc6lZ9GCRPwccucD85UCPJPbBlIPsKg/k4ZcedtLiy
w6TQSr3fDAn36BE0xWD5RG4ZvwTxw2Dcl0vGjNo22lda/00LO2UJ1TjsjAXlkLDEa9iOiXSg26ij
qvAd87kHg6O2Q+HKrYpz5Ihdp7xpBw94d0Q8SZhUuV8ZhZ5Z2syGecGMAXecfGGFmerOE6HoOcIf
tFr7gb3f0AD9E6z7mcsf6eLMLfBh0XDAnHqduOoE4UBxd8yCrPXx+KsBIDBcbSnikD20C30ETre0
7CctqlhIEAnQeXI8Iws+uGNfY2l8FB5HbUd3vaCRDsiLEALokfxDpTaowMDHoAOrWGxAl/9hyQTG
7IuxNqHaQl2iJ5LHz/lHfMzrBP8Tg3XDpdJKsf7rDDnaFTv6ak6UNHkoO609Jz/XJSuCQ9LeA4iL
rhRRUmmTb/nYyh3N2rcbWodcAzK6oOSnDtq940mk+7pesqCGFiKMTqafHcc4hxPmc5SuAZljX1UI
mkTTFkaMVt0VkwFCwSkVNx4eCJQ8uY9XksCry/BHd8oLZATMgUQ12zxIjX3167Upz+Hb8osXFz/s
4uc74VopthTvMTbRqkf4lR3CA+2hbdn9CTaWi6qV7Rex/WvvOr/nr5rwT7KFVC81J0WXEI+81LjC
U3ns8gO8P8j8AQopWPrmDCkLPp5m9wDENOWBch265EuUW0mop5KPj38AuihB13gpSJz7GryE8XdM
i5qrMCg15g61mwxoVPDBODv6IxNftDQdZnWGEs8S7SNM3qVPilGuZBJum23CGNDw8d3nBmKzGzbI
UaTs4BCIGLkF0HkLGAbBTObcGMuAvgoh2UTonTqCG3Q1+n8Z/Og5aLzlv7um9svn32hyyRuedvJd
SXvCoiQ/ZQYMCrzCVqUbIcYnWj3e2Wpx9UaUmQQIQjPre/WTFOnHmFVAbawuw17wKaslP51AZ+t5
Ilg6IBDTVglq0RuC2di7pxsnkPTuzgn4iN/IQb/6xqU6bikhNcFjm7b7OVqhPY4Bqg6llbALvT+9
QUi7yIGAs+LWL9Na8bM4FEi0Pf1a1L/yXAl67kh9vorLvieuyDxcjMR+rIxHI+H9Pj4r+GrDGz8V
8KaD1tuFtFqHps07s60TufgngANeZvPTyP5Hb+ViDMbDJhxpd4HhH2YRxojII2d2krgTx+/uMHLb
JaNGOicSJbR5tyWjZw+7DPqq+3IIzHhlDEEQ+6Uoyl9R3zTrk6BC16eCFleW9JdQsvA0ZL/FyuQK
GrdHAhqDcsdJv6tue6hGgFCVlXiMa3jsmUoaxxx7XUAJUwkMU5pD9RLhTTzLp+d5R55Fpl/t3r5S
uznRE5AMP48FysWp9jRrr8+49RS5OvuECV2XZE+eWo0lv8LLf3P6DvdtKCG2Bme987f7kt6fKjss
ha5lsGUSaOIcmuJjY8otYhP8vdk5hwMkildHmfQfguX8/lzqexj8hshXhKQaW1kkrs0IS5FHyLzb
jYqClx7991cA8pCJaRG+Opfmibps2YFajtKsO2R84TrHOEo5hGdX5mkQqs97ldQHfJTF9sXeS6iO
N8GXd1hYFC90z/i6zhjhGddX7Maw/dxRu4xD0Fa2LsxYTwl32aGqPMS99tjaLxhrVWkaaHJqqNnz
iL89pfVUFKSGU1+wV6SaVFceXxkLi8vzJaeUzcoBKpqHuVgS5ztE1hNhR4+YmfL8tzg9A6cqYs0C
JDsz3Bcemqtl9GdkNKXvL6X77endNfTLRZCZbtM70pfKj7NcGsUqG9YuNE1r3qVaAV/ywUorhCcZ
Y2k0KJ5SFsgyD3/xy70N3aFb+tOgkdF6quuwI++TnJi8GN9pJ/u+1ejx0hwg+Y/5dmLIspGK88h3
MOo/1PIxUhhR5+BgtxJn7XRUzz0D5r6Eg6tRlEs7p9ENgiRn568yDSdhC39K7xfpXj6f33xR0Zn8
/vfF/6z1/zybTMcMaSjKSW4g6HQr87QYMlVkTBFAvWkH21JPi713SmoTTGzed1b3qqavAure2k2P
Gf7QBAeJb5jhAsWc7OhPvps4ctbv+4mdp7EUSpMVJDvu1gIr1vuJdyvecuEYyIlCsAFswYHD/C1E
h1RNqleJ7enAdcgI9KjHE2oWuXSrjFnDpkMCjIYetXOw/hO3oLTScIgE3zGhQ7Hl/y2aIOTedtZU
BNVyq9XmITybOfZ4ZmleEJrO4RvIpmRtlPg17Xxwz3YE4xuyOyNPrgWdmmxUXq9bhMd+jvufMSsY
t+GJGy02TaqWSNHZ6FfWyqAIyeovzguxIuuLzC207nQ2uBihfI7XOZ9Yn5cK2H1GkXCfIXaQ8hVt
tk6Gzl11Y2XXlQ0H+yFmSRWn1tEihEsl82+PoFUOGJLyn/Sfgw79+ToZ4ngs+Ha/VIW/kt3Bfio9
zGTgezekcUrgnU4RGY8eHiK0pfLQu9jrysoYdh43VuIAbUkJG05C9MSlT94Vnz9yZref6zJkQGgv
a+125gKhM68V+BclmKO+/mhsCvC+dN7YjmA1xpuzHeIUCyUjuUAdcVBuEGOzeNLZPMcyTey5UoBe
cP7Sx0flROzHvRKLRKaKw2xark/pUX9nsMGWeBnc66eiOFNaNWUS7MpfgAp0uf9hqVfqwWePBOkQ
lZHYqTJb9yyQYjCnY9uA6a4d//j1KTEU4t/64D74iStgEiZ04wDFa63+yVYTVJ6cSpMWIcq7k8Fy
b1SkwlrYXvW0eajFzt1Nu77OkBRrgFCQp1Ezh1iJ274IUrCoJptOksM3jKelMjdzbQHjmHtF+qjG
aoLR/vgrgwi+9WK1bo2R/yVrwHqBrymW0hnkgbLMq9rf0sgoJGZLQnRDBYmok41YPZb6AylqmRno
7D/+8bX5OlKRAZCs6j968Sei4pjrL+n1JjLVV6Mnw/txVLdCUcBJULX2+VrBQSQOxXY0zLhr/kVX
hieDXnkxKNOLn3svmNbqFO8gHMUAvk1lXSdbdIGzc0EydC7yv33pUor7n4ddX7w107pVpU3Vhjpe
aytSZNCPvIx9Ri8gGhyTyiZFyy9xz8HMoLubzcx3vNMlPmzfZSnSNqh7LexieaAdkPGxPxZPSCtz
VEHwQKkf+22UfI5ckUy58cIWc8FEmwV/Y0WjPVsun59RkHfNUff2zmCnFo13nt+YbL1YfjKkG4lq
IW7iIdSijkd7SQS2aOOHOGEyDAC5LAvn2/01VQJNrgGRXBGeL0jaTVbOtbVTeqgBIgyqLIzR1Eq2
uTYjmkuXRj98fJDZJOdKLUow23QzJmW8jXshPMl29RfqPDENCq/PLhmGHYOX7rtmgZBnlVe9MCe8
JUavhUGpEZW8lda+/rapbvLgZcBqWzyGVHPUX4hcGfnUksvPlwuQDM9RXJ98QsTGJxFw/8XolGYW
a9Qb++u0moppewmJ0i/CgsltbROZMoZwnWvgQesRkgSZ6xvAcmK+D93FAVW9vmCFFt1OiC9v6SbP
FHZYDSdH7NCVvioq1BoAJOx6bE1ZGNXxt7Ukg8cbLaqTxLbEg5uDjGEKICDdbx8+F8kvYoAS/fO8
wUYioEmjGEI/vRyYYljCrS10xnC562ALLRxN07Tqqo1aCq76wQDlENurXu5qqC81+rKmzqgGLOpu
a6e9XxlNLNl/5o0Q2iU35McyAeI+ixzhpGjTJJk9lSl818gcRuwFwr2Wm0rjN+YXldruFcOvGp9h
5cWNJiiM8vMOtdYPouvbclslb9yq00/ESo0ScRzJecNHhGNJR62JqYDoCI5mAPrB9i8vie49N97S
YAa+2xXttO4l4NwiHwaLDUa2JE6j5om57Egkc1vOqCLcwFwrB31zt6+R+bNMVza004SvWeoMaxJ8
krNTP2a2mNqENP0Ife1D7oLCUBkRWTSqsaK5vt5pvK/NUGZw/xCfD3nyze9dfPAPDa0bvTA+dG4F
WT4Q+woa3dfQVL0J9uKhUwMAQziIslgy7mSEi5svxVXn7JEDeI7CNl2LhLWQqIIn+AXVE/UgRyXf
e9Ls0gHweOUPLjo7zQe5Bv5c69lNhOyDRXaXSAr5ASdvWeKKjNQmhibQMcpezgDCIYCfTBbLztWl
PRiwCRqG1WczfSrOaMwzRjZ3uJc2SV+K5XHIk9ECf0jMsSgMZNQFDfZw6uowWxc4RDfYF7cnyaps
MNh+TEebDk14jY4H7ZQFFzzm7mrShZHi59fD5ZBY7jcqN/QSb3OYYDKgUJ6J950Z9cVqJkuQFjxK
TITB+26JS6IbvgByDdhjHQMP0tZ/SRqktNbVCjsBy8bS3e15Ix2Awz+qRWCem3y3O6mfl3FEtT5j
fc4OFvEOfo2+4/A34JAJr7zwKaGQXV83Zv/V4cf5j1lpkUAUqZyfZAg4H4oqfZ0yF+J1iNE6AF7G
L992MFCnUG3sD8Wiiz1s25W2ow7jLj+63cVM53r8apTAzDYTxIYv6ujVth94Zirz9W492XEoP+an
R0CP8d5/4AaXiBCkRGBLZ9mj8h73siVth1U7hWVXQ0/6zLLLc4qh4wXQpCg4pmtF6Ky4kPZophCD
yfGVPs8r9T6ZKayB5IHV5tpPwmvLFVU7XNvAuX2vFdGd+gWmQJuoe1SByqn/b5q8uEdekL1pPYv+
9iMXhbB6bdKWLRG6BFSKq7fx7bG93keGqrY2M89aKEhcN+D08fvdh8RmjVLXOjviYU5l265ZWcjD
/DBSnQs10Ao2658rMtH0tkg8D8lSLhKs+IhOm6cVCXbIVixdvJClDdtg+oEVnn5umU7HZGQ19PtU
byegJVX7RYNCjf3GsT7y++pFY/++iCjcUt2R++czsfJXDyvUDTBTSZ6jSra1KFzYebiS7zx8BYbP
zp5YjCYr4m/RzEsvZPEx/zIuWlBMoQ9Re7Ff1ZV3o08xhQFwueIIODcZ8Z1Dcn3jFsv5LplpgvtY
px9tdbpE/Omw/dsX+Rx0JlkAOuH8MaAppSlIGK5blnFzJExMVYjS5kdlB39MlN4f9ZwvK2gwJr+X
V0i/DaoXqUvmChXaka7SQk82PAOp6vtP91e/cOC+rSj6C92cC65w+DacN7eUKWeyhMuYAI+oPHlq
7ZasX+1s1gzNlPpbz0bgGO1rXDIt7OkIdRu4yruxOq7r1e5T28Y9VwIDqgEhqoTYYY4FY4W81ylP
KDWbu6Ulcw1/Qr7GfdTW3t/X0fxPOHC/MQzmloKvibsLP8RyNqHxZyOQNuwrBDKjzlrp+KY5ZxBh
g8K7iNDsfh/RfUT8U746LdgqdHfg90vADPNEdG9NjW/k00QLjJjvOnjgDkbaZcf517IAwBd2w9XD
H1JvlI18pNrT596eKCSVld1u+GWSfaN5AZLc65a6Prb3bwnmJSJ4Ra8HYSTotarajLO4TN6FY1eS
luTQgiM8XRd4WfIwZPCabw9cXv4FM7foX7flQNaaRDD9xnLleEHLcIkO7Jb7nnIs/1iEHESkWBiG
rQ227sLvG1L9YTlVPgKBhdPZdiubYwn9WCFkw4YyEUqUgDRA6Fi+jWTHv6SQZVoOi8yQkN5v8yxi
gwjpiyWdEpXuYivsXCHStW3Jpz8ie6655V8tF8PePHTCsIHV6AZk3+qyf9WQkkH7Dn/ZaXYBA53Q
5v/hvnTBU6x7dSAPdWMZMoAjPPvmNdNItx4BiSwbD2AJuYW7XChFLOzyihy+66iEsIVwduJH+HH+
KslZf890V0gPTGxj9ButMg7lmfvNocHcWYhFGWLxRNdRZWI8q59C5v3k6tUQTuInPak+gEcBj43J
Fhnz+9P33VclUEVnEbwX5IbbZKOJtr1w7OtQbA8a8H6BjL6uT1oBjfYopihQZbsYSgphiFMbi07M
100XRN7yuXapBZpmbJT4a1sqp6fJ1GETVuooPE8L6w3XP7fcZloesH2YAZKy7idcm744sQMU3GXK
LjCXXdYyCdcD20iK01KaCbfmNTOAH9AX78pC44gXZy2dTi7afSQA9V9m7reDrd/TQcATSdNUtKFQ
XdjKlzm+70RS1aCgigU1ucofjCoGsusMqhtWBYwmz7MsWIWk37/DRQAgpxqF2QpzIEzAzkTjwOSu
zGiWz1ZDI33QT5+riKssOwHGG9FSc0kBaFGkU8c/HUyKN7terQbc8EPeJw15ohZeCRd8pkRZBwO+
cOXCWHqfMpJ6M39vpC5NK52gtP4RZX98VJgMIHrmpe4KGCbQkWFhqi3xIlVTpvtSNcZ5x6X20yJ9
RNiUgpa/weNK/keg9ntWZTYyPCtjbmoak5sYlqUEago4SmqgM2Ccot8I17PZwvE5mi9AnOXaCxYO
SM5QC/QugyxoZfXIDQwiYqy6RzGPjSCO4vtC6fYLgY+Bwis0J3XqoNdcgKtYzZrvFbahwdFWZN3B
dDbSmqg6cRES0FHQL+OHI/1lMRQUusAXs9d7zLAdDWPzi87SbEtByge27obs8gC1IY03Ir2PBsYi
jX+YvUKpMOj3MZV/D7o0rblT8rV9jC5uoS0+meHI50inuMoRRyZGlF4+hPd/KuhR00bwRnW8w4tV
8l3p+nh5gz2L7oY79Ev0EGD+xANVvuOlGeQ7l9cKUD0XbF7bvIOuodly9idf59b2gxKl1mmDFlUa
iMVZuZSdbUnxq2CB+SO6EPbvEtFDyb9pK6eYViqBuHuLIjynCEkc9OntKW+XqgP5mDAWN0jh2D/e
LTVAqQ4wZ5SqgL3uchGkwd+VZvkBl3rELhMGGWozYq+4dU6Y5fhGAp5dEv4aXDGcwB8oExWgH1oD
wEU+6fX4ypKQMJK9tCic9BL9UHPCkxt/ieUtlqpMxlkxiwx1qm1e0PGigEv1XkgBuKO4pMp68Q7G
i0F6E3oLPqOYlXmxwTFFeizkuDhJQzlTWI/Hg6LLqUHmGMAKWhH3a+oY59D6pvGTNuR/dQqjA3QT
vfyIK1VOIAkkV3BM0ZeVBf55HPgoXwqfHIKyaUqCaCEB/3zc9vTAJafDBIMfv1CCe51elZRGw2lx
9NPYggYVWS44Tg5I6zR6KH1Dk/Df7jaGBCCQ9vJIW0C2eOf4wsTf1EiPImq0J4dGK79xMlcToKnJ
gYR2wnP+o4FHzXgHU2lGgbNh5/5+KkxPSuqeYbz2hK4ofu9MJsK98oJ0Sb2K0s82MgG8URBiQpy5
jvEpfRTc8cq0c2siNT2sCJAT22u95CLhaqKWToEf4+sfnIvzB2zZcY6qulbAeSf4dvGguIqozCng
Pvmm60+nXVQqB0mhDF4vIJozLowrdBpir/RQ6hrYITUYGcrWqSGoQDLX2mvVoJKa1KvlD5STeWQq
Xw9qwqvTnfSSFs/qSZjdzjNM8qLQwYqh/JgjSWbgk43/wTdqYhnm7QhByjVhx/jn1wtPRzl3C12D
QIqinW5CnsGbn/MPC55RJHCGaHpSXxZWO4BZ80cnw88fcumXvDeQWglZQQjrbGhrBnr5sYtM1ad9
0OX2W6vHIe04m6ulyna94XNuGAgsHGCLaf5BeZyip5gAs4I76jGN9uE4JJmHeIEX/E0HR3OtthD+
abpbD9cMJDpgX/BmxTXsJMd8HggyLQKhAFFqBngY4LOlZtrqPOfOWC3T2WcLhS6st4YAbJJ8TRav
uXV9x11ZmWi/l8Vi+100yF33Z6Ip7MZjPO/ftZp/Z9M2W3N6Qq1CDkcZvWmmby8JG9b7BG25dPjO
rma6wlKGubt+iU8/weaik/kwqW7VjwIVo2v81BbCvA7MHVZze/IrwcIKm4VIBjq5gaLNNdnLcAI8
PG/4h6Yp2XWW5rx8GO1sjNB0cXAf8CmMNZi+IOnu8XV92rP4dyJ9DE3ZcvF2nWM/Tv/Ebl74w3Jl
uXzFVql9Lz/WuPQaEGCcEWs1EwTSlWm6j0HajWOh/r8R9oWZWfoDg9adxUcCLckrhcD1S/6Li+Jx
N/FwSSCZupdGDXmdEyObI/+uWOO0yNq8Ozpg6lflkXqfDC3ytbjyR4I1r9QwuWVYAF3pDCZ81ght
E/OhWWuIvw7+8nbi7YNgubGQTtxPwj7IsyaCLEbxkdzzED83yFPz1Q/Vbk9Rwt+RC7Q7z/Z6ga3T
vMk8/1F77DevDouWlf6FlZrsNUzBnLoP0UGMeudGVbevoKw0ayVKgMyCVVbQ0KS19zHKpACdxJPm
vY5JKMzK7uaaT8Q62LFSCz5CWGJ/bniwstFeqxoXLlu9mYF5qgWhlZ1zsJNp9N5YDwf5e3jBNy9F
uuSmlPdiUyNWZYTj7kz5Gzkkn0rNJtkq5Lpg0Ox0/MydWItnfqh68A16ULRGWRVkDKeZwtf0QCP+
+3Lj8jWx+YX2g6tZIspAAb+ABUpNtztcs6AJm3kxS7hm4ML5PGnf4jzOUb5yz/F7jyNZ6IHfiI7U
oouL2ztvkN1wk0ps39FlYCjWD44YTavQ0YYho2TqCS9qNnq54OEOSlR/SOPTUNCSEbK1jwFoIjJh
YAtQuozjKMSIEgWIFIYRNeB/u+h35Np4t/mUw0543EXhnMgjzqHdjiOnic3v80Hcnt8mIDybJlWk
rYD1CLlAPeNeBqV5NrqcPuHet++kLbJD917xMrqtHcvN7NLTJm51j6QCPipp0wRHHteAbvZsL7Lu
2nAtGNnPFRuJv/STzAnm4w1XNF8FTf42Y24AwWXbnUizPwy/c4hUakm8/1/4MWA1KTgC7QR0umFO
qfccdkeJb/kGEnCKGtAOQ2HyKKs17Rnm7i/9c3pIUU7rJPUgxTmQ00ZlnKs7lo0EFQcvQWW1idX/
lHcOejT2Y1quegPrn8XDeKeYhT45zcVBCMF7Yr7iG/cuKeu9RN1W11bR8CVDr/BJSQcZEzznULIs
yJ0Z+pguhe4jRM+NA89maY4yv0Ju3hKDKUzf+kwbUwIhJHTf95Xm2dSyu4qgo39oGcvTmlfRZPlm
Kzr6zk3z0JbMfkdZvwEcXpd/fxlg+5NUlwUebjdFbSZmKkJpxWK3uZx5SZ1Qi0Zd7PkAwpD1Xj+u
odQGQD+udARawqcxm58KXZMJ7G60GwuaSJlbw2UILqyc/wb7mG8ftBtVxGL6ApRTIpeKpwHsre9t
OgDdbK0/5PwEJVcafp7DVwDpXyIwa0l+/6VZVVi2530NbHN/54TLT2P14+W2ceDWPkLQs2/ohtDx
ufAFHCM8PZoy0GNTVukVGmbMiQASRUg/sKVBkcf9GD14bv2osXYSqETd0PZMZ1HmuopcWgLtjvfc
ovuia7LwhavnTcqFaB22t+FxvOzzjABTtFi7j6Rr3do+M9yYRmc5eUHaGWC0Psqg130cCALnTx2w
OXVDYqYuoq6WMPDXrx9bLCEHezGhjNYXDy8kbPioNnAhmLv8VxGULFUdCIj0C8LV6mLIRMIRnSmu
sGYFkjo1EEVqBGFJQicqq/E4dMgg63mlt0KygV2Rg19iVK/tOkf4Top1MZHxhs9VcuFcCR1c6dvo
PMkGHRMVAkbjcUd2u/rF+YO+88IpDDI1q1q61dWW5+yiNlcFaYG+61iGWBhJFXGdixSTwHaWK9kc
icux163EqF3Uc1D3M1VQ9IWciBI1Tu2JU0EMfD9rWiehzo0if/4DVKlU/YwrUmWbBvjueSV0MiK5
1KecYU9Ecj+05m4BcYNUhD6YKBqrFPNq+73D/m9aKDT4lIoSoriqmcfnpyzFfWpOT3zh7T42OPYU
mu9sDpURpuho8xGPADYmRZpEt8uQ3tU0cJNejc5DSzCY4IZeLrpBQcKbaq05sQAIZcY8THopZNY9
hv8clf16FmQrzaM2sWl2CVI97yLcPdZ4ciuM2lXxERrLRmqZ7bSPcQ7nBWcueKYLhu8m/+YjPDMl
nK2wvVxVWpeBcW/R7TEZe0umsrTsOkN8Gy+0INKl6jwj++mshy5ckQZiempGt0IQvLN3on21h01l
dnjoglONlwFyvrFrolc17bDmaTwn53zGuAWGQNMm8dghEQ205/yw1OwM+IvJkqdoADarOqWRFNrV
VbP5tMxVKWobzqP8qeFQSs4uyqePZTgmjZfDqTn3hE2aHJOE4RyH7QbOKN4tOIiJUAaSnSMw7moY
wweyhryHi7wUOPWGT/sBRciJEdMCosfmApWVKKxXZ46wzMaNMmxa7DctmvYhugp0DxasUKsNrzsP
hlGemLqzwa4chMQISBhJT1KIURWyqOa++sezbV40qM18Vxnz0JiSvHmvnFuT05QsK7apWQr2gLcl
3r30gbRyLmnrPyQzp2j/sebvMKP9qlMGTpf5sZmxKR175y4tWO3Js4rXuY0mt3MmwNTbmWiXySxm
WRCXwENo/e9cmNz/chs+WJYXK7liv36LDNfmtFIkLy2wxvlia6xD1dLRNIa2kWVvoLvjvAzpUfxY
KT4ZQbbRNwthLL8nEONQZNj8KwwomwhwIw61tIp4nXwd8poe5L4mkeXllvkpnXq6s08/D9lzh5qw
lFPYwJDmGFt95PijCUc0yyDqcOt89VXtCngYFSLbFXML8aWlNUZKRWeor4F+2pyL26ljBdBGQm7K
wPC5QZ63JwfA+OfaSCRhVOlcmjhhF+h5fRMZjOR1QOoodeDY9Nulpyp7L4VCkLzQkF17czqUzCVn
CphxNRvXtXQzz8NJPz2IVhXhnnBU/FBcNlIZ0YgXeSHZsu9M8NG1lNQbm4YYM92VnzQmqNbAepss
jI2OuAaz0OvvNltW0lldy5OtBOjTfeTpWUCMpfFq9WbIzbJ7Q71D8c7ONs+kpOuw0NojHOH4Z7Mj
XQ4KL0by/rnF9iBqbFVaOruMrZlfQeXyy3/oqgf3534KPnQGXAuiP2HLebpkxCeE0t6x0Uy8DAur
Jx6+K/bTulAGd7SzozB/eApw1WBpdm8f5hj0Ghlf1BCYd1QlWCsuoEB4ih34DhPSv+IdP2HcCTYV
7xVt24ssQ1H/PUvmwhAd4UyiId3Vf2NJSfyzgdGh2vv5TUXfXjj+cOsUiPginz1VskDc5Tyil3jO
/NL67+5a8FBgdEIMMN0GQlSZ0E9yDip/2AYylHfhYWLTrKO7rVwgRGeb8rsnwzGYafe5+m/8orXb
VmW3NVKy7lKX8xvX1KohEQlp9xavjhGkk/vrDgg5vMWlTlsg1CHgOLyBjHXw622wy52C+DZiLY0U
tVpnBKVV6WMiSAeEngesMwBHDUPjSLAbK+zgLzeQ+JBJrkW/9MmsVO5tM5McD/hPH1Cstq1PPTwD
h+bLXlwfsOihF7tH+TWem0YTVymVyrYCJGspbrf+wmyNPN8bNcwQ7rF1fsBXlcJwqzPA39/eQYm5
DYF1jLTK0oUEdptl0ehbPBdUJeDbdbnrUyK4X+Ob+Hfmef+8OhnEjVYtW3QKDCuBHpcuwx0sDQ2n
FlG7eYmGHIWSIZk1qDmWmsO8h+l/ojWxFu0X9IwJAAFYNG6apOOdjDmjdFi016VzFMrFE23vJbER
RvwAhTYvkMT+scR/aqzi7djyyCfXLQrZnbc8FoGUNAWRzBHaz4IWnJbtihmn1tE3mZrEScfpz5t9
p6ZvbN4lWIaTzeu2xfDZcsU/+dG+Y54BE8GYvsiA4cLP2NaQDeziCt63/AVJ2v3kBR7IbZA6fzX8
l6HIQXSS5jOkdHnW4Ibr4r9jZ4HPiiRU9RMtgPja3qx+d6LIvcxbvkE17qNljgpNfj52CejAxTSs
Ac9A37XfLEQkYZPvmbxa89gjoQz68E5fkT0gprnBU14uuDgs+MlOpcwmtV6mDSCvudNfktU7jG88
e5X+bNa0TRlkYKUfk264vBRPv8eZAYglNovOW8yhaTOU1wI9+ybLWtGmlUA/7Kd1LiRXOCLOugeJ
1K0VLBW+FlAmd25r5wy1SEoS8YPXiiLAtQj74exRJSi3ANcrDKuxOrar4nZlOiafg9JnxNIfPVDc
RgttQSzN3WtRJKazuafDFrFLH7cYAN9iaA5LhmIlhW3bot8US0Omfuo0K82UNwcDE39ZrpuDIkhP
OM7sowdtO+IG2UmM4R0pf4hjWkvhqD8+Zg365VEGLZpCGtMw7iEsLXH2SXG0tSQ2XTNTugzJg3Sx
M1Wy2HJ9U2Y7RmjDgkl3xTrfaF9346OqffLA7xNrgfif/NlMvdsCTY6tM702lk/cVvpFK24Z2xWt
JL54Hc4wtUC7Ib0E6kbeC7TK2gc7KNZgGqERUByd51KWqZZ10mKoJY0qyDGP/69hf77MpSQHgNCN
lGxPfm1zFVY+9sFoUTP7SCLGmqQHQD0brC0URKKhX/9YnZVlEDC+8Df4GaHA7o7jFS6/s3uAL+XB
0OjYb7o/PMELY3c/0sQatf5V4CqgwduS8AU1CKevjZdCZ09jO9ye0ctSlBsjyQqboho/WkKdU0Xu
40Gv2pCfFUnVPRDjrqlthBgfP870iYjdVt3tDxfLuaaLClpkrOxoPSW/UChLZivQyVPdqkAtEK9g
lizeJ5CtgUWyU4/UVbF2FWqOVnNRHsr7p4mIKGMLdPcT2GvmGu7fOgBfHBH4X3b52MfukyTRK58a
Pj5pJ4XFQ+DCVMhXnSb/T78HJDQDLmx6KkxPPEgqenknF8LRUGx3JGrOSkJynxpVtQVJuMgLJJrN
Tx0Aq6avy793DTFx+VWWzkxtWdKAl/9Wx7wBTLkQxocxoFDO7gjfPCE4PEUDzdU9wc4ki7KY4tSz
74dWuYg4noacdnFoRr5Dbj2aHGSWA79yp8rKa6GMaNAZn0IvqV1UWkJWToSp8Kz6XG7aOIG5X/Ci
qlqgFfdgQa/dyjoAieK6ZNF6CxkYMKRPyUZPSP4OdsL5vt2ChzqyhhyGzYbKat+Aal3mSXQ1t5oD
7xOralik9CdyTzEGvqvcgaShGKPyHp5Bs5i31m1y7bcTAtApjvOKF6ncV1YWc4Lt8AWnD2/+ugEl
DMN5Ns/v7DIR/tCP65Eozlth3VrqC/FXNmsdfXjZpVkA84qfEmzxnspXEsd/eZdsdHskLTNgtMB1
jC9z8rghOnVQpOQpn5oMaHEz6q2/wigIZfWsEUb0XxRuwj8dUEtGEouAlxdE8XRZty6SF/Bk2OEJ
whoTlGCOY1wM3+aFMG0l48/loJXsNkRvCZJoGI0JMzBrm3V6vyCJPoM9iFeVrGTx0rSoktXckFow
FUOYFq9SWuV67K1zUV/LGp7D04yxAZc/sXRaYwd0Wjct7HrDFHDZNw6TA6ADzpSNgn/h7P6IPthK
u9diPIxo3P0B5oM/LfBWbml+XRuguUs8TIgNq23FvQRek4fw7sQ2iDwFyHWfNyI4B3/4V+AL5bO3
l+OgxHcAJa4KI/WANujF4/r50mpt9d2RcCxCw5rNTEE+TbAPcz5zSP5k2KeUDaabpUR+qUia7soI
sxenS8ExEPXWcY+Y+BwvWCH3XV/WLdHH+CMhdxuc2yEBW0vIy/Y0RjFj6gRk4zGRqUSyN3pT1/g1
11j+M4+O7WMr7ex4+s2WY4EZnwMjXv+MoPgzw5funF2ReAJx4WbpBGXtryNKVK1KkBeejQQs3hS+
N+mDaR+4fvr2x+oa7s/7B8nxQ6GK0DIL/H1VpIq1bCALBAhjSoT2hsvPbdqWIOxYjn0qbz34W0VW
GJ1FOeTb6afCjUBCqT2ViYbMENxx+2EkgjKG+1j2ukqYnvcMMGun7B3lL9M0oYQclsbQivgwNhEC
RDC4nsNnsDnkL8ViW15t0x6zPjyYgupjRA8zINk/pHKci5mysl2vJGf01e6d9B/Kp5caDjrMGuk+
VSU1jBr+IxwO2X3ZFlYvwWqYbwZD7/TOsrltEQ6hFWcUaUmF4kqEaQM4nrlY/M+ct4UF7CsAJbrV
24wctJm5cLhrn2HtET4270utXPv2Y23/r1DaaAHjqIW97sqmWazjnEH1tYQBZovIIcdLflPffd/W
aJPyz34woAeKYA7zvWHH5AWIzE5O02huiYzkXbhXjpKa5aj/mtcMQMIGj30OwhLPV9G5X/IlnjqK
uU4+pEPYaPFDs5Y8puOq/l+ATbaQZRODMWU+SuQ5FmYziOsC9CfZglfhUeg+2mfv65//UMX48uct
AzqJTrIeuyn7XZ0i8Zj2zaHoMyFMjtEaufAmOnWZ006G54eEmNU4CXG4cGSBxUQyDya/92VSWPEA
Dk5fFeN+pHk3IhVObuYLwiX0hJ+ByC1cI6YwF0+cSbvq/waTthuSvMMwfJDr2XgmFvuWh46vJyyP
AIPumjBl/xwNVKy0Q1hO31UofLD5UrLu3MpqM2dOcm7DXlzgVS/XGMrxMzNF8h15fRn4WVlwNw0+
EMpsJVZ9s36jexSew6Ywz1QiYl2sc8FYfUVsFLH1x32I4wXquZdOItmO67z6BWKMEgW07eIXPPcW
m8Bdvq2vPB4BTCjnouuNsnbIujN0OY5h/aI+ZkNUtShM04AMr1rDOZPkzIXtYFPhqmSS7q4YOl05
RvcIdLHGr585+nO51R/RQxTzcx2mELNTUtKV1uSPAPvxeZSk5Zy12h9lu3t2Ym72lG1Iz5PdiJxd
LKV+TTDX7sjDtub9bBq6DoSGHKXn1YFkZ8X5sUaYq2MjCwL3A11EF6HBgjX+EHFCIekkmLCx/WPY
fyMosntK1EGUdr/ITMkyRVd9heAsS7l/MO8Pd1P5Wff3ZTlhXYPFu6BTfRRurkejkAxmLjM/elEW
EthPs6PvRhPvwYMvX/hLwNQ/FVhB5Jx1v4UoTBhT/aP+u3qpRqWGnngtsOZ9hCqbi/69B6FWvzMb
aXa/wzJ3Psp3k0gndw1hXVM3Bu4sNueqRM2mHlUzrnz1MX9Iu2DHGXVzYkQp3SdkngJVhJmVJHIH
E+79N+K+za9GGlqwJwsKdLwZe0w2hd3L4mgZJQCXgzwrOjOeiAcdjgDnRADGxDf8uUNQQ5CK2IsA
67zvnsv9kKb9LtVGFiSMmCw7Zka/sdnJZnQtSEH8RYjqa2TUi3jhc4AMFbViyRsfyROUJmmepKQV
3BHB6sgv6j0WxoYtVeGOyXskml/dBqybArJHQDHsINGfjQ9DkmuwzOl541lBCIWyF1q4qPDfsI7t
t1xSRGRVgA12jSQBq7EFpHEccsbzV7zbU3q2hokk5VV30PpvYF3JvK5v7z4GEowFS0zJbyh31lGa
6nRLeHErcfEauWOcsP5W9LDKytLuIl1YcWY78jAxAK8g6Bw3mXKIRN1J43ZScY+ZuF67N+I+G2mt
Zsdqm0xaTrRWphfs+QlXneYrq9eEW3ZgwqPrmiakNSi9b90ZPjPjSNqoaCZkF6sA1F/4Ap89zS89
3BSiohtA70crF/+qUOYdAdV903r8KAU5K04TvhEj/aML6xCtDJ2OSGjvcjZzs4Ra915OCEznblFC
lZRcIxPiTsLWJkqqcQ6HjWMWFFQAhrnpImOTWSO7/fWrnRyJj3tP4F3tCKv8fhAJB8jcG5ZOOP8l
16KvNpG9DSP7+os+kSEBR3+1mgS3CJoUFRiCTWMuhmn+UrpmIqR/R5MBnswfQ5NWYCZOp/p8yLug
yJ4OZy29Bs4WEub6kU3X019MYgWaEpck2upO7B4Hb79ANQgqzHhR64JSdTmoP3ewNn7b9a8DZtIQ
mil+VVKhjsppvprEgkZ87Ye7qk6/PIDZMQN/x81L+hDzKI6PP4jwtwShzz5b3WgpuDRKp75r4qhm
9PLde2ItEPNQPvtVJQU/A0TYNm5j2fa+cA1zbSZqTH5OufP7TWeE0DzNqtePFMZBGJCJr+/0F/sp
9m0VwzapRm2W8DfP36aBcDX0+IvKbIYv59Fi3T2v3XyjKt6LIE/N6c4l7etuDGVpU6aIbKmCTmzH
RYvbZOxu096MJoro72CWuJSDpllLF0imDPi70aABeinb1kzKUYkklPD+u8v7I4B5hgbVopVeTRCP
aOmeujb89m0K/o5LZs2epVv/KMhlf7h8LaltiTMdOOjLb/PISEV1mtsR4rvHNn8SdCDy2LtkHNM5
jcPBHRGAscnBDNkx3CgAxmhaHLyn2W1H/g4Ft0y/smdE5ZPAaYo0J5d1NhiiHsCdBNvoGBbAmswL
o9rosZoV18o2vghsQVBphDgVgJNiWAd1VOFzS57NJS+hXxQyG7cSALruFnTpqKxijSz5/ZiAFvH/
uadKxkln5GFfQ2fHmgV08Y3BGflEF4dfawfk4gSEtE8jcpsBiso27V9gqFJq/6n6wDc2C415TgS0
sdip2wZAGbQH70Zs70+mkNKzybBE8qoi4ajBi6CyB/2rKHM2AsX7o0ZAMp+cm/gN6kADPWNxTlpF
t9j81h/KtFu/OE4JK6+4WRP3WQDS4zBL6eWQwxtmpyjhsHzRhPCxefnpBTpA4kdeGHqQfVbJz9DS
Xo3zA4hhSD7iLLrJ4JvyOgClaIODi8xl/1ILgHM1TRBJtQv8OTJ4qobuulPl0ANKOktLkJS8fxUP
1ihOr5Fw+xLQRaEtechNpfgrtRdxfGmUXYgL0TDHyZfgpZNhTG/1oa5xy26LpEjSrV15Pinj2Fv7
Crjh4NArNdtwaiWAIWrQ5UYED+cfgfS6M+QDa+O6o3GkQP34WLahmRurm0ujbhYzjWJLjqWPooc+
/UhWxTkpy/yXk4iJx46EF7tlh15IMirBMldQ3RrAArgs4GY+e6fkBS0Q1lkSkU0gfP0WIs/dgRVK
xHKFbXc8lupiDT36NkuHqGSnTzyx5XJQvMqL2tHy3zURiboKjm76/CJlugZ8gXMFtiLQVwpkKAmk
G9GYl9hMkr+Y8VFTRZXUm/+b9x/qJO3GgAu823HGz0BHv9UuQfqufVemSiq4amu9+UP1/ChJJ2Hw
/Vlx0kAI3hVUt3p2sjeCJvDX1XDP2PwnALqZ5ZQcaPxqkCqa0XTg2Gs5bGanCfR4obAPKH6PpdLs
B6PhsH8GkCCVlyTclYioWDz9V65ijqKhw2rNbOpArFRjUy5YXmzCvLrG22Kte7lpaQlRXG80L5Q5
NANKKh2KzQBwu+fFCodkuG5ZD+lz768k2aLyoL2qRlU2TMfO/0lBQatWTi8rCjWex7IlxocCTUVf
ysUM9YFhXoHtCT/9sgh1xM1HaPGZnGlpQUTOeI2Pj/d9SsQ4yIMpXdHmGvnNH8A9QeE9NwNCvAr5
zNXBp/GQgsoijiwrOk6sPDkMwJskEG4esVqOZian2U9kxqafdgnPs0iYY9NN8SalEyMi74x2wGU5
3W44uj0cACXEVK6NIw2vo/seAUGQxXue+AKeHwCzg3V4ZReSYXFkIGXoj0GraglWXc3CRFybESbO
0Ik7CX+OCYUDRQnl6txnEDFie2v8rBFzoTZqn+zMLte0PlLGV7oT6X2uT99samKY1dnoNpmrSTwh
kxenG9K+8NZ/H6TC78TGGH5tvX/QWCCFhaol/gt53ja22bmHYZsj7AkLzVwSvfZflnRXruSwWX3d
0K08tRbVjxEjmGzduvw0Z9tJUxls8IGlYKqtYE/Nmt0XEYmt5TACd/8I2hNHwIw29qA3T90L5WGL
oV0Dwod/EXyzcVc/yeMAdrbVlq1E32A9S06tY3AWImGIVqUUheTJ7Jl8Vyzmh1n99UP+QpduFAfT
6Bu2agzIQqJUta93GIFpetuMa7wcPC8qqH3+Cqm6ogJarsQY5/IWxEN9TuqSWXA3vlR/aEq4jsst
5Ivtwf721GaY6532HrTbk6SydCdELSvuPsw9KCTEAahjE7soXno0AP2BXkp5hSYEb3UC6PNxNBrt
vQ7+H19+ZtZaZpifN4We2TRKPGxAzm6aRHgGgcmHJ4jXpXYNpvx1UhaphKJ9CXR8tXv8EDZQbkjB
yr2dU5pZ3Cz61wFezMKaTtJR0VTQuqfgg17aelgDr9rOzS9sfoUyhHvlebREO7jj8+SiSKptWpWk
0s7p8GxgwEtd/zKmk2Z2plH6uyWS9e2yS4zNr8+y3YIO2yZ28rsxtJ00bXP8mj43onfslYh335EL
+/eAOLMRVvHM4W1y2zVqXqfeh+/oI3Tx/ww8D7/cnrrRfilGUjqqIqICawcjVEC5nN3UbwcSHhPQ
n7KhOYyytETl4vTxiK8MuGTyhqG48a9hu0oLxTgbr/ZsPzD+TwGLaYS8oudxb7u/JJOoKlisKRIE
/78+ItyNrTWtHxmkogTXY5pYqwb1UdYd8e8QTWpONar7neDgWYCUahyoFUzPi5dtQUob64IkARFw
t3+GiC7Guz/M14f3PoCA7X6ru/SKFseq3hon/duZx/WeH/z+2t7cKRiLKCNUtGnjr4bL+8BsLi09
NWKgUHyBO8dKeys7AwQpeSDtcHmOn9Ggk5l2bl5HqmGcBWs93EmEBtmUZpGSY/wN9J9EZdowrYlH
NzMgW0YyX5ATRKVvaf5tMEShiQwj2Fp7jo1BJF1eK4UWDNpnHbw5x1btW/H1HWSR2JPOlM4hAOc2
9esfL8fnr659yqx7g9Y7zeEt2sfO+PGQQGvZdxION1xJetjXQHxGvGorxrFTgZu7ru40ptRuePGO
+NpuuRyaz/Ohh+BVr2yK4q3e/rLv5/MEI4hP2Zb572tsrBWDGZaXPK1k7PG2RbUftRNQrufRTPdH
gpqrKyxOagwfedSaVnmXAn4Z+JAQ8VLCJloxkV67pRyZ8Asex+8GWntar4JD0m0fZynJYkbYd4Of
Kfdi9tCkOe0ailF8zNRx6tXshjks1xUqCra/kWf8jKk2JAkXQD6+tBcPYFDqFuX3EedvUOWZYnOV
jqnvIm00G73C7WGOJdgqiWwQjpnY6QGnDFW49p46AxBtau50DahmMaAOJW7jKZqjGYuifE/y8Xy4
+di2UKTtRHOG0AkITlZmLwJ//NLX/J4Fo9hvAlVK66I5ETKZpSQOCzca69k9LSyHCMAoUlk1cQgh
raOldN5+4jsJrc4dEMSL7uhs4UiytFGkmFPb5Gk8oP0tmHuuVWL950zpj2w5LcIp4I7aJ3Dw2eWS
/Eg8YJpU9j81FfnneKC7cZz07dVNzj+rPExDHsjiLjbMW+b3OOcp3oQo7XWW1pdwNtvKLQEDxTiO
AnkKUhgyEJIfsiqDNAVfvBs2vlAgphzdE4uGCq2LC+7IehNKmPNYr6fg7tu7wECw5ChBGFvTooNT
d/e9QUuF9mppICZWol5EFHoOXL4hMEi9TMZte7iGXk+M63PSgTiSjysihS1x4cR3n/qrveBzARgA
gBhentG38poktUPG0VtzIYwW5BPGBI4jHq01KdesCP5BLlTgyO4hfOQApjqF1tQgUinsOGDH73D7
Ijym/s17KXhblxzNm0pQxYXokMqMAO0EY+jkWpYT5OXPO5UNf/Q3UUpnNnbabY0/CAaoxxnTyGjY
r0AJt8ebEjw/Fc28Gl3bsZ9BReJJmA/CxmZU2Y6uLOyy9OpNGvZAX9sk33j4QDCW0Grg0KOtr5cN
wcQqy5ygf3eO7+KWbRuI/1k1RMSqOiGMsL/jFRxRBFRvP9iT+DTIDRTjNun5bm0x4Z1FGclkAqyp
A8NgSPXw6JnqRZBWM/c3UtIUmP/xy3FG5TtJyNyfJqmI7ASiYwR22GwsSvensO9c4pXuHc2d2t+s
ylBF6hs76EohWvGdoDhylEyY2zCvvj09p0/v/XTxPyIKSaG4dta8WivisHodU9MiC9E3eMIQFjxh
3at12AhUcqYZzNRzP3UlFvR7z4XigegreppHAQcjd/YKrputlQI9q2CDriI8orc7ARKfZoAtnOOH
ZBR6t1F/dEmR+bEcfHuntpUUY1fIXFkAYe+qDC0DlX2CF6oVLoyv149v0DWTO/5G/AZgW+wFXLMi
BSgIZNM6Oyvi8EQ6w00QZ2+zYINgBXsl1WwbSOorRbQ22UBhQWegE48MijN8hIQ7hjTw8tzS29e/
Nl/DdwcR6z2ZXokPur+u9i1B7zmUWPvSdZNOauAosFbiPmhGuOTa6qxhokbVTDCjJkV1El+oLssL
jE9pAq63Iw+wTPf5drXH0R/pqslsdAJj/nFhwv1lqzCbEWyvbQrhlHt5RZPZogdiRcBTu2B6dE3e
CtsyLooMO1F50pFD0Pkne2DH3fjQ8P0zJuL9xQJoOjHabiZGfUOwjz6OqE67Yg1fwXYEDT3q0AQR
aB5NHM8i0DVsk0VxDJIF2ag+S/QUA3pCgEwGn3IPyKRuqUhbUMkGHyZJeMD/vLMnaZro0090yvVB
4J3MhyxPo9vc9qyEsZ0yKQ+VrPRivnBRP/UKZ4Rm1/WhtkceP8Lyffa6UPtY5sg3rRJfKWEh7frq
lNiumiNH4kHYl1RInmlq7QoHqm9H7GH8FgqSGLwGD6qCK0Qw36VvEiXXPZUGa2pm5iSalLPk5E3b
9Fij2+YQhYRqVzPQEofZEGSkPglhyi1uk7I3BesECAcGk0BBMrbpX1WRgd1xZCOA4d/Fz19Y7SzB
TMf8aYiVNs6Q2XndcGiHqj8kfZjz/PJqWZVA+8FK7h8uSA8DHjzcLCLHWX/nPgSWNDExloS/jp9q
WabDOEf3mb8WcxU6GuoCuIPJRLlO8iOqMcVEGt0e2ThL+buhPAj9kRJ/8896e6lGDD4PoXF3NTL7
a/NqzpWZ0OwGQ52jmnHWlFQFWNY6g7sKMTEKYQjrZ0cbED7xP6gq9KmLrx7X+Z1R2k8MZp6TpN04
Wjehueh3y2/WhQ/4d1DvpZk5CTcet0ZKf2PeTqqIjbNoIQ1lzaMAMtwoWXLtjDdWg5gHijMoCNGw
/MOWYvrpg/icFhXuvR6jtFbA2C8m2p0QcCzdfYDY4cKI36e4U+NOb4gjpmmpCgBc0z/GAjRDgdR0
aoeOvIKSuS+tW09LG3zX2OhTGCGM4z0Rd4k0n9+lwLK6JKuNF/on+KfjUQObzSI/5odMpn8Lxb9n
dnhWYVX9DzbRrpZf8RRAH4jJzhx9saN7q6jUY88npcc6t8SXJw2o5FXldxJHUL39W7Z/M00f0vtI
sqAW9DIWVX9RETSkE218kYbYTm7p11lEKsiOksUbICEe3ZQvB655OBmiqkEXiHdxy5yjeAXMp9P7
X7j931qJ7xWzg5gTC3vC0vpDuEQOTtaoEx9OeNQZNrdngDJh/McxwhbH33NkXT5+Xo7ZhfMWv7p3
QYeskdzLhvaHhaZDx+Rce5iquWG2S8ipoRVRJwiXEoQlJe/56eewW4itEsEIIiDgc75I/HHyta8S
SnnirlWNPesqAeMTXGjFIyKNXckZybsSGisQGWkTJRD+O1CMHX4ZHQ285AGejOXnSayTrlNAN7F+
boVHEzQJR0ylNCtWfU1Tu68IsiOdo8tzDl8UYBFn89ApRDHdr4iNMj9t3fQrvSYmq5z99Wl/pw5Y
1e9uvpn0RCs98DPFcpRl35eK2i+UrCSmL6E6MeK9y3VgEAK2VWctb/jw+7Yv+QK5AO4ORP+bmbtM
AfdbuhTX8U/S8QJMtkMRB2N/aAG8wPUVB5MP+jC/14zBeLu7OYBK5JtowXsb8fwkPI6uw1Q6WWSn
5pdQcveSB8kcN6NjbPeLW838m3jpcjrG3hOUo6kDQc6zs6/ZbYy6SkW2IUPPgy5uPW0zdPJXKaz9
INRO2IsvBxjlQfDPwKu/w1jpvRDAbBN3cpAavXV46wAolhi6LmiJsff1rTxJ4S1UvilOxmkOMc9B
pHDSNoh2bJRrmIeVOVeTne6zoFtREaYRwYsIe4TOo1XStVLiSoHF2GItKQlKqZfRelJUgl/CVRd4
ZdUULtjCPrpksa5pcst4lr0WcuSQraYzthyycXBq94WxovH9k4R6TVmNXfVhYDpDjCUsVo5f1GuS
QJZ40ZW2WHmRxIy1xXszNiRhzUg79q5qI+QaxQpL/Y4qnYpOehwofX0YIMYa9GKFGHcnI5jgcaQB
+V5h6+iwWr2x7bML5FQTlRv40BZc5fwfPhzteKQ7Tk61XgtbjvFZ1kF/hL8zvlSeqPP2RjXJ2VRn
5J3QJOJAB6421aMLIZjCFxERFI9Snk+ScLM5Jow1cWzZPdd6z1cg6Om9jdsn2H61jgmdDmIz3+fv
qAfn/Ni7z07vX6cPRAJdCajTRSjFJr+1etorpV3rGZBFE2POi4z/wmIL5VWioTIwjLhgd7MLfbEP
ZNSqEC8Qeo0MMvpfa3o4EW5kge+boSJD+9plrP0w6hnIrWziBnoryrzncuG3ut5LU2YVVTDxmE/E
uf/wo8tBmBdWXC40ZTni4DQUNH9CvmyGElq7A7FXi5mYjQquDS0F97uZFIMhlw82P+9QIeo7dvLV
mjrSc3EQJ4R17NUltfL5CtNCX49O3oBijk0pD9agr188W9ujbzeV7LHC7IuggF9CxSBRl+yNnBbt
Owt5T9Yjnb0P00cyeg+T1sMnruJPBwZUkK71Gc/MNFNobjG1NKqz5/V5/hSIkreXpB9oC1XKNn5o
rOuj7MiNXFjlataKnT/6FQRAgB9uH7MM6duLVfwR2zYyrebUOMahlLP5UH9gaO+rUBpm6tbHecUx
WZmk9xtWRu2q/lek/gs77La9J2ebVwgt8S7zEboTg4IexyiutveN69wT7Jl6BNQ65kp9O46HcqLt
AC+2YGb517PTTiKeY/+xwF7cSEevZaPU1d0fTiiQrjp6zm7U5I9yUJxEgHsIQhH+WqrwipPOhf84
Ik9QMSSvPLt9o4t4/xh3gcWMmjK4cXQ0o2rwdhBjhVVBRvItqy+wuJCjHZerXJqHGq0bKUFI6EJj
tuoXc0NsmJ0DmVPiOO8/gPTy79aA5o/BU/xNjmaWWJGIM2tBj+CjDsTG3cuNSlojV4xTE8wzi2E9
mO9t0W2cGPAcs2GYP9as1J/5ILS94zwOGRkpL5MN05ifxR8d7osXW2MbW1ZYJbtO+H5+O93MCpir
8+3+CdbT6umYMrcUbQFMvinI+EXjhksBbgo12+1q5fCYfIHdSRN1XKdobOA81JaWCU0w+o+fpyrk
7KbKX91UByz9zf3Ych499lB4KpKXE12xjQTuP+UHyPxDveZDt8DxHHQ1W/WLiLxp+mdjKPInBPFd
S4Bsrpq5Qx5rgQQAVftB8hmCcbHVNCUJa9LOXabaYHBPP+360jLxtnKrKdon9cicT2Z0VFF6QMjJ
k/jUPmgHPS9jrM9Xl6V0Xhnn7pShYqijsB0XKNxg9b8NsvDQ6aMZbolRCveQuIAFBNsxD86ntlBq
C1KsL5VvVT0DebeDXo2/3FMWMeaGWLUiT+vocVj5WSIZXlgNxzQ7Y8WOFVBQ5tT8hk2+luT5U7A5
QsEJrATfgCNvuojlttWoaMBb1fI2/VffBlFiDcL4/YQFnH7iaiCUyrF1nYgTrIkFngoppMnvR7o3
hquddHKzHiyjv1qre56KA334cr4cP10ziWQcH6JeNLpqLD0cUSUmZOHUhaZTUN183XFYS3/2L/lq
zqLniyRPRK+x4dSMkfxcWvNGokH1TZczmjqA4/U48q+Nt+DtfhSqoQQsqOgn9Mv5GuRMsJ3/1DIf
1/UHI4M3YA0kEZJgMn5AkbiiU4AQkS//sgNlzHq8jpT7VocnY2lGx/BNxcz4ZlINyye25knSE77r
JrrQcdTVTepM+VxdApoL3ZTvVZ5vly1RN7c5qKtMDqa5AEsI/nYGr6yWk++Wv6fq4kImpEVBmk/k
1m/ZCk2IcpkkdG+JxDttw747w4H9D2jE5w9TsMdHhMHvjcJ3PybWyIVbT2na4NOnI5SjQTWCaLTe
NZ4J2jF2S/5Mh2FCcKcoo6RSciY3uB8gdTCODapJELKmAULBbAsh3Mwi8olyXEDTbpJn0/PQg4hi
MvPz3C5ZNRCGcv6YsHqUqoIic9/n6CqCaBgGqZ9N5gb3o1BY7XTNPBK0yFAbebyxkS9ILhJvw+Sn
1wc4SGYLRpjjGHgLdJr6ZL6AmfIg07qpoelW62AHWVe8Y5fYpz+4NxLm+aGdomq/VYPaHy3Ha1cg
Xmq9IS0XKsuoMyX6CA0hWqtRxQ9a6LpdROmsbWVdrbLxwOGYJ7GlCZwhKgwP4XweBHWWSitxJkg+
Zzp57x+KOfQMQAgxgKq8/xzGlPGSO0qx7slU5MJD0LgJDMM/DSARb6YzaoEd3gAPYCSUBJQH7epB
S3oYYC9yJtbQxbtuDJrpxkkRjMLKlt5mRlqhzeLs62d+Z3DFjM4vcLKXb3f2pq1aXfKH0OFXv5NP
Yothu8NGiUbkK3Sv/kIrzbdopX7DSdKaY8/38e1pM/etAZ7RGTom5D98jp+4iW2X/YmzdB8SD0Na
c3wOMlQMJWQc0Z3DViJNba5OlosauKGVCqd+Rl+rJBRNZmkcnrhFWmjPhJSFZ2ntP36HjkduCg+e
6Z0TTDXd6zicwyW3oAR4KQRWzTSSIXb/hbn77UiJqprDbkWhIQh7xWc5n4hQNbV+j3hAwhR4rAsG
KjTAhCOjHfYqWI8DIFR8CwYp+iVa3uU51F2m6yG2S2TZdt6vqhvWcMUZfIOg4f7g2ItVg2UCLA9+
oq0XH2aHpYIqwrXIZlBORiOzG2jqYPI0/ioYWFqslE1OOs5dMmznia6Keg578MpttkkCbye1cMCe
9sqGSk8N9VsIqtkA3O99dwYVIt4XLp7CMPXtjbvdqh3zJc6nfgMOxkbGZZ1PveLx/9LZiu+Nhot0
lqGle7YwB3CXNBsWyGTNCmmFJ7TdDce//KUt4F0dKCAMElkUWqywt8g++Bmtzg3cdckX43uByopu
OgcZf15/+dg1kE3zes1JeROziz2qH7Psym4y5iNv3KwPGPfzOL9YzSts775NxRzu/zJVWHPIoiSe
Mz0jCUGNFa1vmxmJ9xZVGFJiNoCi1xZC4b+kEm1tUXajho32lJ7FuSZIaIx4ColotwXdmv04c5pO
EI7I1xFFZOUhKb3cjs8tj0eNgwleSVxFasm7rXyPg5mDpSVhdZJ417M2ea5N3Kjfqbbo48fML8wu
ZH/jtm7XZXemsCrubeccDI5WltIdDqlFOuE1GUbAqQobCLsQors12m96yez6ga5IQTVwd+D/yPVT
n3mjaQTND7F6rHO3ckq/CQGqTCxjKAXkEsX4kx6mh6ca0H951MhQhlGGam5PLmrOf5lR4OQcUrj2
u9crHKi9PzrjzI0F9N7ckVb3m/VJ8tUU/19z/8T3nRb6YDPiH0BUOMt1YdnGWp6g/ET+KONdwFTd
PVX5I7eWHEcVlVTxIZleJJWjvVTLq7VHdIgA5iJRDgyPLTQZJ6XVi/YcE65G7IhF137ZogjHnsU6
H25KaZfq0oEQd+VRkEvZT7w6Nq7HNfnig5Q53gUJ5cKz8O6wEttg+gzbzMtwbfdLMk4PFlDdyfy+
p8RSj5NKItURA6WVju6ly+4RDerK7yYrv1pNxaB4vQdsQ8+pr0uQq2f/CoHfxjUfHnWjUREbkEEy
TPx6kUQzSrFPul94YZM6HmKKHsI3lzoQoAmcmSJysvCfUdHCpo5np5POXJ9apviRlh+cg9L0AriT
3JBtYhJf/Yij/xjF7QSSk3OPRpkOvuQMcnBkZqXx641sr3L0nZd7rOlEG2kEvG2ijM1ZhGnl5VRm
b8OcuU1bvytHaGUGhNisyugD7nXjl4AcVEezXNw3kbtui+yOenNJxOUS+cOhdoVh1pguvbB5lF8u
ZU/dJZXDhm4O7sn8RaDQ7qJGW78dM11jX76gqj6WLfa0Bbc4Tpo2hhKqjhlbKvPTQm97/4gn/W+x
a5k/G+GAcN/Em9A27m6LuMbiyCRHXqUpbsMfv28RYPtzvr2xeXQ0JvtjfzR+a7AYNy2+SFy5UWrH
gAtD8GugOf1gPZWjiIhI9rijjY0fenuXdFBrHqivutuYgjETnjj95zuZhIgnDPWtaU0lV0uNMxEW
LbofTIPMlxyqt4ryWRI7YGSdWZNdqfXGNnnn0oxEjI+4ncJNy0ZgkMuHdubzFGTE6J0WZ19MSuX+
yI6CptS5SpJEpmsrHmCvP6n0jsrf1oVbHQ3rJo3EUC/pDmdV67iSwdpXJk8p2iGhs0MjBd/zjlpD
0I7xu/ubLc3XkcrSNkEWA+58yTwCmvhX/057/qx3e776gjbn0eDr1Glu0qU5DHXhWt4QgkwrBlW0
J1Fohi/gBo5XRolhk1xXkewgf6TEmzW5EVDGG33vmm+WNFG+mpALYGiJbdEOeicX+xDBdG/WSv/y
zuy74/DOdwlRshHUKSxAdGKtRuqiDnOIJNjDfzUvU2rpKczDmz8OtJ4b5h8thT0jyIg4t2+muZxu
tk7Ck4anXDO9RchCW60Ld8aJHpos4pLwLvphU8EI0lZmpAbhvPZOnOuXZ84nDOiatFf89H4zqFtz
v5oVosNfZsB0VhgBiZ9tJPgYHu4XiQrDIiujG4ljD+hVAarj6iM9trzOqo3cQZBz3CY1p8QrMoJl
mqJvELI2Opurn/CyqpVzth/ezbqZjyS3iTlSUhmzKXwlQG5B/YrCAqVEX/qQLtQk6dl/mrkziuzL
ENhgXXY6KPWDUWLnSlZH5Tld85JPiL+16Y41Fx67NfZ23HGIOnVipgZ2GpAPiaunN3ezeXW07h8L
KgraJVzcccpnX7FCAKctv0351yQw3AXS+y+sbK1DAhnPBPdfgWv2Y+qxTXDchqLcNNclX2q1CFEB
cCl7RjyZwkrcRfZoA5ZuCKmSSDHiOOYUnWQZLBoI0Q2IPYbn12mmM2Ql68iafWXQC1StK8HvUEgQ
RfbGvXpwu1v1jotS8/x2Paf4+WE8ykDvf2B1bdDx1noYEcJ13ED+vYbLqgz+TQw2wFkaU8DFeTOB
HIcWPttT1gHGoADCzsIe+OaI+XvcENRATh02RRM753sFjGUwYRd2dksYCpNVtxYNs4IU1ExZbM9O
JfTF2KY0DVd25jHzmhgxheKyYR0Bu8/7w/IX13Lc5Y/mwg8pAS47mnfUQQcPWIEGWbxs0/vv/sdV
ovHO/MF8EZWM/xi+aTTHzFIZFBra7JUyOoe7TIAnIsg9juUC0pvbFOT9J/XB6vP05zksghAzwVJE
DqcVz3Mtd1wuZWENQceGIdqmWOwYyFzLe58L2PTv/Mnia9fEV1k1sGdEfZAc5IjBCjwRAQB9MB7j
/vSzD14cqZZJaXDQZgcLDvud7+xeKOBj7bH2kcx9zNBM2Yd0f2nNlckz5dzmac2N0/JyFJyn3vNA
gJ7E2jmC44noXUWmDRtbcHBECjcFBkuGqlk/mX/pW9av/l7e4I1G8pX0lT38soLsTs4dQUzo9Dj7
a3K88GD3xy01dB5qXpSWU07XHlfiKu+yicfJAord4XeFPlYtqyFzHjf06oOGN3YpCyRgYeQVyghN
M1k0Kd4bXLGpkWBTFTIollA+VXGgzbbBVeVRAECM30+N48wvY8C6Ea/0itsSYoFuyElhiI17E1SG
dCdIV/4XpLfpYKU9V1XSD70EWbpwLJcg/hZN2Y+G4bWBPttMaQS7F74XTI7eEVc3ok/fRINUhlN6
iGsphGMRQzlRiBaKCpPG+60zeAti7xx7ObO58LlvXMJqFl8yBLr2XYsKdw/4w+tZKcsu723n28Rm
NugSssyHG08pWX4YgbLNL8htM8VAqn8Hd5I8K7TrpeZGJS/3LOdoktKB1udTM5TZAWV/EVT6bdTz
znt02cdh/Tq/0Fk4uQUPT1bSNg8U2KoVbdu8BdGH1GoJdiLmgcNzZgGSUrvlfMaNPfLDFQ2SikZ5
4UU+q1bQndxQ3qJUiHiiglyDQySYiPxAkTKawwGMknq38ZF4bk7pD7XkdbekMmap2FSN6xjvcXPX
HdYutcdupeusdYZnF3DgRuCj4zp+DbIYeTvyHMPBY3gvcgayYzo+55f7i+qTVRlvoxuXF7OGDJNg
tuR4GfpcL1M3I9WZNRSLeF+7LhUMwy3N2fiXyA1SxlooqLFuIKVMgyPJn/dO9Oi8jdPGA3Q/JQ7Y
0RTzbBnRP8W5OCCnRIyAqOM3k+BB7DxEAY/KNCd6AyBy8B1dyoykC5Grc5cHmHxH5Ax29/n80mm/
JOUNm1klFd4SoSKUCGTVP4mr/NFmdyRB7mY1CwoftZRCcCmlrHqZtW+l06MPiYEkediXpv4d+bOD
CRrBBOOwIiuB343iGLZLlkiTEYnYUOe7bSVyY2lav8sXDIpZ32KbWciAq/bkfueL6B2ebTPeeuX6
qyNsVKR3w31UlwmNLOncgKUpwxV5pZYokOjcJzx+GpVIXQCEiIRsby/xNl2Kv4wQHKQfhjhYQhFK
GaMv2OhRxprPWVlEyv4idkXOWIZKNAvIpTA01LdXsIrmeoaRKnqST6bKirueEcvA0AY07dr73Fyd
X3SRuU4MMy5gZwJxP64CqIx6myCpTxGxnFI1OeYW/P/Mw2KE8OImtCZ1QtbHe7iRkg5qFAYBsi2m
jaydcQwpo4xEvmKJk8kGMsc8mY47aejrEmZxlFONZ+CXmemt7b4RkkmWjOBCd0AlFaqmkQqmMmMs
5jJKKP+k59CcpCe7wPfS4c73TY67V7wkJdKUiwYD4v4djHDK2EZGmRkUWey8o952kLRqq+GUoT/+
xJcbacMthFf8olTr0DJvBPWG8i8U/UJNYp3WfPm9nWvgsuGyTlefKLcryTsuJlE2MU19QfHUyNbC
tagKeREHfihLTvpxPT6yisBpktuHXYoK2ZakwNRWL7u+aHO0418gRqLL5uD/fAKF5YL7LfduOKVc
1jnviZS+Buc9COOz2CJCuztINE3/AUlqvv0/6Zn2IW+LckhGa+5a5zqUgKYAJcHsrEjSnLEQMuYk
t0xrQ5h5q1KgGFOJQ8kCKvc92vfloO+Pq7BJVlF5AtkQ9arD+8uhaMQoCZ3dPxoFcELyoX3flgVB
+scmmH4FwZ6KSpdYYeiES5zQMtVTGFtqDvRbKdVhwjpxpTmi9jq6hDQXVtlXfujF6PYnBh6IVGLT
dq9eetSlKzXuuS6HPA4Cdn80w4yi/H9nssMgQDJ9yKuzzSTL2I7bNflm5IT0SrBCVj6W3Kd+7EjM
xPpHu0xSo6B1UyU2Row6AeHUT4fEnEdC4AVMiGpFbWymkiDz/91GHy6p98fvQ1/uTlfOc8zLQd70
Wo5fWLOauZwEL6VvI1BX72nxbLDWJE0BWpu7owVtCrViaK5s3iqxAfS+YpnlIgfQYruzbsoF3j1E
SFDD1VAL7CGORT8mWRIhOy5IbcurG0RU/hgjtT2aCFQvMcjF36uuHGVnFInX0F+QA5YEGLSxztAg
bLOJp7jQVXhNVpQZQoedlXPx6kp3ZT9t577I0q2GaBviWiofEXkKq58GJ9UZp9tuA8cMzZp7135l
1xRNKV/YCWrcMI4btbqzP9xLFm/7i2LG2vVuBoAe5VYiWEQ18ltLfHXjd+63lmszTKJtnwOtioVs
6qSmdnMiQDRQBeOXvivBbdDYrgvl1zdMHx5DzcMFaZakdwzfZn7CGruv90PT2a2iErnupTSjgWTP
vbbgztYMOiWMq1jhL4vhgn2f8A5TffE55NBLRmIDy9EjOoXZ44+6jM+dLJyr+tIHeCWW4/bKgr9I
oXQMEBKES8R5MkCZBPSYbgmlM63rTM/iCgQWpt8sCWpLDovgciYderflU3d/mzSZByaDCX7r7Ej3
ZBXi/bMc1j2hC+fgcckpdoALEm+uFMxAO7B5wIA5COdqikRrRXVDY/zhVkh0NA5rVKkMAC6Jm30p
QBgtVxxr940PCVlD6kTqXXfByVUTNbIou/Ick7Tfu6Q/E9kXBeUTNbb1KyfXhvcgakSx5JyEnD/T
MBBoHAqP5kuXATPg9NTACkqB+8Do6/JVKQ1X6KgPhQ3SV2k8VZ6u48f6TVLosm4QkWXZUFaT/kKM
DKuizRc9dZZX0QOdMq25N79ESqQGO6/DvZtnD8LdcQO/XcpzQyvoxDMCYuNJkXB//D8J5h8AVhes
bQQPdSeaxZavk2e454E/f7Uq+YhGlJzeODqCrZRTv1T35PTUJ28Wa3IR45Bl3d06kwEhzNqiMmdc
uG0RQc9DClsBKZWi0ylUJ6s6YzguLoMu9zwWmF0bux2VgVKaAkUoUpRerSM4D5n7kVz3ZWVWa8Li
KtFE6/fHzl9fslHcjCKhXGD9A1nuRAGI6DHToPoLrAfF9U/jbHoUO4g1ypZIsUvmHobDjy42xEOB
vBu6aUQWjtCHHliQuEGsCNUaTlpp2KtKkyRtcyf4CsOE0PTNAi0+JskfL9sej/Zhv4Yrb7Z8Z8F0
s3G+V/OuoS4/0t15beMe1e+l3NCmMqqxMXM04eW8t/pEaZn5CXXqL9W3ik9cowu1MMJ1tFzoIBv+
ksOSYlnH7Aqz2pWxcAsYRKYi6j+feQ5yViA3yxgKf5BaM2SZFcgKGhCUc1lPV75vrCAjOY6lTpap
mAyzIZ5khZ3bWLVZE4Ztwv0Io/97aQtnqE34ZRrSPhpluU/F4fSSYZA2NF+HjmVVgVNJKNHyUiVx
Dxp+8CBwokt/605mp9qpNT9sRkqGKtaAJb2Se3b/Pw3Kkabl7LzQhbkP5F/tsI31+wdNsoHXNcZH
cpSl0CtQ30LOgchfnDFGI7TDYzTpEHrWO4eme1DJl2dE6KMQoAiMHwItLWv0FUhkis9HHJsCt57P
gVDkIKKCROWEAMjZckXl5PV24/Z7uALPcpD9jvVEO8jdojNMRzAbLeWua03PLBnsVgNYLoS7MeyW
QXdVTB8HiIOvp42HMBqV4+aspouSiaJGi1AtHORrYVwS3uSB1bz5tWaqsuVtdGs3muLzBsffnB4Q
A5jfAko/l3Wl2qEE+91wuY6IuExqrlh6TDK7bm6ndV2EyHb1IrYd/YiCj2bgiex4uqPtb7CwqcGn
zjLSyHHkjhV43xERuhkgRZ5x7QJ0kLySSaeIMO4OPZpDGRVZQN/axVAwv8u6Mr3GmxjfMdzQlM83
gZ3UnBmygDNkciZ+5mVaQbyICPOdcUbjSeQmVdP/g+/vLO3y10wmNhUFZyGLYUEF9Yzx3LHvQt1g
XsgV7iv5xTVEFwGAe0HJpCT/mtVO25i9GR3San57HTpbbo3+Ad6ySZoRLiSftd8OVKb1HkWA04Ki
JtOc30eA3fkulE9YRnTSiFE4JGSUaMUANJxoV7sTP6vwDCMOBM8JZGhuUtVDtQfxgJ0yfTmAxUDd
eapgcNjMRZAD/jfGb3gXke/rUEdW2O6vjqXExSBlilA2UJ6WEkkXH0LOFJjn3J8ikEatlgCLl7BY
wE8zlMt+kKbtwyXUCfFbvwxRwEDQMbiMV7U4Hi9PB1l+/pjIZ+twdjNI4C+EQBkBXvwJrKaAiAU6
w5CoMAlPtTHYeQQQKw0BuR+NpnWphZZvni6PnD9osdmTvji/+tWOGEdT+AE+ggZ7FmutqKFf6bQC
YFz/QLVWs1dEoeaupqW6zHaiZHqxPTHz2yERmwso8l6cT6MFnWPrqriGTcFgBcuaL9/Gn6FahtY0
Vm6ARitdLqZCbZ1ycSo2ZBO24XQSvIZh/9KpKxou1ifeMCAWGlW9Nes7xX4tfQrKT/Ls2D0Lak6i
DeNIyojXPdUdlws9uXLIvVx6chIfIeismU8r3MqggT0QRv32AQO2Gy1jpQmUyJzGIZHohFHwxtEL
yhWvVXtQjuBLV2RjnKgzwgEqc0H2udhjpbb78PdO56nOCA7tiseLdqnGEZ8sX3WzzJPgWSnG+xmh
VSQt6WrRGcCYoSmhgEqoXCi/2l4JmDfkyPSlWqqZncMxNusrhpIhXQ4DT5txLd+N9ZuJXdELwBz+
8XGO6rwOwqLCQsLQF9bnSh4Q528auaG8/ekb6ghC08oJbREXE0y0NzsYOWDIaMJReHmRijModzIe
tyi3WTYQFzLy3A+JKxKiAK3WDe7EoJmGbBm9rJUu+cDErc/3IfAUQEgVC9Pg+2VNRlMw6sTJPBAv
LHEdlUJwTBO+mCF/I0fp6Rn8rpSvG5uNKaMaa7ntWpIcr48+8He0P2mBkX9XiWhUoUMw9x2V2EkD
i94uuhl1mra+ufNjeKcV24tEqsOeLeNmdaSjIU3X0B2DiWtgOoqdhnztdbZlwSn1NoTzIBjjKePl
UwLv4M1i41UCTPFnC2OJFFOmZqn96QbSRP1fLq88IohkaxdB54YnjXP5BiyfRArTTvcfPcG2yggM
zM079V3mUJhzvbLw58dpTneIVrC7jQ6PU9hESFBR1sEDNSFNoWfUSl6VWjyzsJBa3iCWvBLpadGg
3RHTF6w+fU56skCsAANU354ZYId06W4WwwOp5N36+/5CvAKyaU0K4QQueagtn9y1bQZGrxogiOE+
SJX/8AU1VxI63s8BP+DBjsAnpQtS+nnUtJhmXvMkQdjDZUmW5U1Z5W4EthBUpMst5ysqE1A2i7BT
IhgVt++9RJbDejkbYtOExoTzgX7PqFkUsMrVz11xHII/SYEYafGR0OaAzDK5whrJQ7KPIcukKqVd
2qNC3U+O/uPb7rSEqVfGz2SaN0W7I2pbVXbnUuFvsEqwoK2x3qKXO+GmljDQ0AOhXO28AR4CLXxU
IdP07wM9rF0zHfVPGh1qUWlCGV+3ZnhAT6pbWMjAO7kviDLk5BQYVJBsIZHgAFUvyaMU8sGmCbLb
oMr/nKPXyobUfYJ9im3NDcadmlUGOVBtLBBpnob6YmnmPKLx/gxVadRBIarLsaC9MCjtld76N2Bq
eAv04NljvbyigoKzSixYgWbeAe1WApPYm3mrlGsoqHRZPZaTYOPJint6GGxqhT1WnoPi/ZR6wuh8
9WgGouJ5+ZtTfYYXdQlz9nmdOHvjQvwWCABky0B1Au0v+YENfX2zH/k47kJe1arzBEQxiQfQRAAU
gi1V8TiMVn+4rguhaiOXGwdg5gLs+8Z/Req3oh1Bqx8OPDVKHYZkej12Mbj+8/mySQUg0RHsv2x/
E8tnbdMj9ffOfPkkp2t+BafTfrWljN0ugs9GY+xMYNernBTmgm3buTB/ekihPnFAf0bxcW0C2C1F
Z4geKJizYiUQxpyu+h8loD2drpzXP9LdDn8wdNK2xJMQp6ZU2guZ5mfOUePdBAVliSDlkEqzq7Iu
lqzyE3cEaGQbvICd35cFxn6o0Zfw6uc5ra6WXVd28atc+nshI1t6I53NX2ETKTz/VxQ67s/pdKLF
C+dMO8k3LRttt5hQFbKAs3q5foWx4l7XoZIxlkDFuKGcwLWIKHxUGUE4bq7XlC+nR5iFkWuQDxLx
5Z7dkHmWfNW+JDkhWkWCvWj1vetuGR+qx/AKacAdVPUh/TRUoq0Tejgg7NVgNWTc/ChaGG+y8v/G
SJtnJkxssX/7VKxh41pRRgqmraxPAY6vSYWwWDE+einz9C5yxxTCH7vBlKWt0nwQmpJhIojkyaXS
MNHMjAhDXVoaeqy/Jfs3oIOoGippS0IhSpGRYPgOkCyyKylZcAQ6QU5N5+MzJZaxsEowt1v+2P5V
RSOW40chEMIfz49YwqNcpXGGtiDBfTB9+mXcAkztBONffxBPDB9IMryqL6S9b2S5qBAqpVX8AYD+
88RE3dQwgsiTBceq/s4oiVe7dnqMtny+nflNAI65CCCf6roCc3MlJx5WaeMyQ1+/MRR48I6tNfp/
qojWrSLbu+Er8xnJ0fkUQxds/nS55buJrZh1a8E6Yw8kiw1JRLbVVQ7OpKRxRpjbMYiiZ0u9BOns
ELIFL1V5Qv0bYP+6IX5+fTUnBXYm8hHL0DXWRKbCQbsGL4mc7vuFYk0sDY7pmtOaQ5vwyUxbqKUC
e1xVCs/zTdzjJTrdHCUiBBq2+CZlL3yy3BZ+T/4yIIrQPwWLGPXJ8XmTIlDd9PIjb5jkI+kNaQ6q
hEqev90gwH9gKGFRoFCKQeu7CWDUMatuU9YzZkzH8XKSHv5z3nhgK6qBIZjQMc35NALOtj33iYI/
p/w7vT+Q7n5jBaJtqRdE/x17kTjLHQ3Md+zBySlACklRkUrY3jpmFPu5X2r4TOtjAIwJx5d6htsk
0ZFV770hvCYtNGH/HfdrUiFw7OyeDzIaPF0kO6Cnj5lhN7YUy1KP1sTOt0xgpGYTthhhqzuGofcF
VYeT1Dzvh6T/d+ZnfDiEmPL0+pDfyk1H+64u3CqklsM8Tw6WMqYhxidl+bV5wUN+nvo3H7NHxu/5
dH4tjHNYtEwgz90+p5doO0vnvUUQA52INnQmo1/bdEoPwq8c0r0PHfHKmPqTcQpFNrpaqunuicHs
YE6i1fnBz5wwrKo5CNmtf5++E+2n1p5xdKdXuutf85WUksvENNM/ulOQCkJKvPtlb1lXY08Pkb6P
Y7nMQeh7pgECaXQAf7hNLHngHe8luLHzrjNHL4d+eD3qDqWQmM99TOyqQDLhIqlPCtQLzqdIFjU+
L4cjVsIOPWXIdkGwMlOYupdgBaB6ewxSm5Gv02WDagnI7h21rE/nik5TtnT1MJnbPvaEGEstMkWg
e1IhnQcTmsvFSV56cIhhE5UC2sjSp3kaJ/3MjK8+mbGYA+H6qx5woIf1dGh18n5G+229yCMHD/4d
dPkhfruY2uiGuH0dWyUO6A1PH+LaKBCuF1AlU0wtTm4jbCeGVm4ouZJtGEPLu4sdXu/AsDIu9EbZ
F7c0WB7rPAyJEY+K2Scy4oAIZ4sdsitIQVYDk029ehmjKg9+vOPrXn2yUOseU+8f2JwaYfRryJYs
8urLUZzsHeCa6oj/w+MWRhIESxrS6EKUdHtiwNCvTD8rHD54WhCn637g1b9DN/HMX3QaCI6BmWIt
uojNbZN+I6wdUIPI6DELy5OkPlKNoeoYEvM0J/mJMAIi70W5J+pWnvWNqwu2H1CQm9o6neflVHwy
ZqgXm/9J5InArFVOQZkMpU28QYdcJteVDAvgWGLjv0SJaB4i7PCHHYpW5pPGMr8ehz0BSpL1VI/I
Nji33FkQWT6i1QRPmjldvSLu67HXqFzUV7nc3DnMv3QJ7GiOCZU1J/KLMbXH/TMXCkh5ittGsbGT
TN4BU/Ss+4QMLCYEMV03B04QdjAyUt91dxmplWBEaAp0UlcUalFFSKeMtIQ5lrEyZQxOpAENjr3G
WPif8mRAdbErosyL0AotPKX4T9yhBaxyOWJQ0/fZEkvXaYTJB0NOCcDEMqz8CdqCjLMF2HF7E0hU
e1C4TdZG8OUzyQH79us1O/lw282oZFqKWhnAXg3nGJNnrwvmPs9wQltdTcnwTEPuppUQXamYvWXN
qvU1KayVLsPWEFG52p4IOsCcf8dID0gMct+Dt2hMLBsNmXfmW7oVdQWlwVreO7dSmKI3ep18DU4S
7XCeWBZwAJNfyVXgDY6PzhWM5IU8fxIxfGspoyY9q9UkqyuAs0jlqQr1AzfdhzqxIXlYPAOkuGZo
Ys/kOiXk70kYerYbG1O4v/40HNEyG3x1KjtR827REhaLSqHLZzFrOmgN4mIfaKdkNFn3bpS1mufG
vROAlgXguUrtfRqb0Z3HuoaQLAbkYJbKjmcIZkoacKxLDPwd2K09CmKfgKStr3YJVFncqWqlYh8i
4pjgKaCVbFB4Mt6MlSLfRv50zMxr5uNpZGcaeIme1GxB4KSviuGnocmH6Tm37NUn74BAVcw3CuJp
BR40/MTD0c7ydkkoj3k0QF76W77GxlTp32gAjjVD9ZCIqYkmTHTkdqRf/S5qPjsPLv7DuTMiaqVr
kvaHSq5Zehia4FGnNxARPJFMz8Yw8xV63YzGfbMFFKt3c7nMLRPhlpzf4qqJ1zaLbWAbOr3ap0A/
4Dc2AMdopf/3U/H9rr90XMVVOZOSffHl0wOFC/oH7XF3tQ9wyWWiIeMbgjZNLJhJNpvX29Utl0Sx
yUlIY3JO+sT56ecFMnCHDtnXZnxCaM30PdPxxNk7OGztdh50S3EEVnmVMOC6b50r6LC1cSUcXLwN
6rom7o8iPh9usH4lP8bFai0SnYh9fNk7pIoSm85FSsdhnxX3xgmf4HbFpWGmW/miJK1EuTY7Xpfb
hMOW2dzTwXBsQDy92gVZsI9TocopJi6+h1kjakM03l6FiWCiwHXyok6bMQo+QI4lKnSWo2q/u5bh
rsNbVztbNdftNhH458wRbsp33GUL23j4BAnyj3FauYuNnZyWbfBgeQQU1xdX9dGev+lnzlhYNLr6
QSXaxrWTPeAVbf487iNkajzAk5ioAk0rYCQxO5u68c9AZIZ+dWKOYcI0KBjojahfm7spG557Qfma
h6GXnlXMonWGY06qOcsmGoSRIhGiAi4lqF5rsa1RYFGDZm+wdLv7j+6b+vVw3yEI2MKpvgPXc1Pl
M+9OgLkSNW25UhUEGStPJupUVl1GSV9GTQCofiIt2j34Rt2IJFxSUqGp7ko67KCOyD0ch8nJTlgu
MLJBWL9TjXFjU18PSwFanyazJlf2FwYrfK3KQYPuU4iwVLbdc8DfkCrp2e2wIZjbdzsBEl+K/CY9
Q0wpFXeMtstZ+KbyxIgdLy9ARnyOwRvQoaJLdvUcVpJkXx/Va1T0SL/jjAOi7ALgDxO+BBPP4UdO
dHU65/TNCG0lI2zueQutZNIfgNSJGT6UygVvSEKLh8fgWDyMb8NXdiJ7F6oP2GHwJ2Q20ZgLNWfe
Z31QNOT7R0OwGIXlysE37heivuEvlrqrUUClWsZrE39YiY+0N5UhxgpD8WeY3JccjxD7J4yfyhIj
ZzGJTCjGVd8YibWqPCScjCIt/fHnx4lCTiH50RYs4Iqz5FqPOAGK7Tv6XkUhb7nYzcG7fr7GRkNF
UfVVNRfVDEC9l1Bio49lljTVmerSCLnU9uPqe7hCLgFmDJyBGeriIrB+Isjex3Ua4PlYiRGrx1e5
h+ILBpV5aFwmR+To7qjnO9X9hmi7tK1glayhwkPDKXyXKa9FbYQp89FG6mv4rxqYO5r8ckSkq2C5
QXuiqDw4t2TAFFalWDvlibavCjGoMlTblS2sp+XiOJMmW0Tpf7fLLoyCRsyx5LbrQbY9Ol4i1nGG
EQh/7mQ7djt6GxAdfg3x0dQlMFn2+i7Ki+yT5vEfQLhI3WAdTzC348lcJVl+IN9wQavNHQQ+YqiH
bfVHsi+DgM7C0pGKPkW7JXF6p1IklixWKzTXK0tyGVIUSLrMoUBto2MvhMlCkAS+7G831zH9BT4+
i343LFpqK80m8zlQoiWgylnzf0TYAnw6S9fC9XIOnuvKWclXM/j+rOX1xyLKoXETSsC3DciuxReo
VMRGNjCYQyaWEHHAI96SYLttYJLkF+sCIay8DMqUUgYWwaRG1qEwiE/ZPHqeWinf6rWSOgnoYo6U
GDRIwByNSVIIlyjh8zgC9Mi8HfjbEod/EdZ0hOLALubOqcesEShijh1iilYOLtYYWLX/GWw5WmBE
xFF9TFGSKmf2KGkKYRoKhrU2PgyqQLz4KgqVZo03tp/8rIcJRnrHVfy2wfh/4gjiLKp/xBzdckMo
r1i7H/a2HRUCMH9guq7MoLrtiFzAYdPM61xDPBPYzH16jh35IgU3GBNmYLHhjoxfkTdA1e16cKcC
+FWmWZbjbU7DjW9GbUguvf/z1/CxMQc21880A2dnE66u0xOg0AEnKzvYI5JQDaTx4WjXnL9Pn7f3
COr5wp4sY7+DBkDp7KscXkLWk/UZUv3iUNGVqNnmw8Pe9HkN15+WzyMq6BZFvAoUr/Rz/zezGufS
kzpnoEbd/hwfEpDheS5CVuMrIe61p5bMutNM6YgKYy/99kS+9I+kdKTnwA+Sl5zqUwU3qOe9Hx5H
VRVzIlnkFIJp1cQw2Z+jO1HF5V8013VCtmv543Jad5VKEMO03Xts+0UcZafQ5d5oGCdCRPMmF8eN
u534CorOqNyNSvJgDCk8dPHJzHMAp/J/5mXPKDKVhIkCEVI8/s48m7NcJjCr9QQzikkwqAcYSGZW
RZFgpGucwUT/wB2VH+SkaX1fMRnPx0KycqGkADHYmpjbMRWZ77aYmGPcXEoqks3aGunmi//gr1qB
BkQaPW50n+B89HzI3ICSuAqNxKGEJVFt5D7Y2ygAPiXkjHAWTL31DslhtDAgHdi4KYbwJoJ4LUQF
whuxKdfSN/iZqBJ9QszDKZNbHS1iNVCR9Rzz+U3M5rHZ0Bnl6FuNuWb23azVRsgnrRt7WcOnWCyb
CCsopNDUHn5RGrOawMCo1EnHRSrm4pWEIfTpZBtxyiQYc2FAiz9/c68SfKoSQL98hoS+8rmNTKwa
plbGxPz1NZGavpq3aiaIheRkwhGn+ryINWtHdScLtFJsqk7UphJue1d+LoEs0SHL/uVxU2DsMTOQ
Ug+uDs7pJ+nYJr4MdwMU6kAoEzEuA9B65FQK7yszcBRQXpwCqASFixtQBmoAwkFbIKDYBIGMtqni
pO2fT4oT0CquP1Z+rh4xPkjaMF61pk3sSgstoqQgRUBgimY3gaUreTFpQUc8rAAxJIOfR9E4ZQJI
MEjPlYw+fIyvexx4/f7da5AQs6uZmXUPXGYxJ/eWXPsqTm8/Ksxzhpkee4hYHh2FPI2fWX+54Lfd
J/81Tp2e7F0dkbFA4sP2A6jZDtYeOVDo5OYO9AIlSSv4lPvhZgHZaQQ8gbzDSjCP1p5a83JzJ5Vb
UzlXMPkO1ltKgn5VB+t5PtMwSEDgSBlo8j39KZ6kROF214umIbeKIn+B/rH6LkA5q7rbITbsMsZM
uEg8l22sY2mUcfr9Kf094KqEOaVOXTMU0x24lYrsjp/E6kdwVaDSQBpYpJr3riWcpBsr16QHeG+Z
NH8xekM4pbmU2U8DDHNrLdu9Xwww1dCc8vWGFjs0GWjeJI/7vK7cQtA4IXtWkgn71oHtZ0RPKwfr
x8xKSMfKxSYX9F5cmORK7J2ZaCz1mA8DZz5O8dvo2ctT9ROkhOItFslZn6yjMH2eZ9OCOQTxEsjE
lj9z9OavtjCG3/iXAx09FHJzt95TYDgyp2hNXdNdTG8CuQg6li/6LFhg25WH1ZkBlGORqHyA5Hu0
3E37hh5oVwW4iLIXh+8EjG1r0rnVPH2zMuPXR5dgA4vUcXMr0JVg8NNTBmAbR5bHdJ6tHCdq+e2j
0f+9/zV7RDN3acN6JeRlDRZb0WsEHYXQw6WtxeN8ohhtF03J1t7QjZIOP8I248ydFAAuvq3IhjLs
wsiEbUUZom3adaw+UvHXGX9bPKbBEuZyo5vxI2uTFzH+NAQteGU+wMRr4Xc+aBcSjzjeQrN5Yw8k
1roadJ8dRMBB80x+aMIJSSEs2vXnEmWdbZ2Smp9osucrH/vqBxM6+zrzrxdiZZkW62ZiN+88sm9g
9McPPvjb2M/WKNQK2JusNU0H+0nfvQunTB9EykoR84qZ5haCMX10cg1I6OH5QosUI/OsGhspYjjN
6TOSI7rLvmFpdjtJn7EA2JjzC3RcqJ21C8emUIf1taFPXWFEaf9KExJuPK2O7gt8EcF7yeybgm8s
4UsWPmVDv4FA3ZQwQfMaH1hUEm64gW9Iue41B6UcB2Op7ZlKlauip76A6pVaEXgLbvuLcB4SswDX
CcRPsSZFg6tzH2e6MNoVEio+RWlSxt+AUDA5ZUh2DCtHwwJRmP5Kmoz6pcf6H/5Exsc5bIEiRaVp
SJnoDkUjB1Ys7vtJEwG8XTHHDJhTG1QOL/4Z2+q6fyIxu/Lfa+Wi30d9gqydlmGnddLTOZ+DfKof
fuU+mki7sWyIzN4Wm8+L4Fc4dIHTMQwp8LBKAf4Zn2nRlJRphfe7NJ01v+8lX+ctNw1A+97P5l9/
uZEPGGfTibm0nliz7mknkcUgNVOMCknUiV4KGIJjxJsV5Tijq2tSGrmaUmgRL703lHQmlnFu0eUW
QbvREzFl2rI/D/l6jMXXbKHdkiYIvutjJqFdNulogrRJfRAT05D01t44veBDFpqAUnn7IUcUkHaQ
JSxsLiM7+Do6yBdDnOXY5EqExbXteOtvvptd9WHnZAxiOUhKrwMDUJhXONz6ZF9UEPpD8p4OLvpr
cnODbJIWdg9bcN6T8t9VzuDxToEwMkTO62W8qCq5IOrD5w/M4AepuyGIkToFho/7sPMPFPPB4zkP
kwL+RwO6F0bXlaOT6LMuXbyzW2ZvIF8+olVPL9zs7KMbTazrAYTwSIgyxdyElcrQ0lHbl0AfX6Xm
oby5+Ghxcm2CfPpcY/q3gGi0NP5z7Av77gxNOCet5D42iEIwGguXlTPS8iO9BWmTnjmLseViIoV0
VYfCY4hsoZGp8IYIXE+eIfiAtTZbiKPUJIEjL4ackUYFP9tTU52B9Xd0LVMVumQr/hoWfdQaoVO1
0uWLFBvmaU+NGQIhLHMH2wY4BpqbWbNO9S5F8EBkNyGuXf3/Q5gnZfl/Ip1AB/zkW6Mexo/PiNrD
l9HmLOtV6t9fxhlJwU3hWNMi2cMPJWdl+39vAk6WxeVSYs6HO5HHrkkWwMuW0QtRBTAeNJIvzg6N
grXZFYcJuoDZdldcCzN72X3iGz2Gi5X//ppcShYkl80nW0OWxyyBMpLKSihQjdSEiNzF4aWk621P
VnEKfptI95jFnVbukmmBxBk6l42/Xijm/zt2Kva7QsavAJBS0tXV+ZmsCAfeqcEarw6QyuRH1RGB
f69hL2xxM7pdggycW7Vjkm6r/B2bxeN2JLm2488g4FAfm4yYecXWWANkXYyTwTor81JY3KE0cTin
xbO6SQPoD2J/57SOvWTlhfJTAneUD884Xgwb58QfurGlcJqIiOCpTQENvtIihn5dMTnM3EiraK11
b7kvPkI5m75bdvsrHanq2ANrmwJlYwyCXkSF7XKOAmDaX4wXfyCkAKwT8Ej9w1tHp/a60AC0GWuL
Yc8qjL/5BJELbu9+FXPPQ5WPk+7hLYuvrIn/K+eJoAsiRf1dowAu/vPPwsmUi2mz3LrcAP0SgWOZ
VMras5Ro9mjaaPV8+00sw5u/6Ou9xvGWKc3HnJkVGVGqRd5T3vmN9I18rpKAyT6a5smCF/7I6XAK
I+EOosoiOZvY3TrGmVHmScef2++3z/9xUMtIwXIgZ9FkUYl9kbaH/TocxLIBXKRhKEXMuokKHCEk
hiGgTJmJ9/E11erItBuc7Qjyuns6cTP7N79Jf/GlilWisMR61bojRi2goQ+d4fDNQkUIMWSOSSTe
tBh4/CwOYQ2fhz86bk2ZeUJVcZeEa87vgVyjDvfuy7VKGSnEUc29Tf9FzwNxs5JOXH8Wzs/2w35/
pPn2ITE44nU8J10PDbCvuKbUtyBmXbw3TETeV9b6YvwdXshpKxJ6Zv88DXS/T0VYrySIrQ+xEXyC
5qoa9mEXdrd6w1DeNjBIEUUGRZULLq2A03zoVlFHsfrJQV8SIbIB3imEayNmmlcy6v/vYN85+8t7
az5Azhr/ckLK06NYOc9vKjMLIh7k99M6BXj1fGy7rlOc+HYsdXV/pvd39xqYlNLsNdsxpLZd7kV/
3NXtZZzlFP805acYXeSTOrmEAu4AYR2ElSBzdWCjXPDK8R6FiVUuTJGHNi1p48SGUudAguJTt6Be
0be5HT6PeEkwZUd2ju9Wi/UrtPEeSjTrPRoqbHqqnWeXjjA7OblSEHEfipPj4V+UluDBijkqbOSH
wCEDYGiE7qw02Yh/XHedSTTaNrFLVTDIUfA4po2/DNKpZ+2F95HyySmPem5VoEOyKoSHBsC9Ulfw
Ukk53rF//Qcg07KdFgOw+3C58vMEBuKqozXVSH5CpAwr1oxl0BqZ2Pkio9uGkNNJO/Igkahic2L4
TO/sW0ZFQZ5zRRjOhk95O06W00fSN3FNYEDZy/K64WvSXp6a5BAZF/3D4eEHcNA5PPOhymjwLtWy
JqUrKwkVHA8tELFQujAqWzslk4JRYXz+krPttomCO3ZOjvNFD0pH8lj4/EFB4bzLUlvOkI4W5z0+
EjQep0Iymx5aukx68jesjBtNuCpPvENrXHBh4V/lbQBoHenFK867NHQWe3/L37pz14dvqfeyNbps
ws46DPFGJfW1/90Vy2XEbCUPGUmfTrsQAb9P6uGyh70JW5oyOQyFnTutMcPtlsxZzT76451BXfTg
KnKC1N8Z3EBnhljd7VzbbJCfECI4aTPRKATtkw+2NxQjvN2aTf+vDLjLA/uwlXj3Rk2JaP4R41IX
W3SWS+SoXAp0Gtp/MJXdBI3WR3pDgBSoEqu5LWygjUvJWBfl6GJNf6bWCs5dFtK+D0g19DT/HNB1
FMClzV2bRAQckLAgKOZqxD0UWgxeyRzi95I2uK+BpKmLKj+eftZAFyljcgZb+XunMfvVsKN2zcfT
xxKT4OOf6HNkZS0SQceiBcy5ZMlYH7eOC9eGnF4Yc0FIpJw0ZS+hUBjtRWcSuH6tQrwaOgDDEudf
iXmJAjvxLsdS87tdXdz34pCr/GEWXVOhSvYX2GBG0DvfsWJPIPFnBM1644/6rxpgG81ueTR66YMa
IdSOO5VRiJYdSHBEC2c41OO/o5avOOj7YSgl7/9rlr7u6F5almH6jzmTGlbmOC2Xw//31Cfs+ZCg
vKZMD2/XJv7NlMb5KC1PyfCuiOpmZ3WoB+pzSs9tKy7zkBOt7jFOEwmkFBUDnxtaqrt2Jk21hPuV
4uu+dLarEzoInD7ov8/TR2CzNG8xlOFDik45PBhqkUEmH8Grc31bC3n46qPcBqlO2gk+2Hue6k5m
qDdODW5zqzBVvshw6pFDErds2QzBy2LiFwpUsd5NxbEYw2bUjV5a+rkWaLGSsi4omMwSU08cq2xi
Qj22ByY+R5zeia86o7xsNwBqy/+F5FwFAp4/3BYZX3I44wLiEI+MhjAruj6608iRiV+2Ec+QWWvQ
Xk/uLwYo58k13KVQlnfqe0ZHCsaLPPOqU51OX1mNzXhR0ZYb32YNH1bvUNqoODsG4Kg172QBUSwh
8Tj05Mr0jMFmidgf2X4NDwBwGaukQyawrBtNyqHWoxI7ommadccuP3y5dFP9Hw1mAn/85x1f2My6
1Oh/gx2uu4qinv24pMXmOTCJzOJSAxgXxTIhe6ys3AMePqqwrUuUNxqmRmAyLhWYTjTpKFm2O36S
98x6QJSbJnXRdBvtrHn13mlbavli5VvrlqvK+pHcUc45SS6PIPV+DcU4aHXu+aAOetwoKsYs3eBp
GQy51ih6wwzhmSrTKwOPvB+9lGnrIlESOtHxM5GTXts4wEIhet18FVG7VzGIDVCq7QEiopAGrB+r
h9rg2WjQ3IpmvlpdSRsvbSiEQ5kMHlDStXrVEbZjLpL38fwqcP7gJrDsUJ7z96I/oYD4bw4Bkt4x
zEMDKBi9JxXUDhQXhfBCWBouK/WpLcCCjY71FuI5RtxpVDvoJKd/aN2lfwyVAH+f/kaSLFCXpHIu
UwWTrvZlJHWY4P+wAF9wqqyc32oHOu81h/JxYxBm4Jsw+FJYvlKfCAoNW+U7q2tbi5xdvWF1nley
2IjD7ZHkEFPvqtwfgJ//1lgEAFknUnQUL7GowkjZVQ5Z/ucKr/D6AVh+Q6fK4Cigg6TTNf80fTNL
eY5bzXmWqXp15tVjZTnXwJYBTxI5YK0bGZTYcahyoW6z38u2xTloEw4y9DDnCf8uGssTWIt/foi2
U5+U+LjvYl8yCQt8MUju1hDUuk61iY59CI2MckaRpllZanNv5qrIdOgFWuDXy5w4hmKiZl7GEdUy
Fv2ucllotGAKOW5cn5GC93TDv+I2aupx4zkcbg2O9N3CsPvw9wKkzFSqUrtlmhIBFF5jphbBdXD+
m7kFSc7vFqX6soS/ZRSGMj5LdG0O8vZVwgzdeXcgRbHmJl51dJmw5JsHZxXDJJRBLiJDECzgUmNv
eb55HtwEwzk9eO6zCHBuX3pea6uc9QTkz2TAykN+xHHa+3wg2OMneW2iNyFuNnPGDOmvd+KP5R8s
54axVxkdiNEsReUbqjgkMmfWNiBAy98pnfzWL7AXWswmbWLPDfK+ZMfQkozKI3NuGqfqvnOC/LVw
eP3U4W/L2dunl1n75jq9bFAvNbmyQokwgAIO30yFoFhTG9GpMf9ljLZ2UyP8i3971/9Gg3tGYwvA
VAnjzRL87E5sqq8DRt5l9UoCiAlGyhInrTRz0rgyFXxXP76mia0js012oJLexXjmPxaWLNwTUPXM
ZlZ/aNtuaoZ5FI0ylw1M3LPFP56+ztkKvTySuypsd0VaXMdBgEYAQMeOwxigcueabhqVm4TTr21X
JKZdo7dhcv7r+BJiLLmWXiFJY6J4BCTI+8twoL6xUFwkcyZbo62hTe3eoOnrbg9GLVdGdVxAh52d
5mNZZmoKHArYWhPdaj50hVQYJUT3rrxKSirq3Ao3VQ+fSDsbZCq8Yr/JWB7eTffo0ouLplnsC3aw
jH98lHvbaB28R1+JsobZMZMdrWplejoyFXwD6Bl0ErYiXXIxZGV9LAyzW3ma3kzB0DYTxfx6ca8p
PeDFTT77X6sr4fJhJ8IeESlWbfrvzhJ5wh7seGbV/qAk/drVmStbfauuyxk3koTKrYAiGR/Dne8c
FCQg/dmuBI11vzd3YCeUgS9vnHGdVuKhmB+lSXS6F9FFA6cTLiJzQgmV+hI8p1+QQ0GALr9NqMKp
C/cHNqJq81zOcSJw8wxkDYsSNWUbflZyddz2CwKVlPsuw5KbHuhqUOVQKOsCMztkk1oXUOdhRrlH
gkkQ36AJSk+ELh2G+vUMs9xlUyF2riKuAbn2IMiKTY2W4QIg+Y0zpMrVoq/eBoOSjQnQh9CsqyD9
5fcNx7yAM7OaxvmAvbf92n8cChVmuj3fm0DTK+ArkLmlBLfRYtNboP6K16v7tjaUGKcfMBSwKSyp
5scKPhk+i8AV7xNNTLhRKV2zsxiw1hTla4ZshYqBfaizUfGJS8kv0LLJ2rL7re2qGhJZUSo1stTp
atWcd5Tj97mQdDgNK8gF/v7J0BhX+G9ljB6h1AUB9TaDu/OU1UXnk+hcqH9+XRNUB3HocuRwQ045
P0UhwWH4qNJa8fFLNZ/9MwsrEybBcFo82+4/ook6FmCmwR0GIHkcOLoZ7mCe5CitkTX8TI309xBi
yUtr0wYuQ05N8QpY4idunJuhI1/GNcdUXa+9xIfzbbWHspg/2B9jDXF4kB2u7ziPfR+Q2FOW2h9i
Kk2OQcx36Oz8shnZ6ptz40NrRFiwZ4dxPISkInfLg50wTpl77/IAjsR3UmDL52aFMpzIoicYtulL
3BxBoucikFh2iqosA2uCsNH71b+fVfkv9vFR40Lc8lB367KqbtD0AOy9RVNSDbtf9yA5csup/eZr
BCI7Mef4nTdXedzSliHT16HsJbYCujNnS+/HQD8BdO5l5kuIuWUulQDE1rzGiZcRNq9NyW7OsU9Q
S64a1IFmc1bfTcVjqXwurTf+dx/JhabiDWGacdnAGYWjEnpMDyKEkxA1ub9L2IYJAi80QMpKhEi/
LFjEX58UUIZYlDwzja2yhcBQ4DxJomcGkiswhSBvM6463r5y0EPiZ8Nk7NoNgJsh1370GSDPnCm0
SbpTFHry6gVe/ihtEYUI6t12LEQbuY3K7/cIdl5I9UcGl4FN6r9F5K+E3u0r86liEsogw9+q83Ei
aNI8ksngp3IJ28bIaG6p3v+iSCpnigJF79u25qU3f7EmDIKuRGfFYdnR6kFhgru+KLpUychu7EeZ
7yhQq43K6Jkx2xzqEAgQXH7RYvX6G7W673U78abZDsBxcSIRIV1n4IPHyqD2K8BHbUy03nTZRVut
KIeIaofGG7Zm0Z8a/JQbALbCA2dglSOKQFZ42peKzqDXs4wNFA8ysQwDEwenZfZNOPX7lWillOUd
HXj7E145EFvM1hD6vg/r2lMiBQWkW/0yQZMKzMBZCdm4NCxaHflzE6FPbEAcIiuQhXazBtEI/r55
RtMPp1+3BpPwhcJBcWTimCOFufntpthkP49dlm4XboXsu3mDvrJvfFjtVfXBl5RArIgYeyA8laRU
pg/TBtm6CF99jPb4zahW5uTYRng7VJ4fn6OlH0GHMrGbvEN2BF2eO97vNnaB1A7DeO1Ee3PHamF3
s3YrmbULTNls/pReGuqGmpyy505V//oJl1N8B8ssYaa7ntJM5l2Aln6XatZ+8a3c4HRE0lG00CEi
7++g8fRojbellstWrpxYVI6jxXss70YbYGDfH24fugO+F/fegpoPn16OtHA9mKlWQHs8iYMRw3A6
kyefI6X3riL9wArXaSbmXOFy1iqxpgs1WRtL7fyQ4RSyRajTCaZVOt1v/QQta5Ru97FFfEW3h/kA
l+yg8Y/sU3zIF/XwUm8uELSHmzcgRIbwuX8XxYK4EZg320eafTMZ9qFPp+E7npMAx1UMhw4+/JM2
rviLZTFoLjzZWGOQxFx6uYOsYv5Hhxzo3Y5mdWjtXf4zGZZMZNlGgZR2W9YU9xpmLQ+tZghRbHRT
y9hZDgiUnitzUw3gmYQ68iykMUw9gpINZ6rmc8sS/JXMplDFUYQein1Y74bFcjY/jCGiXGhMRQkL
8wPOXTwhXUsCePdzlwCFJqHt/heVDA9q5GGOZD3fnbOs/AsHdb7i8OLqZZptqwivUS9ZOqUiT/Wp
PS3zrPDAyNJ6vu6TwTO2KdnlNdaj3bL86K8PbVhL9K3nnjGTvG4/cFKn1t4bwpU63irDsOohqy0P
mD+z0XCBEfkfqJQ2OEz55gBC14YGJ9bz2sw+zeeIP8Pz5/4agmVQmYPXvBIDBBWUFtzt3L4fSjr7
760eRMq47IefYs2WX9ZVdEG6/Y545FUTSy0KPtHWUOa0Kt10twQdVxN6kz9tTrI+QZobGs5TJgsd
fLRdZhXg/iLvW4WX4aqx247M7TDdpQQAXJFmw5+Ky+1XmLIU5AYkKKFTgCfFQ/sV6Z5R1yT+Bqee
SKdnOtuNQUem82CQo7GR+gm50x3NX2DUZfMxcEeZWKhLPhClPB0PD+cCOnkM93jBdEndZuFcTxwK
iXU6eBjfcgpCikGCvaDZplvz3fGVOO77Tl6i4TUQ4ZwwDHD2x/4N2GsvMXbX79gYvejxoaJthP2o
R5uQvwqVoBLqNLhWnbkaT0gr4SNhzCLFJPzKjIi2Fuf2tbTXVH5lEC0JvgfWX7KYlJy3D60ZGeor
mdWHwTKNapCaIVbxn4BRF1Guw+ttSekBR572YJijIyDqEWnMMQFA9PJQNowItcaIcZ/92Yc4aOsX
osxHJ2WqeWX77acSd7pc2W/UslL22ZoFCHpo/tgUtxzb9F5o49bx6dg4mdNFfeByu7Z2Tl/XNGs3
vKy3qd2QA38Y9TxFCKNLWr+Kwg8ic/rfvErstQsUzhnkUfvkiP/ZfCM7779Ex8u3ZFQfCI4HGmWw
0NoPchEx0veKNRUNkm5xa1qakcnoGDajDl9wqxL632L8EV9kjJ4+CgVizMOr4nKIml0kUuFiqaPZ
meU/R+VeHgaGPTdGrhhT+RNKRuDm3fL3aLevQuAmLaVFosnlbL6/WGjxL6YrAS7+zV2sDBRpmXN0
n81ne1HDQGWp12s/iUht17KkT2EbkeAm6LdkfgsOsyHZmvRc6P51Sd09O3u4XK7hyj0u6m3UvWJC
mBlgHh4EZPzHGY1ewhdrnjbDBVYRc8d1Yu/cM9Ijl0qNq0l7Qwq0HIL8rqYsOh7IX4GTKit5whrd
A2CMynAwFbXXQacfjpJSzEHZOJu1C158//pbOqvFlR8Gluu/L9/8T7SMJd3WJh9dxqUORmavJWUE
rqXxMC95VdCbSFKQ050UoU5o/KBI+oGM01nwGqYrQuOulEg8JT/PxdSi19tEWO/Nehb+6hmcRsO0
j5aF8txuQI/aNWjNj5DHMV7ZEhISiO4Sj0V2ekVUoYz67dNGbxMB/ni9b+i/DljcHuyvga1dGjQg
VNLQyQx7hU+1y1rchUSrlKMlzm5cHitX7GJwE7hzwNyxEqdJGh3/9qWwOWHGIF8+4mD+voa7MVLV
vw7+fuyaZ2NCyZnAziCP0NpNanTOuSCFldblGGoEnZXvDQbZZCFcRBef8kqrsw5AUkHHaTGunT/o
RizaH/i3cOOemTFL8v9EiTaq3s15nJFq55zG3OFADLXcBfBfhuMbGgWcqdIr2Ncz9IFkg/RFmL8Y
CcMrr2g85tqlEjQIvJ5xk0bOOe0NCI5kvXVnKuUUX4ERSpSZQ1GkqV692GbonzHJQxEz1oNVNB+w
bcLYaOtYo2/gyEau/fqe8TGtGd01vxOGLB7jVaf8GI3mJGrKlVePwPSarMljZsnTQ58FPodU1442
snGdCUCQUCFO2Syl0pPoT+Xz82Ea2SruI8xA89XmSel04XPy8+tvUFxzPIoXwBxVHrEdcv3/N4xu
b+Y13KrFhuixsEpRtd9o+blwGBPdIXZL2pPT/YiNdqmugWbd2JqIX/8LbedcoxWCf9KieNRfUlyE
F1zKFa5OPAMuTCWsNCp0X3pnXPufwSIlEvwgbEw0XdbbO7NSU6646XoS1vVSHVnbA3bVJ34moUI1
uyfmTDsBuJbf3t2OuDPMk/tH+JPpsCI5nkcUjEv/sCnmH3ETHy9+Ar9LxIRqiOvdcBq81Oa/BvJu
dP+5u16ebZJoyjBQOEequMzEb0PmHla2dq0RapZx1i2mBosJ5KzlZ/Tepn92vpUrmzuZQfby3DOt
htep0As6NEOgKINJ8kzv4at42CCfJ2MaHbp2DVYdrK2xAiHSx4EKRinfixDnUYNNpZM7AB0ef2Db
J1Wjff6Eb0HE/P5NrEZw8PkxDgS/xKj4nDB6yG7tDZ6u9T1Z2MVlmJwHoxEwEgZQMHWok6Ozmlf/
UsrtYL9sxjZePFAQV4u19Wilgi00JXAM+sjtMyzK+0yp1FvGLMVOivGYAKPypkhJA0M8q8+a2tCT
iSEMHcI8zAhnGThJvyKa43T66tXBV7IZTGPuanVjP4znhhVmHhRR3rii3cY5ZgQm/RjfGnQr7Dwd
Q19bpIJxuPdZu6pMWousMVwy366jaxKcDid/ovwJ2C5rCpS5af+MsQzTWxvxMVEIhny9iOe43TFg
KCxWRplzIjIj7tKhTA7ccOLO52LJPDi9Z9ZOvDfQ0tqC9QtLGRVrLEz/mbA21UkYJX+O5/8qbt/p
pY0YMPJikcGmrx2f4Q1ZfIFkcuyYYJE9IQIcewGyFTlOZTWvRbuBTCabo2JeZG0oUXB4hgcRNjcV
0C1eFlXzxVrLVZPSnXbCKPsBDytH6chhs6ajN0UPprO6+L8hs+h/euWDCERwSuUoqM6pac9VaBdR
3F3oD60jO2Pp/yXEB3dw5DYEpE+xOdztNAsGXvZNlBV1hxpCtwmCYu+xTXjmojiq+2SRsM/cIEER
+x5VOQauPiJh0uG2Qe+85HZlva+vNplbAMuK6okYakEykTiaKXwX1pEJBU3F9XzK2ze2XkI5a5cX
FCOBPGcvJr+KC57DvP2YvxwSCs+Fk9H4HbkoXfFCNjnVjK4D7Xn1+M/3A4L5r8jXrCJsUmfS9TRx
hGquGCDb0aG1a5eGxUC6N+0FpF8DzrCH0866Vvx3RIYlLAt5YwtaR5Ns8VHoV2avOiZXYKdJn1aq
6BA509FvsU3t6ydqwMBUIXBAAg5doG1XwJWhdl1VkawI0C3p/Wj/FcoBrd/ov8X0YSoBHPL/Safg
1koTBDfZFb9Zl7mTPY7pudKg0ByEa5yIYT7/iOHiMvmk2xZlTSioCK4SQzLg0TGaxg4oBdzWggRF
/w0Z75e5OLcc4ZkYgkes42Doz5sKTlzNPY08/EGaQPz5rZWGzV1f/p1DDyGA+5reXFtYJ36PlF+8
yeGTVXdWZZgQ0HRPhnOvwxcuXNAHoV8ve/ldDddNl52cc420cgTsxgHejYXO9rrFLMpGmrDJltal
YF1X6bfVmx31SgYLmiUkQSl55CRgEToBw5ufBz61XQGBOmUqeHWM1SHjh+pQTlTXiRKKZCNDRrIt
a0vIq6zu/jARjweXz3R3MRkcyXsi5MlMGggUqCAQTJAhIxsXR+wqaYr78C6HDr8FWDnine+1Yqkv
g4ICjZ/nPw/eWOHni19YeczZp+ynpg81hpVBPMpT1mc9g+2H1I5vDUUku/FfFj918FjYRba/9g9s
zCjS7oPzkCdf3AYxgMfOWXGKKIkgHmoy1GPoNpHIlCzfuRBcj7xhbeujLD6pXz3qIZtXbnuNn2oK
qS7FTZMFroDDKKlk26vQ+1vxb5lIjXTn+EVb+J+K1jydH6miPHc8j2nyWyjRjkKg4EhkebG3BfzQ
CHTeeNis30RX9GAVw5OwRpz4g+ti3y19vYSP/Jy/oh/XOUivilizpSaOwIQiRg7WQW5fW7cUM1Wo
2Gd0mKFGFejjPag3ixJwqs3stjK9+N7f4T3gGBHrSUj3P3lamWoGfsStBJ5i2AEywPCABOQL9OOZ
RFdq7A4lelCBTL8c+crgkBg1SceKOyv5qVK8G/0wL+nsL2BgHAceXcg7rwxGFuGmwNtEaLSKegv6
Tw1B2oyn/8FbCixwV7HMCyr98vFKo2xATQaqEPcv7GuA7tXscLv7+iXGUXu6O20rCGU1brOoJhmv
tPBfPaaLYhVAnrG5V7y7jf4Cq+SRn9v2EZRbYpESW2ZgCn4C2MwKZIqXSltITGYpzxjG46+VEV2g
jUNwuaf4MtWeE3gb7iT7Bd/rGDW/MjSXT8DDhMcflTHJ+xmWDaoMFc3sM5lup1Sjryi3IQDKdNFJ
E8fxqI7HF6NyXecXfdV1D05xam7gtgbwngbZf9D/dvMbs8S8nnXxV4DFtgkuQJihYsCUld0CtUnM
HxKhFbnnTtao+u/P1wUUC7ySyW1ansGYud3JAii+wVcGV4zb1dNHdUW68xF9Y9fxxTvzE2+CGV6B
aAojJxyN6z7jNZVaA3Uifz9yHj8ebYrlZ+HlAPpImcUQrxm7cuTEp8dC7sRv6bBnqHVSyjxB5LKA
4daYNn7WrEdBYSgUZFta9S3eP+VVe5FM2KYC6xE4OIMcBERHHdRpsnXavD0sfnyOC+Jxxs47eneY
d5yVlTxRy0xjalGA3VMpzyR4MbRC4V8swTLXMvYQALUwWltTxz/KiHVEdiAGl5gIKq33EAEv0Lof
i7g+lsgqHNK00QBS/Hbqmz6cDkUPG1uw6KlyqV+slZKq4zRkghkbENw7532ehQHasVF4CzcaaylA
/vd2qjzvwAdmLQPC93SCfDnje5MlG096YMn+2tv4/TEmvXeQFPqMp/4GhWjZ5AJfTPG1XROqO+bt
Hazba3BBu28gnFSeajM3v74edw4z2Jb9f91SAO0MRX+CVXqcGOsc5swKE5OAUYv3leOos0m2jozI
dacSDd/1k/L1X6Je8V2Kfpbvfo9baCG0Gw5eoe31AVGze8dkTrdGrDvBe0IJEKdMVoMVxCWUK9lr
WK/mseuzX8XKKTUlpTIWYGcDMowDICbqf9U196yOO74nY3ZTAfHk1IfsJS2pvTVYAGxITZBGOmdI
CmG63XzS1LXpTf8vmO/J2pkYLe9iuRm7kIZzeWu2KyeXyvpT3/wPQMAacOR7EdpTTV917KXk4PbA
ZtUCtCFS7uGrBjJ+u2v0WbGAClJi87khyC8H7uYGHBN1QM3J1MDF87xahdgFVzStXhTBLv4oX93d
OFRg/gCyJOee7iXQZhfnE2SteAXQQlQKW2j7lo+fNgJyyhiutZdTtT00NrDKngv9eZNUCLIlkZQi
bP6niecadnojgNNIhBZX6UNZ2b8kQAEJhZN5sZop8pg1uKXzcQLFzOgmEvtUo6QRpfuQiEcT0E2X
dDozqP4BFzGwZ/TtTXv5ehpddfPjXFBRlJw1Es8B/XY8cvv9gmwMrJejxy0MoKzmSmCGlSKTCssH
sc4R/caWtxshIp7kLWSlVgAEYQw4rm2dpI9/br075xOiXQV9ThUgSOC0eQCi+KMmHyZp846fj2Zz
HMubrkT3bOuI/QzzSDNKejX+dANFi0xDEHnmWqGl57GxWp29YDnvebY0wgLDBA5rVtQidiaR+aaQ
X5fXw2v0hlB5pHLmBBNpWwWBmQA43jAo9zFFG9JHD32c5ulV05edOTrrxbTKg/llKhVs9VWo2Tjq
+I0XgDBiYNHh2li/nP/EXW24lQ+kTT3V+8eMGwCGCiL3YnRzs6I+9iGl6p6tPnopnzLrY8BGbal5
ogV22Ec0iX7iuNWnzSU8qLNqTCYGbBzmA08jhKv81x3Rv/UKaC2eDdjgQW6q/0BKqTINz5Wo/0ga
4eMW/6wrwM2hcT2F4wIAU+RgutnFiWDK3fCAUQXHj9pPjxtuV/VOjyHOCv5Gu7P1F8BsX8vpBz6X
Yck2G6UTu+dSwBy+xAft1QpbIL2s3hhCnaCn6F7CrCXXW8HY+jWCZxvs1OuCP1qQOF8icOk0cBz7
0s2gvPUWXec2GWDUvDxOv1UrwbEW/weqHYhExnnXmBEtnO9/QCImNlGVVBG/3QnIVsOxPyhhmgph
ths/x9B1ZZj73+EdX2IeLpu1psEUEUZ861SaqGw/arXXzqDgwrgYDcclCvy8N2A/2CPDy+pBOob2
W1O3hG0U8ZwkEiRwJm3fjsjgLw6ZqbYQH3qt9kZ1W6RKktsJf50y5UmD9712xhtDTDC34utUrDHG
EUk747AKRWnPpAz7Bsa+mUkvotklovjAvSEQUFmRjxD347m4zsxE6x0qBrgjicDub7LXG8HKG2V5
ECstwKvuUDvJC1zF+uT2gsW1DWLlWrQ3Om1XBL068NEHiTuMRIRNhra9fz+4bHK0mIvOILcp/R/1
/yKCSIECtm/jEWWoi0T0qsxJvdJSG4s07pqkt0Mvq1eQk/WnPwDKdE7xUGZ49+p+fCdZ9sN6AOsj
tA+pPSkpMswVIghX0BzIyhUQ1ln6vjVX3TmlO96W8NlYY6RdbqaZizRUeE85JypRtTBy0T1idDMZ
ROEJfNHbNvLar76pKoSsO9okT6Ysj1FTYGJHPWEm+61Fmp1gpmvdzBmU/7xEk288V8FHNViCNgrF
LPXvS6b0GkU82ShHV5bgfWfYFLkSP6nYu3PZYgQ/v1Zxgm6cTv/Taap3KCZViG9PqR1k7QSgM/6Q
Zv6aVKGNVLp/g1/qwW6xjQwOpz5laKf4R3UWFKSbSjMUurvf6ePJEim7g5HETQ2+tyc68uevOqta
aVHmiYrKD2RaLb39Nx43ORphOU0bOd+HulqfCndOhL/kp1BwqgUbisLVGfaJxmZjs5wU3fs4sqFB
ck28bRNT7zMA1ZXjo7zNJz9pawiwwfQGq7SzoqavnORt3F8DqY29cqSgUNWP3ZB14FBTKz1FXOKg
/pJ5clWKPNhJU8ORmEMPRnWfq3QSdT4ayoB/GhUn8uGpLt7KsD/EazALKYObwae47TPE8+mM6YTP
G5T7EqmzHQ9FNg2B1gn5nEeZwwHDQyvRpmVmjXC/jHEmd8giPwnxePzS4bSU5cnjYTzWdKsblpbR
i5li0ueYB1RI9LO9YDpB/gw6u1P3tjnM+M0N0V/0ook+m3fR84QukB42RbB+yNiYH8lidu0S9sAy
hXDZjH4PkDb4CsAqz806tSYe4YOMJV7symiDhLN/LeayhwH+Uw7+Nprs0XcWPH8nLxqQyjXc00b4
Pj5NznLJ+W4plWvfQwySQpTdZO9RpIKV7rB8SrtXSYlZCNN4U59h2a7uDNm6zpf+VqYuBJ1TjCaS
SJXhn5nw8RtCoC19LM2GfAn01g859iRK1wDOGHOL7O96yFRyCdxU2DEYFtQZ5uzTOKELSr9Em8uQ
cjckDl0xd4X2kVfpzg5Ts3XiXToYXKnxW6pU16pzR9EjTu98G8d2IUE/BcRM2r+owTQU/q7svfdb
64LgtoaiM6/qiQWCJ75V0K4wmi4vjlkaULxl4r96vb1KCjAF78TXEbAaT/R1u5NSZ14wJ116szXX
99z1TFAa6epzCPRQwfktKU4/igTRmLzeYonVaBhu/anjFX3B5lMjF/tHdzMkr1poOrVBElofL/Vt
FeLgfNOUUpofz47dCq6OwijBsNHhw/6v72mAEWYBK9ho7Jt9hex+J0D5QL/yXn9rF2i6AcUCmuuE
kcUVs1gsRXIHFT9pWXuiAbycxm+2ZNiNLlModFQVFN7qiWM1BKO8HgAqSCjs/+3qNTToYqlNMvnw
V7RG7MqpoDO84RKMt8rqOqDeKN99xcKWs1sBewmQJ33gBPcl4ja0mVRYlyJAtvWyL8huX5UlzX87
c1RILSYPIwiKA1zfv9EUW0YxcbT5ENEoEU1fol4G5sAGdBUHHAXPY1IoWfRKJtFdGkknlF3bIeMV
b7HdUB1QhTFSt48jpWRYMMY1CvbnhCIDKV0mkS9qp12VNKI76r2qkyqUbvuN6ukp0n7tlH8qDFfJ
JwYDnhsySAj/a5EQ+W/iyNzh+u9IWTXYNW1qyszjqh0OvzMqGO2p7RDFN4U9/MHAXIhVEuhq5kP/
WzbFsJ094QfcGlb/Xyiyy6aTcA/zoIMF9tbmUNhnLZ9Gv8J15fTYS5nxgES1pASDdGlOAB0YqMi4
FFlVYBMwvwJ8bmduMBJyICXnqkPzQLE9PinJqwD3tuq9vLcdO6EA3VyF8kUGVHtcKZ+Why83JoDJ
8ppQav3jW5lHZY6S0udOIpnjxQXiVt4v7Rhs7JHTZsq72cWD0pEvC74K2xM97KKyZ0d8EbtolxrF
iw0f39moGU4SbhAuc6bSAgmOWMtOhM/3ZltAZhWwS+Db4klQNZDHKg3D3p8inBobyU/HQ5LCmV8P
Q9OZ77ESf7QnOQLPj8y2HBSHXeTS+T7ZLiD8fMnQo8oyYZLOkPRiTjK3BDVEYpulSSeIezk4zfTg
4Wz8afBB198SYx84cU7oHhFGAxYZaUaCaGhaKhD7jAvunEsKeUFAR8utDDulV6bQPP5euAbg8dTZ
U7pUts+WFxyWjZIJLrD8Id9c7Xr5GAf6qpWmnwGpicgWHS0BV0VdPYdB9cqi2nreV4/mb4tHYAey
lBrtimd6Fgeb5vicv0NPLecmN01JJrJHyp00exj2vjOes/l+PD7IwjMBxH6OnlTsULwPMkH/9RFn
nL5t4TzfrLcZy17sZ1mZ7fYnaPL+WN6AxMCsvQY2h3fpg9EmAdf6dpYCTXukkwlm3G89Q+yvQ/K3
1dRZXjTj8i5RFT2rpiv+C+fJIuWU0+AZM9yQq+PzytV397BFNIqwSCyhql+2oLYS3cCSIWAAyHph
iFv1TqF5O++aGGvS9XjEuGCmlwDn0R8Y3bV8p94W4VHI2hmlOz3SFPvvnzIYIoXRp5v9wh8rkMWm
uILXQuO38zfGsu6eshZZr0zbpHGgNQFosrMXlIbAi6JZ8DlDvbXA3Mrz2hol664pcz861A1pmRAI
EXXEt6Nb3HRcqYNTEOSou5uSA0CoxeFclgYSYLJOESNJU597LFPKL1Jti0rx01pCfdALnW7TI2kU
MzF7fgkKgG5NXnt/IE+KK3NCyxLtYJapkPWcWjWYrIXZDdbhhuGzgh4Cq27pgOkgn+LvT0OF7oka
12Cn2jMAK1PLQn32QxjWdsT8I1vJVyNoplPeGfs5yqJxYS+cfRYjCWEuAX7d3O1gmJCzakNGih6Q
/ng9wMKNmq0pm/envTmfM04RK/N5VCK70pFadtC567aF84gGYcq4Am2RhYXL+lcEYTozuFrIjoz8
ZQ4Y+2F0asIiC0ULvNrBfW1abpQ0e6ISXnfDwU10xAJbY2g6B9VO57RbFs43/b+RxY0ybN/e6QPw
PFy6S4SNAEhkH5bdGKM+seAb8Q6B7wUwmK7+AiBAKgY1kN7nx2mxaUOnc2duFUeN00xh8Rub0zN7
JAx0XTXDCL3Ssq203vAuE1lE49OqjCa1EXpyRcwV2bP1ZEh8tS5CCv2RbBKAzV8HVZVTjPVyU7Yp
uTij0avOiHnzC4BuTshVVbEtLf50FT1kXjsPp68sQrdLOJIy02iGbALro2KkQ/mc350aOmdMCSuS
bni/YXh9R3q9iqbpKsX895LNUlt2XaUSImbAXPI/zrC/eOOChWLdvRAjSYfLL0QOtDdPL9MEWnIM
TbHNvIxrty12+j6Ef4K8XGxjsi1XublLxI/SzmHJv4AiFc4eJ+I/0LFS1CMA0FfRIwiynSCvqXa6
pixbZ/Zt39fZXMXoGDPv5VpROuczRY21dsI1Z76FjSplyKbHOycFAxczsQ2zpFkFIknOSjdqpW37
FIkrS0NjyyLXGuhae/uugaORU6N5Mbv4KXuEdK4CRpbGE/exSzwDy8qMXDX8RicGPfisQEiPqTku
ryv9ygOUWUfWkrK51zatne+i1sBQH1dGb+Xz88HSxau8ESaYGGS7pWMCz0dgoUmJgpnupGt1VJci
r9JPNPsRdrx7KS6ZbWOszryGggZHnCX5WsaHksJ9owHbViTHrWDu4ivj6E7X3qmFSlV+xFIoWDS0
13FonFxBOQytELVWvYkBYsuIq1reVh3SNXDxC1cHi6N7o2TbVBLL3bBEoJPxWzmC8JPMvRMF+ESe
6tziZV5MoT/GtdlM3eDgH1DT64Wa53l02DqiU2JUg2v6YTirA8qLgf34tjLYSv9T4LJDkvLeir27
+iVtd9pA0iH99qqbGP5lO3xtHcOy20u4w2NI187EKkdnkMutRUNgYEeIV+s2HgxPwYjPRmA8s31t
z9Do8xQzHd4DBvFi1Eoq/uDXyuct1vXcZ+Hdrku8SOHZEcyPiLsHb1n4qk+UAwk71QfUXqV+eazG
6M+t8IntyULA7Y2iV0A3JPQYUT8m2CAi4Ca+FvM0XUaoG7zxWpDIJTjL0ss6QGha66r2XIypFfT4
wbRRl1ZYgX3kYCvQ1iVd8gbq935HZ87UhqVtzRdfWuVCJkgiX2fePCeFDF/1ImfHADofAxjEtxri
JJYfhfpE8Km+XGwai6F6Xtls0aG0XvyF0UV17ttHglZNUNBJ/j1uobPYS7jv39X2FWMF2qhPA4To
S4/DhwEmGV7csZi/57Ssd7b0PdWpyKH6LXqp4sAy9Ecg21GuRkCPr9IpTn5rZHizhh4MdiaZxLkm
LRihHRqm92EZJ/pwHS3+6lOYe2yy+fDqsYMJY6376KYClZvMgHMYWIprEzynAs/GDt2PJO4zLdKs
H7F4Qm6HiBwyTkOj+48sx2pj+zBHUIouCws1LMGx/dOZj8OlVeE4ARza7WilUTHSv6nIGOiKPHp8
aF84Nat88mr6ccC9dYerVMSHgJBbpLQiA0OorGWjnJqtl1UIU1qk66NY6AcllUgIx3Uq/KUBXvdJ
0s+TF7kmV2DcYYPJrZaumKCvGKJlzwvbXZO+/hsMie1fEuuArNMI2uhrdpeqrjLy3ugM9/yfqpbk
TyE0cPQMpu9tm0eVo7YeF9NJkC6Lq7zKYo9Y4ecTdnvVO4iejT5rMu2dBQ1TrY29Gmf5/aYP5Tj0
VONB5eEWnEEGyZTKTNNauId18B6SON41fHMzt74axqP8gtKFbCBoiud8izuIn2oS6SnLm5uQvb3k
ftgoKfBb1KUX9xv/A5DfLH+16RZ5h2lFspgGYciGEPOK2oc0LnVtoZkp7agUhyp+vxBqZRNcI0ey
ZwGvcSpDP0QhyLgJnhf73OjK/zXCPT3/NZKRETgMhZwjvkdssrs1mqCaBskp3bz7dgUvmNo70XX5
cC+zn0v4wbnMPKMgbkPmTBR8JqEcegX5xTXX2jiEIIe7cp/5sAoEF8kXHCExK+QxdZIaA9N+UQ0m
+BSVCbFXO9EvQEPhLtQSt4j4fb9Rrvw8U+qMaPPOytPs4ZqFqosN+4K5O/eSPqywMkfOLfE6XZwu
y+0YfIVgh3sciVxwg34BZDxHxWJQ+B8bBkDsD4bjtFOY5fObkvA3zyh/ITvrP1TJ7CH5BxFd5AVu
iMQnB9LKS7/taji6nNzpyuFlzOwbb9/taT99aU+eHFe1bmvNKAL5fSuQYXtucp8CoBgbtKa/ilNq
m3CoWX7vUg230nEs9U4djLO8pUGeHIGalsWkpgBcJ4/jE4XHLvC26PJGtnb9bDpyTGZrzPzQ2NgL
0QhAH2f9T05IZtkxZ2mHzdNp0C0PDMuSufzHAKX1SUZKdVrs+8fzDEpekGxTELuPiLjXC9eiBBRC
GvjIVZ8AxV4oTsYgExZ5XpE2dBT080I4y+Gqe80xRUpqRY/UC3Bn+Yfhq19iy0wY+s2yFUP5tKrO
ASF1eCmQmvDifZBF2x8iqjkbnXicS09+Mv1EnEJnmS5HInyvrGWI1+ktI6tMkSMnGHJk6tqHJsHK
T0LS01LrrcDZu0xuPQDlkS7aqWdcx0kQ7L43nuigpmZy+u6NP6kpMfSVbAnfjMUSnVaekqzAfgoU
Uu02mD3AavMsohIDYldSh5l6aeU726oP1v9qtjyjyu7vFypnoaiCBjVzCh/pjYlPrnXNUa4liHLM
4xDX9Lz83zN0T8VTkKnO6XS9Kh82yDSU3J+hJsHJimPDb6OdcWqFG1DIcHf+X6tt6DRwAyPxMyio
Jf7SuRVe/57PsDpltSrrir/xxsB4nxkZWhN81EPP7NBRKeq/rfYVudCHraBwMsEUhOO0vT4BveZL
rcH5mS2fweIclL7PMxdWqTLmNA58ktpIa2xiGqtsFE/SbSu6wMqBeIjZdo/SUdsEaLgWasiAzTKe
l5rjRKoJn4hM7yzeFe9oNE5XTwrmuqTSjzPaZWuf6acLI2gG/8BSQoAXWasW0KfnXqrqa34f3E+B
gKxpV5kWg7H3IzF3Td3rtDonKBgRwuv2KIOd7uKwuIFtItnQCIHHzAFzp8v7Fc1U8v0NF7KvDfbL
7Rs51o9OoUKyYmJjHq7zWu40n6JU6j2sCUWIgT8xHFo8ayP99C4EcYCyY2ConkriAb0+9PuzxoTa
rPQToCP9o2fpLcUbZ5T0cx+ah3bAU8Fw8g3aG8atKDErKXYy5I6cA2wnAbRlZIsiWQ+P+G0O6QIc
qZY9Kvj9peYNQmeNUVDTF1MGkj24Lxh/kQtg3A4BwEMZfcstU5RNt/OC63oSh+Z3E1d9YcNN8Do9
MsESX5beSF32QLZLTvvu08P9jxkdqMpZePwT0yHXEeW2Ch3pTfbFXy1tQxfoAVKrC7w7Roz9qbai
QtPCq6rS9a3ajZgiHGB98aJqBoM4KM2gXouCjW3e6lr6UCsdSG1EEmQ61lfsK/N8qlbIwptOPUg5
dXus6dJh3R0fCDM9o0I9xfqJrg3P61w8g+FH7GX852cIjQKH4/W3d2SAUrJfCMNebfxffcXw0CiS
64ctPOKlxQXov/J+Y8PTpGGvMbqT3rPalzZ9JVEZuyBq6bsIzkg7gLS96Yx0Qg5lmEwPqc6Tzz75
zmONeyEaT+efxOrF17FfqPdGJY6ISJo7sqMRwpZ98LsHAqmZiW1fjk3nBRLaZygO/p/npI+vpLYT
FzX6suNUBQ+G9bTT0wwQ3ZRvOqKPADimzIZLeEMoDQdqYcaju8pNM4NB2DUf1aI9nyR7gOww2/90
fyl+LOlm4Xk2dcClu+wMmF9nV0b07MfBgKVgZJlctTWuJTbZAcdqmDuQjhSDA8OlMwPXmZkWn6H3
8lHaIgBaYqEFf8PFcheMS57l5JUK0YpLYyLXIx32c4PhQBgcGXgzmEPvaUPXfEgtkn6dVvcNtxiH
8S7+P7+Z8UUSZMwwe0nJWc1g/iGH/h5CmCurpbrKDPD8K144VaM8M2Pi3cbsRqi5NsNRnvyoVE4I
xU+RkhubouUxwz2A444iqOUFtcDGzgm/K1q89wGCMaPbJkNgt4sM08eVw4C1o6ZAMsz4pv8uaSrP
m14dNv0RDFIuecAesw56ROH8yqlg9inb7Uy8r2qXG+ubGyXeJMrow5yiUc2CQbxvblLUioV6KWS2
VKApoMGWUVz6f0gkkY9Ax+2qw0QVDRlK9YVG5Dz64kCotmXrelHJ/EPnzk/5biX0/jfZ4hL114Kl
cWpu2lsEJOubQQt2sOAF9C35HZsPVyr/BmBz3n64mNUBcOHA7dUQxyzfhQdz2xxHu9YueQF/oIvl
GuZN/BmdEJhzeBQqN3zXugszEZGDSL3YwyI19Tppmgp+jZMoQSWwYt1D5C2SsmzHf2hazR7DXpZM
fEWaWa0/XvEylLRg7nQXmSQTmPA0/XVYgoshWsayOG7LFNky9GQ8JfOOU4IeUpuWHewEJSmIFHl7
uIykQBcNFSmRiW9FG4OCpcJoCnVZx05eBtxKilFgd6ihHUehNCQHflfHxI09dtO1HDQ9WkQlTaBE
iocc0O7sKI6YQkbUm3VKwj1n/VYJI0LseC8bCYs1y0DJmlOYfOr/pfA9lSGqjUwrSG5oeqN8JkuH
aWzEpqHlYeM4vmNU3hWu6vuO3+McLEthTI5YE6XfbtOFPsyxp5NIkNoasDnDOdtXqWLG7KG3la/f
Gpetq5VX3HZdoudU8ytXt7deEl2AoKQyuh9unASBNBDaz+j8ETViHfehgswZ0VvMixJmOxeIFZ03
WRQuAil7Q0TcmzswhAQKkADajsHCICi6rsPHGaZGFYSsjPGpUx6f3SrVbc+dRxO7f17hZTlEVjEp
vxpEhkxYnu/v3j8vW5LhylIqndHnTSNKqtizMHardwta4K6fwBwgweSX0uFvyfHPNhhmJH9gFlH9
fVyzKYUtfTL5IVMc/T0ya6cpa7iUdEu+SH603YSCbKqTF/42pSGbNtCwIShSxTnDsxDRoEPhk4uL
mAGEzv8cXj5A048FjgCGXd1fSOgzvGCmYkcTTBFNH87IaDMT2uBSL4CUFQVNpMaFEhx/iTxeoOpq
k/iHCfqUmfibTggkaQL+3agBlGYTP2INmLhcT2a8ZQyul2MLNL9y3Hx3F+MfMBWMuZcTotFX57Up
6SbnJZlIMj7SJmJ5/ElXANwYVbt3i1M+QGbtzLfLz+YmLmhUknNkBtYXu1eei1tevjzG7JHB0FaR
tBSmSL/6sqR15HMNczx3G+h1xITQ80DUNK63ImCEJFsbXu4JR0PYq2hDGdou9rAmoNrQoU7NOCtm
pOMxfXBZBgZBQZ325wHmIsoBAqJxCujnseNs2k/lNFTEop9iCRPBzgSuzuI/pKsJ3FwIPBVBlZme
4UWgQL4PYZigjJlUsHp+p/s3fGQCIqLZ1S3LBWk2Y0O23I667qgnyBJUBUzqiWOXnaeTFaQYjXj/
gCBCljO+pApicWBMJMkIyAQpCA1lPT8geHaU6cGNt3R85S6cnUa/wFIPH5QLOfBwUxVwgM+YPo+D
fVd3VXj9JP/RXUlgPHhObSkjEUFW0xCQo2kez2mm47UomY0jdyOlD7d4Kfi267yq7I2oF9hL3kVK
1vcqbBDOMIefJz+XncvWO9HvfR7Rcp8nHMbvjgEAM9mDtsBWkUqPdjNpEK+G0ODMjtt+2MoG/0XC
M9aTzNGXv4Mpx6PIY+Xz/sebmVlRrEU6/AJUPrS6VX2h6oJZG6+ecy5vFcRUDJcRVXApBmGik1Vs
lNn61V8f+jqDLYKkTsReU3tPLgaXf9CT5vCgI01Wp12wQPd7eZPp651RYg2teMUGoLMSfEK4TwKn
q3s4ONaJRi4rADaiEpF9QKwnBhnD6hJtU0eYc1LqJDpdLyWx4RxENL5NOSKs5Q9EZhGsfS0iDqjm
hET8Xe/La4i6oSiu3n+q45u6yfhjCOyY0lN7vRIKtuJLP6cRsyqAk0NX//tUjtdcmGcAznONADFz
5sdcFq415UEjy5l42OKEHIvULQ1pq/a1gz0Unh3t3vjHn9Gp3YIVW6tWTwRnSbdXZQqkS7m0wVja
cWIQj41KIp1B1aLDJFgxJJ8shOcHxdlkpRgNLgxecQ4s8lECYDA7iVoeNh+v1dnz4eUD5D9t8X3t
7gG3WeZiW88v2fLVvaATb/mtCPQnJDnFgkyOd1NOkyWep2C+5TlhXbfMH27PvKizmX3Cl4p4f2fa
solXQLdQ4Kd55L8/vCzrdthQ9Sal+OnUoo3wj3EeyVZNXALVU3mE656TjmKAzx0UAVL9fRfh2SSl
Olw2wlz3tORxdlhqmKlBiV703H36OixenVJlZkRNqmr7oTy+oMKvbyB1ePjo3e2SZQ3xPgKHxTvB
WWvyj4g0Uu2CIFva5gncZsTzUMltApYwRe3bQxy6aCFPO7NJoxs54II00vIVbNipQxPMyi0Z36ZJ
NUSS544qzbwLDvxJ6dCUZZUQFxy+l1eN76VDpKmsN/xT+1LMeIL+C83f0l66xqkXad3xo0vsqh8+
h/duqVf2hXwsDSLb8MvTzcDMO+BLEmtSN3CrqpuoV2NMHA6McQx4V/V1ORtr3lNJkrVGR9FGv8da
gh7lUWdKbNeWgJFOwAe/P0d9wIQ6klPXNL//LYOVtzq/wem26RNovUtieVeHBkiKfSZ5eQFNy7qG
2bIp2FQfRQL43k1giQADVyoPyl1COFuYo7JsnOPQzi6IJZdlrcSUve7t3VnjpwU1IxgpalWMW0ld
AHm5glhVx6pN0YmODFOZmsdwt+LHmaKP+9dDRUxOj9om8Dz65Bd4q3Aca/3zJDFhUuNYr9xCeSir
hXYgXvYMHdLFlSazcSPgFfqK8hLtAAVdQp6aDQUsrmETIJLAhBwzDXjIzIBzvk8zEvGxjfGmDC6D
HRpxZDIzJESAT0bIZmKDs53n3T8BSPDnMrMAzt901P4PYAuIMzcFYLoPr1/Q969u1SO4+xAhJYCj
YO40vGvsV0LR/Wmrz1+j1bNKsOTwspzWB9y8olNte9uesReShzaID1Wk9HkLdWyWwc+pT+rEA1LA
5VPkw5ZXy6hJIniCyz7fcOaKrV0qbbQvQ4XU0FeUEzsujYVr3FyGgxfikHJE2K+8h/f6ZlmijGG/
G1jv6chPzguiaX0LuCSG2KZKJisHqB6/RTHlr5maVxSxWjIsXzMwkCj7cMMAvrv6K3uaRs+DwU+n
yB60il9rIuiATBKA4wbD3M3mVGxOJdSGZDUa73rPhc9knmkBrricsa9MZCcT0iVboKafvxb+CN2Y
myaU10EpldtGGjUlnhrWOlX8CgJn8RM+r27J9maYeYRHRuEEmlkBC9kherdiBUL4EP+h0y9BB+B3
ygCWI3eWSFDpryZIWKir2R8aa9TfZeVNoTNBEtyJweZzIiYCfPaGECTu3W6/wznFUMGPnHNcEQX7
hAiTtcWvrBuS50Uo329W4tkAFyIHVcsO5Z17TqXr54tM1577vqWoZ9HRCc0+9rORii2ygvZTOlW1
gTwl9jLRSFgoZ0XuPvDaOYNLKLv9kZFrZHLdyRQ8i4xsbn2CmeqjhtnC7U2zVNJZN57riImMIXvb
X2gVzNyJ+L5BJ3R4m1tdIEI37a0Od0wIi/h+Q/Y7PoC5stQM672xSW6oz9YbQKNrn/cMBFnSbbLh
m+8ya0BjxOkpHct7Fc+B4ktZQ5HIK1uMFOZ3dB8NkxMQ3SaYeiCMz3Is6en4fbBw/153FZAy6tnh
tr0MI4EBXlUImoXWZzKMWRTvGFiEudSz2Z2kEM82AUeDRUc+yveU97psytdARxZ2r4uavTxJSlNz
OlRNDjEcwbAfz1FJF4xVKjgrIGiZeD2pSAzdjM2yQEVbm9nNbz10TANqxziDsA+DoBbZrvqk1QhY
iQhDDS2oWrnEoJHCcR2tL9sQ/U8EDlxthGak/NIjOEJJ5zvSfo+QxZC0lmo8+oA/8qVXMBE+d9rI
+8mAOhpPk42ZsDXicEQgA8y3ADa0rbQbQWTZWSXcMzTnceljHWLPomBLIm4HFxUlcBZKDL/UrKyO
rA6uY/TsF8AqlXJ1KkvqT59BF6D4Qv6uT2aVvU+gPqRM6HTzpcG/8Nxz9PDGKDvKiaystrkE356i
eC9vA4DhQwObu2RJPXg0zGNxdfDYdYb0GH9IUOD70IMPu9lyPALaXPB7QFMBMbAfGn4ai12BE5/3
ckTaQVevFXjPaxqKIbbZahuzB7qNLY4hA1jztG7sTM73z3bXw9i7mmaSnBAVsyEojHcKNp6504Q9
D16p1CtxAVqSyKhqIQzlsOcd/UUqw7BexCJauLynGnTUS3PusCPl1yHyiIcRF7lhIUIijaCvdST5
HM8bybUOTvPhn5biDzSEsFrYX5AXdca0IS7EVVKdelfxbzY2+kXK5o7XuuxdAbwt2wyfQE544c2v
EBeo1vvqZUbp1RwqduxCJ208tjlPGK/A7QcVvFNgn8S6EaQTB4oi2c7mY1pKUcK+uXjq6eSTYHM3
V9TpK8FP89jiYekrMaGV+GmMi/ReA0MB/Xi5uT4XjLpX3Rw+kFXr0qscpvWJL2J6FkcQ2ZYKCXml
3lqd1db/xJkCZbOzkG9b3d3gEtrzDaHdmLL6szGXgILUiljtDP/pX7J4z9Wd1S8o6nd5gcN7GmEh
95YaRxVrvEBSb86lhI8UV87zed/AVeRH/L8a55tT4wCYMrZbuRTO9jmj4PpZyHIpHP58mltrxIhH
QOs64cJGiaUONjXqzDwTHPnZIg687RUm4fm4+o7qiY5NXqBOdpcuwWBvSFlpK3AKv1f4xy8e6YRo
mvAHC/VATKzJ1y2qzBdY03zW8wycV4Bz7dldDRWS6uT7oel0d0ffQLXuOT1cDAu/jqrs0t7uQ7Vu
7eiP9BUj35MXYldJrRMVeUtSBCh+ecVgsGsespIdYwd8uPSZL3rvGtttRNLUjdMdBIalzetBgVUr
OYAJo38PyKqz3M39n0UDEhayrRXjgOJkhuLsq67D9adtc9N2lh35ZeGKwP7SJNSXrZW8hVr5ycRm
yedH/L3QLCuPvKK+aj8S7PCIvIUiB6IXDJl5hlno9VMFL/1xqGeMPgVxIa/bamtOxVTaAm6u3v2s
kWRd6XBsRd7FDAhj8qmykQ5ElgoMK+OElrgyqgAgxFg9LOm9t1IaBMpUJGrWdJ9VUw3dM1e0M6Je
Z0ham+9+eeE7wkC8RIeLRh6erc4o08dwTMP4lFxlhH/tuVTqqdWE4MYXSeTuznutK+MTr1EUVlJ6
62ve8L+WgulH88bBPoXhS1DJqgY8kZ89JheoQNK+mWcNK+893Y5ywMMdfEUtOYZCOGFtU6Pe8q+8
TDZkx+Y/udVXL9tfF3VvS/CLDIeJup6wNae7+st97PFiM4cIsS8b/smconAwZuhkqYAj6tu/Oapk
Z1b0k3i0VM/VAuXEK+M5wkKH0RcjeTojDbFpNebpaQUQDS5c+bZ/xrH773BKpQnuONxEB5kwazST
rX6jqgAKoSSFT0eCgdf8w9TXxYIuNxeW3zh5gTw0qJI33W5U0Zs+EncjMLufqz44evZXkvZf7yuk
w1OxeNWNhTI5lxyjQ9Ml7rlBmPI7W2GXVsFAKwtTsnrMXCLuyf0SD4Tsvv+lkCNCuObkx0x1xPmK
1eX+CiC0XtNXnMM3Yr9UtvsjckpkSRx4MmZX5ol+svbVfms2a624YiV+akQE/avWOUQ1ckQ1UQI6
LsRyTZB/ml9cjnvXdWX4ObhkOHKm7C36qbVtHebMKEoLmkx6u+Ol2lAkfJ2kB2wUlrejEe9FgM0R
z0/SjOp5raQ+9HIgP0sBXaXB2w8Gwznr7w0ajA46Fv6b9eLrAE26wYRV5KCxm/TwpaMVQZZrotEc
3siKxgE9Bwbi9DBYbhZopNdrv+MtV3f64j1AF0pmZu5YP/HicJTKDMkbJIikONPxY39yV6YKlJT0
/m+9Fshkgbo/XJDKN8SD+cFcYVArK4CzRiwjU8cenlCb4d7i0tXbjG0qSCWaWzTTiB+l85XyK1dq
dtUheozwTgzOD2pjZrT7l2Qv3z2RxtEnbUkFtcS9cB3YS4uyIdTQb5ZZ10uSt19geyoMEO+7aqn2
3HhCLvFr8JGbvT9btK/d6JUNeKGlgTYNKYw8hj4xtIdo64onSr54PA+PJ3kd0UKFmPi+7AXVSXI5
81cszlYQAbelm++TwVRtkwuMR2WZTuT20d2aXaaYwEdbgI7ge88k1vX7bggz2J5dHyhTagmn7Wr3
pjFtpoPEly5/nRYOcsBAxLt9PC+RUqOBM0QVV768w1rueeKKSdLiyixFG7jJj4E0UzclVr3KZMVS
AHVeK6b2oeYD+4BsAUz3CeTK3FZRVQtn4Dtt+eXQCYKTlvsBVBZRquyDuoA1fAzTARHKZtNZ8BNn
0ehV5VQEl4kM/BZao1LNFmYD9EB1/xWBTyNIojCbi7OJ4GNuKeu4YpUbXo3IIKMZgpNUFDMui52n
vSSJt3yhEsc35I7MBAdEAMTICnrjS41aM8mRjMexpFlKqrlxFlsiV6V/U/W6xujmxSY/Mft5s+qj
J8uKuWTUyg22IW0tyeon/BnL32MXUurxvChpD2ctvGjwHoPUhmw0t1PvcEO+4jW57a9N3DTlEiS5
sHhHRUTyUhqjp4eLXlY5VelIbycy+VwO2nGk5XyiP8SplhCwUGer/gn3abgpvyEGPlBoL1XMXK07
+/MaktcWcpsdIJ5tsKYK1J/8VGQvEd7AH97cgRGNwzO8STmIHLu3mO5yqHulS/3yo0CMt0BN4DO2
Gf7p38ZTpdWThFP0qUp3a0XYJoQfH4NgUYHHse4F2iBvxRv88M6WKyTYvd3USLKna438hV+Mk0bz
FfsnZhK+x1IbueXuANWHso/kfW0mDr6Sh0HUCoiLPopCke9bksHN/2JwhvohNTIgsP1/QadC3Zf/
bdTxOLuQd8WzuV5cLknc3WXDFDomBtiQwXRtLWgkZauuybcDTyr/Jdc+nvg+Q1HHC9qmLFmzxaeP
TiqEOl6TSTrXWWpCH2aTpLq4O0bVmKyuEE76k9IQb5XrzvnoAEMf/fiPwVXoUH1LbY6IyKMikl4O
qorCdE24xmpE0Xa920K2sgDbLEEfrNMjmxfDuqhcVTV8Pjf5TE1g8WJEEb34o3jiVr2NbTuedyHG
6dvYtb+hSSL6WbqEwoA0G7dnl7/IDkWcUFXqlzZMeH1mMkSMNAvmFPnUBOT4CPO35Jh6cPgWdU92
wbdhcGaBc8Oj8cqApX4+xLp6WjrIvwS+dTGonyDRbPrBoC5i5pHWhUvlS3dZfzkLw/PQVCqtnxx2
svBc76yXlXmFwH4Hm+3Wtm73PmSG7XjzLJAhy6HPL8IVQFEVkAGS6sNF9Gmu3Jt5X6kHUkYDhR1Y
rAHptrRhxcTF3A3Pvv5WzzjHvpeIfCuhacNgqdRL8CQXhuYNQVFrD7XX6hUl1BuaHi68Mx+4BLrT
KgsJ58ElNE9zYlQiB5CSoobuDFDkpvT9kNJOdBTkK+jNBqBSyHwfH8hpkcE/W3uk6Rvl4uHR8G8q
yqZAdfWO99Asob8tuEgjUUhkZPHk4C6xlJJwmcE8uwVLfa6i2IdXKQEAGY6JqNe3xKOmRsY53Dad
42X8BpSKpc7EvqKkBn5cUSbxuH1XmSz9RU2PPMV7ib/Tt0NW1jynT0iuL+ZJIcY4Q7ldzbkYB4Mm
F6qK5UbNvx0V6yEdJD6cMuAts310v4cA58BKxOErBsbTnIBRAMfrCm0eP+1VoTClvd1oKnSTH3Cb
t7CI0DfXm1LeZfg2Z7qNVsYUeZiS4PZDZh3HNqe7BotOiHI/thOrU+L8h0s1ka3zxs1QFz4rmL2H
nemI39nx8R1KFZzm4hhp3/4RbwMFDDeGTHKQ8FxoXYc63qbGMsm5eemc86TZQCLakVV/7Wm6iI4B
ETRI5NRfWadg/joG8BNblqTcMPaG1zrnfDyyut88Iuw6kB7bACGhDrqC0VhZJ0+wGCnluiUBSMG5
qfnYjSVNpt4r9+VOQRxNqx5mJOSQtrVoyAH0EnkQpt5TtIunnUhyNvChcxYTby267fRlPAj3nCoN
gO+xrVPlo8niGcI0HM6TePv6gBzkV0pT+KiNydZfJr26TzqREODpiG9rH0BHTHHQU8hCTQIZGKow
fQt3mlwDxQ8/in0eBmGW2+Bu/5KkQHzXiDau8Os//Yj06iJuAy6SuHtxJFDGxUL1UAZ8l9g4VeZs
h4mSDXd/44rmr4QmUsDK8x4IxKDnQJwMzlfbc84t22uaUj0g2EpTEmC/Jd+h7CGqbpl4d7yCb5LS
xxRM/HR8Jy4i0XtThJzu4a1lolEmCh1J7v5uc5gdl5M8tqXL6/6vS6tInrVKFSbZGg6RUm2mysAp
lNiijgxOJE+A9qKgOoc2HVsa448iLWNE2ftf0YxtKdia3EQGFmQILwclOzsi7dEOHAC/ta8SKOSM
fHexHJjbEeloh/gqSdgEf2QtDbad3RBSLUxzryIxywwUZNvdXScq2c0OuwNLbUK44ut550t5BUrr
WbL5s/DL3kVuUhfjSNfXyUddp4K11LUt5q/6sH4L/idzAKpjvRxPXF97uwFlHhfklQMC5dixdIdu
/o9z9+/ynrFDfXp9wC33QMyuvMNqE/YrgUkgyFGkim+gW2INqt4OS4TQlkirjQ/XPD0lEftblNJu
gY+I4V2uOBQ1o9NPjPTHmSzKG7mJ15Xn8gpTzZd0KIj7NVAVaamJZXG4QjgPZXAgB4tt2wNwNC8R
qNyWrpsQPVHVzl67DUfNz13kcSJcPkGQUbwpvB79iFv50w16DfbD3K/Y++YKVprFL9uaqCiL/orl
0cTe4Fpbse/KW4zQqMg2iqZiIYOp0Fa4Xiw0g0zLGUjard27BThuhvt51EucDjKIyd6Qn3QgOQ/z
qDjyNvj/Li3lEk/7Mf5nPrjcSXZsfRIXdFCnt+BgljRRVuVyZ6Fv5UPifrKhoO6ZqA2+t6YVrn4O
0elfGZsbKMWXdiV7We6cKGqQrUle2KiTh6mZXhjZTMVFBlvdTKiBYy1CEY/cq3mlRz0wHsJSVEVL
JYcB6CXeqXclnhOh9Mj6DIl9P5gGnFrLyqMjGtfkVYgl2WjUxtO8lT2dknAR/JfQzquyIrOrxOoX
8r5jXmPY0jTA15JztT6+k49YS9rgHeXxfBQRqQ5EL/x2VL2dr61qAR4EAh99Rp9b8cYSMwxxFNxc
XPurD4vjCRIdBsec65HzjbNi8tI2ASUUx2cyLw0ar8yB9kwhrHkRqflWUXM6s04RWgy5clq1USB+
wWbzZyBNXPrAkeiI4arM/Hi6jCJop24LB9Ks2hXQSgM2rySl0a2IOvhxEsUdsgIf6mdU5zgxtiC4
Qmx6g0Vl/VkYSJO32RRePuwmvMAU+XAfcGFh/241fXFJEaSh73pwxhJLi2wBHdOL4Z+7HhoIRZLc
QNrnbD+KVKaTUMCB240+onZsU1vGIizdh3tyBEwGOpSyAYW7oUMbBGZhHbfZoTpREnC3I4Kvr076
SJLEMM1A9ykqv/U+qWojBiYSLdexFj2S32VjnKQI7jRR4FH/QEoIzXG0xg/FHVTcvoPBDEVKahr5
rn1fL4kTDDWvk92NoyK5zmjZCu79M1OnjcIfsgis1LM+mQwEO7rN8tKl3vOBxi+5W1vRb0sOM0/G
7AJuyCp2P2IQ6Mdwqze6fQ7le1QNvIQF2QHgzEFoFSp4KNkqQcLvSC9ZMPkvEEJR7ORJE8MlZOyS
efd3/THgBgcFPkZLPDbEOJalsfKZssAIIcJ9mlc6uWmUNdLw8ZQviwGDL3rnpS7wEZXoHDfrePXI
NTIcMHoDZKdLVSjldEzrgY6yNPLPM+oCqFjMmXKXFcn+dkQbSmkchVb6y8QCPtMILvs6kMATbhP/
6mSM3fJM5KAnUVBGyumZjcbbUDE1Or7nWSs0mXJgMCgUAvcj6yBKZmU2gaplGdk0DYUuTHi5XQOb
YsTjDLHDhkwG/LYMV5dxJd2QmQuky8gMF5fxRn8N64QuhQFP3UvZ8EQ04X7SB7HPT2m7vfMQ+pEW
1LLt39FAHUyKXp7qIpYrXhXNwWP6bvUWo5oXkG1aqf00bJcwSekjladDbIv4BmbOej/SAS7HZGXO
vTyYezyc3CufqU0SGbDy81NkVGSZNcbStUygAp/ZvXAIZymCvnwjDGK6y8jLBUToK23nE3hIvut9
OZqzmEZ57d9C409mcwTrivm9nmtxazkWFd1ouJNuEnoexQkLXmY5tW8yc2Js/c6M3RRaMxbIAMJN
HROlwPPNGx+r/Ft1wvS9P6wjylgcr92/W3nlKGz8IXjkcawqnmlPGeoOf4C05vyb9CssSQd6XMwV
A1X4LuXUghT+qRiVEEl+lPm+PBxgkszQVNjJrO7yyvKgoxzCIufUMrbpBlA4pBlHZamKfU9HZFO8
e+hK8eS3O1bVUVwejjKpRqJBhFuTkt8GAEOR5WC4qYO51G5m0eGu+Kt3Py2nxk05IWe6hLp8QXeH
eijkK6mDY3hWfFr5pPAG4B01qmrgDD+8ebsM9thmKJBzG6i5QqxEtspPj9dIJaJoyrLxAImtxy45
vi7qYJt9ciAo/j0HNmZZw7nMVA2ZWCpjcmtB7eUmhAbdKEHTokcki7W6o1gtJBLmKntKf8OZNhf4
n91hl4tyBfkw8/clXlWKO06vsy46II/WHWYg/geXuYj2NzCpQalTIQI3faGt7ksZluBV6Ds3eHjh
t+xaUZkDu2FcW8Az+IFlRfuxNytIEmFSm+jdyXPkGLAC8IOiZsGQp01IQ6YzSWdPIGThpw11Q+DL
dMdm0lamYDz0WAfSduw+Z614FP04guO9NgpsmkbHVhfxMe4iy340i9wJz7O2/jxO2UlhshkbANzL
ocuiqmPDbW2BUwYeAvAPBFv4k3GT2YnLFVemyUBawRCdxa5ARJaBMsm9ZGiEH7LjvALchrNuThsk
ru8Ohd2FKFDeeZDLfsJJujTUE8aAfrrVF00Xp2E7xW+V3el8uM0tSoMue6yypnEbQ7fbXQ0wQcYQ
AXEFzK0R/62DMm0XafUrnPstaoiG7p4B11ZVA08lYT5lsxSdXuhntR9659xC4iEkOOxbJm7G+fm7
QpbyCAyi4UNUPEdtqQ/h9gBNYvz1Dx6VTB+yb0YGWUPfyZUZXD3Oa17mhTD76du9sh7pJ9yOe86Z
KDT0l7AmIgkvWjz9/I9HsFDX4oY9cjYQWz8o07QxUtJPuqfbxW23DRZFNlx5LqQOGEWZHZLDudyq
6IW9sX0lq77SdIlIbUxk1QZsTbH31p6P0K3MhqaFJz/Q7FFcI4PDPgmeLGyDxrmoefMwKNWtyby7
CgGLr183/a2CvhQCOLrLqV4x6T3KiYNSgnEM+opdptZD1LhSL4ByAhPd2nDvNQYPpkePLCGe7N4m
PV9C4ZDo1ns+6zMW1U3Mcps+YeCY/esNcjQ0O6DrPCykq12QwYaXXu09Zo2IlWHByoHY0RiWYKIQ
pbto2/xBAsMylWr3aNxUeCZmxEEOIgRF6xhUrvaNG+23EKMQ3JI4X/X8A1iZ0RMy416kXo9J9GEi
z9eS2Vi93loamLMyfcRbRLJUuyuuoDRq0Irf/hedZ3s0QzVBl1p75ebykAPOi0Z6laPdZKHW8HrJ
Mdw+oFDLLALOKP2gL+7x1MDXXQj0Dc5c8jVgMGrsjqw074crslu8cIrpxWIwXQYvMZFFD6kLHXco
eCa1Vp33v9ORhTltlRpA9e6rjogvHq3AXxK7UxHlL9l/47CPbio5RYyq4xf0xOPR8KsqKo1aCoQG
uJDfQqNLQ0XoPRa3sxdATWX7rNPeRQH4gkjlgFFC+Fj8b/zGMCDkUMwNFlJe/X0ecFEg/C9UOunx
cjHpKrvMNw+/IytRRjtN1GYCLLpSHbztqLgT00bF7mR6JNnkB4gDbn6q5LHLiH3kn2vJD7E2zYG+
zw1mEGnPyN41s2mXCVrXfDbYVKA5VCrwpPaWwj3dsYcJqYAsTp0moV8xnkscZmhKhZpqV2Q8HoOu
ryhjmBnmOZhRdVGKFgd/Rjd+qvTQTY38NiP8JEdpsLooR6yST/Gfgg8G9CzjUezK3CE5hAl9Yc9X
Qp+7R0FraAdJw2Tv49vXsV5GXk/gUNEloIjzMGqtk2Vird4OxbIi4EKlPAdDDUBO+PZRyXq8pESa
Uh9OABaqsRAIYi5tjM5A8p+DowYsIPttfQNbIs5f3OaF5iYtl5pMNatCCT36Ejh7kbbhJL5Jn+xj
QQaS8MWGJGhUnOVV6oEvYJx/3E7wvfsaQjIPQNQnFpoXNyn/PGbDb7XCCz9M7rAE3jlxKrZkKXAs
ghwqQ2uskWrXFzaIewAiJtYfe6DEWZ/KqTCooPc4jwRwBfTNIaJEk5/aIZoKniC2IB8anu2JhxgI
DCktG78j/8QUPkgeYRcp2iMCr+aBNX6wJBWPndzg8naEgD/7930SyK5X6v79DinX5nU1YYreyhPn
yQdbrFHmib/2QMA7jEbBr3X4s5G8Serd1xha0djSbllc5rDvCqsKS43/LPWXFi4ZEYC/DcHmT+cX
yDThMokrgoO6KhkgiudZaIzilGKqqh4XGuaVhyZj2qKLiXPZoRBWy7Pqq3AHJ7tdaKx+NzNdosk2
EUqu3EWnJQN3mlLSa3lksSqXPuR7bLHECZnN6chbghDd2DpCHdcdDWQBQ7+UZEGlXzaTH6z/G+eZ
BWnaesPC5LHL+0FOsgyMn3uZjQ189pJWV+YRaMgzMQZj1YuFV4E2aTpOh+h/IWT0OPXO7naNfsse
M+o15QUlyfWiVB2AeKn+ySZwJksaufAR2QZpP7RygBdPsQ7+ZQ9UeYpGyRaxQY/UYEocoP+NUQkx
nh0Yp4xLxs1mi4yAggrl0nojKcPT6RIXmwRAVZ+4N83NvI/lj8tKmBD2qrb851QErrp8R+P3ot9R
8m5Tg36GY9XXBBXMZ76FddFRNfBfS1XU8AHsptA6pooh773mUv7jx42ToZXwoyc1LjJNLrOn/4tU
mrXk3nBh0KVUH1Zb7ag65nMexajvHG3cOeOU5FBc8T2GCnY8Ky7ToeqEqt7iCcDRZSlGQ3T2Vzp8
bOZ7spT77wwHH6JLmC8UnePZFxJ/srQFClxVuTKw2q0i3opXojqFA/D+Snb78TkFBo1wqVBN49bX
x4d1YSSNkdi/4np+zfVW3VgIczNXcX8WTPMI6V6gWKcq3J1WN/XxWHrTzltKEmeM6D9a6hM9dHdr
K2CgZaLcXm41b5Qv9ZK0xg4qRn3lCMSmKZ+wAEVFnW7PNfbjAQaTua9mYdbmzcBPSLfuvZz7zYAP
y5UjoFllAdHMof0sduUTGq+mQQRVPwRJ6Rg0bN5aYJ8WcbGNYVEKImG6V8+gK8V+5NuatPO+K+o2
Hc5n+GX3FstSgR97nqaNqF8btwpeQi0MRxRTIupoA9mCXRKDag5aB3h7mVlxOFVNEG1y8NlVm+G/
GoiB9MTLtHr0BAF/NArm36NUyZDaN6WxxGM4ev013+oOvqaI3XE3Qqt2gKiwr0AzAcWEMzdTr7p6
Wp5YXE8+CG7LnMIgKNZa4iWmcBQ0d3drTVMJ/uqpkcpjCci80oFBOpm17BCssJMIHnymbBPQPJTZ
4Bq+9Ak+RPvIbqmAvUsk0O24LvvBM8ndvVe1bfhl/QDYy74eiD9VDtsUNkTJDX85P0dsritYwSL7
jW3cYie18K24WPW5USlgfIWab6I7G15KIRZro8g+hUQere364BrQ5xLuZx1ltqIa0HZ8dh1MWaie
YzWVH8SCxSy6eV2uDnNguCkx7TU7OtqCbP5syazvOsacROvHlfx7DVzw+VWu9tG+O03o/Xtvt2r6
ZQ3mylVYQ75u/cnVdfu8rp5LGmQeIS30uAybC7rv7aGL1ikqylcGZ1KAKvTg8emvLNn1NTrKWM1x
dGJyZ1JZBB8h1RQxJ6aL9pn/FCVatztA5e9TAjzWVjp0Zqa/xxJX99x0YVDkhJBo6lclrVcBnuY4
mURthwmB521fZknUNLQh2bwfrnoaeag4h+5PywDyJl8wy9rCvOnqRr8Yj89MhRNd5+xlIucIWYKR
i2jjNvxULlxRPEKBVojPvdMvvSF/poFu/m5Ebdy1fSplvCVh4o6yzrqR3005kgyBwNlVgJ/ezNXy
OdzyUOjTxhjYpKyvcsxMpSOk6Tbec2VCp0rQV4/Qeqwx5gaCXQFxQ0y65fPqjt/sjitZ9mRezT/M
6dhmbAAKP8oWBGuR6a02UH8rH9wDQ66KSij/qXXAUrGFfrW9UQkxTrdL9Q80sbs01ZKT2RQlGRop
Eh2L8/Ni+wm2szeidsOtf53xUhLLhyjDzzYXdPGu9jDC22atxSC6V8JHAK/zD8nS6/MT3Rra+fWp
fzS66oQUfDowAQl2hgWLdUQO5SaRCA+p8p4PWxFY9831vsgSSHechJ53mXYm9IX+3sl1NX11OD4i
Zqk0U+UhCHkj1KWGdE+qbBOgnY8f9Ki1k+w/f5PVy/kK8rfvnN5R8Z6uJAsXPNvRi658E1OLibwr
LIt7Bdw3gvoCSPngsS4K/hIR1g/kT+1UlGDd7j3zFERuVzuTRfNwg3rEft1og+RuoX6G/PN1hYyB
fbo5eXKSdaUWvRrPqwti2hOyjS2wlQTcQw8LtkejZpqcnyaB2/Gp6olweezMR5nP1i0DiTgB42nY
36Cf/H259Jm/ZDXeUdlcRzvGkNFpjSceVxnt1zIxtKGpa/RPs97Mq6kO20HF/+/LRVpTLkDideER
/QzWU/M0pFyua26HRog7B/i+mT2qhxKFhkPTXvlbZOeVtRVOSHw2bjS0T1A8U+bk3ikA9H/99n54
2HSPM1FN78lhpIoOyWAWm84g/8p+NN+7UsSRD4aaW7rVlUVYRYOfjtRAo9XEIUigb6NBBYTAfsST
BehGwrbFK/6Frn6djmT0KoTZJFIrLN/lMK1DpRXE2MPesN6gb7Ext2ZanfNuAW+e0agQQcEMSeKq
46I5Flx+fr2LujBNEgkJEbgUJBz3RGs0sZt5fSaTYva4csMz79hmtbL/l5UNnQw1wyg/Go4rzIai
/jn6L7UWJ+PbcGxzXMb5xTioCwbDF8ADTyBxR1P6zQDg7n64R+ZIN/4X61P/EwC2dgWl4GxTXG6A
efyhAfqXlo8ZK9wZSMYxZFWT+ydIgHsx35L/Kox3H1zjhmdYPDBR71YYnMVWC1/lAEjj+7UisKSM
uW/F1as4geBWRAIpYlQ+TIKn7FfO2LW5cAS8cJA7fw7d4+3mikShl+42p+eLMmj/EInI3iWpo6rv
xnBmwge1c+iIxflWp/ztalu3La6ZtbEblQD01JNjoMWCAUxAn0XMomzBwW3pcPv8zD34gESxNbMJ
fRoZ2ogP8MaX8wcaYvxKSTr92U6NAT+UsYyCl3mw/KoEdLXehz34NA9b6plBVHhFMbJZm6VgGWrI
OlFkgupsDqHdfrKGiRxwmF77TvLDTcpzxVga79L4BLPwn+rRSmnhVFs9Y68IEvsQetl8T5CAmGJu
hCD/6HNvJrSi1IlVDmtnUUSiGNBHKgybYXFbFlMnDoq0t/BZnNOjAcH6z2OdtlnBQeWD/ojZ+Zfz
gtnIfnhISIUefEmgP8TpLCCQedkUhzcY2e76oQqI8w52K0REde0iy6whA/ZNrY2OOHdQU+X8d6hQ
m7WdsjbbknT02uxKbpwMqs+PlY02jGZ5ndNDQxCFGUxJ8TKsoSyHcB0ZuFg6tqkMmKnu2zzEb0OJ
iOVOvRcYp1rKwfxB2Ep7NZZW0rXcBZehKgISfkME5cFIohTBzoc31+SUbyQUi7j2YZi7Rsa8TFap
tIfXHGvKfQbE3J1s2+tmypRbrasmMwZjQypxOxxqr+AJchLsVBBcBAoIWlI466mc32C/oOEpQoAL
/JydXvVTNxiFmCdKiTItfKGOoi/+e5CHzXVCBFcWRj+ypxBh+NRXTs1RSuZ30XdmfqUVdSO8hIQM
0aYbdSp3zByG6VzjshhPnmb417eR1n99I5H+IdOfohMiQH00m/U1IpAoeVx2+F2xeWtTlDKaZVMj
4f+Y0/SMy6zpt6DlDc017euCwFP6Je1DK0QXfYbw5NZDPJ9jH+EqPRyXBOjrKDttIO2ejbtUFVgO
CIPQ1OHlGealUPsxpASR+pzJTy2TbiDUi95ZUuI8WvuSSClfpmShIxU0veGBoJrIaxmVXLCr9F8z
ZWTpaSQcigl/hNzRD8CPX6xBf3/3r93dpJhn6cgydgINHuqzEXHSSqTnHqOY+L46qBwdKZV7SBu/
HVn0g37NCGEBUtnDaY9cJjHMICbC38Fmqc5o1PTCVa0rLr0v4xcS5Zj03/xW5w1ZYAfJp1Fo68GU
/0yoQqoUBSySZX6BF772mGPgi65w4riyPGxC/xpmKH9jcqzOlfmOnTTGUvaUGYddn7ajmM09qHqD
iZ0RHCc4OKaJd9ghCS5ewq9VsKx1mZbGphBn+iDXkQGcQ6sDIOnNmWvZo19NLrMFtf6NEn6yX70X
rlW4xS9JS1gnLJbM3DPOr15UrISno8vS1ts67AWciSgii8EVeWM9v7Fs9i1wN8kR62qoxXDPbnn9
uPY6yk4BuWuHeoKACnMxmk/HNMOW1o73nER/vprsdOL3C1SXQnjYShQjZfrgFu5mVBcCeV89bqfJ
rvF+u3rCj/Vrg3R5cJ7Q8Xgy8ygdC5BHpEGDzorSp9XHgmBnHQmV+rf7IFsD7UgqVC4VyWk3Gv+7
j013nZo4g2WAzoAtcdP0cPNXKNy8eWMYoPRngrAvI9CDXzh1xZKqbYXkqddC5fgxbHvu4gSzCO+d
Je+sTf13amr1YsZmlq+OkeJuTXVo6nyx/GXirOWBelYiwlulVnuHBJ4Jgpx60VxsgPwloMR214zv
1XDXHxKFBxM2TCon/Y3wZj7K7dTd0w8SbBXUDRKXP5VgSZfBmLSi15XkSCSlMgOoSYpgXKbDsQlY
P0K+lRwVHUlPk67W6LzVnEdvkvq1cRn3Yo6ukZQkc2b63iIH79kepmp4x5ID3u2akgu/kToygynG
DfEB4y+HAcwY99sP5PvzqNAZG6LI//alEUS1WfgF0ngN5DUhpwOwLWtLelF/IDtC6PsnWJN0KSG1
cOuXCcxPtm+NBnSdfhayJL9uhSxo6YwyVsFZj96dsL5LRNbyXyU0ndH9bXSdm2aZ5eJ3XAt4wrTC
5CJTX6D9VkgKMgQU3oaOmFPWDN5iJM3+z0QZN5PLHaGXIK6RCTRSKEU8AQJ5RedW17vOKJrTtDwB
aY1AKy/RVynMvYXw8ECFmqqRD9spBnJiFWXFMf+1lIToia8+3Ht9lIvL32dGP6zDPTEeQ4JgxD/J
/y+Squ5KruFqHStDp7E3uzzcq+wmKAh0IwTwoaUoRjjNTL3cXqQbxYJ+nvV/uVwEgqGmwkrPfLUp
KP2IfEQw7/PYNTtJHAUsMRkl09Uf9V2KQBx2tlbLId01axvPDkHhfhQie1ylcJ9t597rubkDZVF3
Cqk6mEIVBRfmSCBpe/EzN5KrGTpWJ/TrRIh/VdxiwWlNKv6E7JZyHd4SgzyhT17FzAm82eiENTlN
y2mIc4zw14Yr3leKxB5TrtUPP1Ps62TWmkQWGZZ+Rxmlw3CTvC+uYbjs4d4aUlj7WAwRJ4vli6Up
0/3k/Sc1uRdxJ6Iqcml/CrZDJFF/Uamj6aankuyqGQfNueWhVPae4kj4yl1cut9kbI9/5iR6cWLi
UQTLrpwBAI23gYuxf4Aj3SmUjS9l3yoSGub/zUR78XbWyKf55tEyklTqYjy/RKmA+RervwUoKTmR
UoMvXLVJygK/CxKl8rSNHkusT+/sNVqV8jK0I6ZdjG4+4mtTBa2fJpcPPe7bL1FbjXPfbjFSPXwd
wSZ9RXm4yfuFoafZBCrNsm3JfDWDcXsO96pfhvE6JG8yBth2feCAFzgmtAD2z4T2Y92mYsChzJbV
YoMPpEvT23EpozO4h2XtHAORfXfgAoR1z4P06Az3qJYHrBDsVWYy58FWUzaTxKExhktkNiRIFLbw
hWc2YUMw7/FpIUaEhCaqZ8fC1u/Bq3ot26qPI6BhRUDgwrSP6NqAbCwi4h+vQCS+5fFLwX9jO3FU
BH78cgsGAsSJaF25frPK7xFphljWobKFmoAui9DG2ZRIg+aPkQHMyFv80nug5Z/vy4zNeIK8ny8M
32FSO+PxdTNSgNyRa5ePZs4GbbwMzvDYoiOxgIXAExBolgX5XbkIGX++U2s8KJvqqeR069YLDBYn
uB1wReR855rpY8QmnYkXD+HnqtgYm7gDRrV+by1jPTIiYxDaG0WrqGPwlmFw4f7yDwrvxp2TRmB5
ToZMVzfDymF/fCqvrDE9F2u8mmDZuZ2c5Wpu13+/FyczFpzIopabFIjU+TDFK/5wfPuykI/uC2hl
nvBTGzaXSvsy/INJ+SEAXsLmwdDUYrgvSSSDUZPP6CLt6C8rd+dieLSq3zGUZ+2qhGSbHrIPF1Im
6Gaa897U2Jt99IyPQBsJPx7Nrl/sPFRSg9fcUKAik34oJqEotTAtnFM9o1fkMrCyM/uq+eXTD+XO
gC+slMgkrGD+57bJvFFQKjQwtiRUMlrFeWLMkCuyKKEJEpDruhZHV1NBpCluOwMi+TqWt3qR+L9D
MvPC3x3mNe6rZBr5vKSBxhIhMdUHrj1OemKJtn3NHm9n/vPqRFm8fJso/526SQjWaNbl8lcGPu9q
vc+SlTGG0ppFq3jEHPOMGcOUkieXJqJSYgsuPuqH79SQjNZShhV365q41GPI1ykNfJkzUrLkz4Ho
Fmsr36jvL80S/YZGoeaTjWWwBEZtOeW001/i/Jku4nZ7yWCZGeSPPAFCBeYkdM058/efRBc8jkvS
CTjHhXRUuaUTSryTJ1f8Sn9hyyeVVLB1XEp1M6pcNu2Mh5Ol/A8vTqR+vk8XBgLT32dL2u6TPWeh
13rKo+BLzeuqgpW8NjK41EPbw12RHzu49CoeQDMnZqCqudJFqj74H+FZFJ6obULdFgIT7maqfT5U
jWA+zas4piYYfattP30FqrdKzYTglzt/B+ShT07Hy8ia+S6JhrzaREZGK+1vLkjxvZ90WjwU/Tys
a6ig7pZxo+KmevxH+pHl4PKmphuc6CNwHBTGf4tVW8784YL6+8ucABfIqdPkcedD8ywvr5iSydLu
tk5qxZCFnfXmVu9PDjYN0vn/475i+ZLbAz/oxN5OZrBBlweel25a5RVZH++5QaVsQpfkvMtI1Sx/
uwH4XF8FqgjRz95cv7u4jMZVLCVQeVlRBw9hbrp2l57jMrcYIlW15kkFuTzMvCjhJe/R1eexjf0N
VUbHTyI7nNOP4WaiQvVm5nu7qdrqNPAYI7u/CNbVpErwEama/onT6EaPtYzpB1AY6f9u8a9J33y+
j3ky7VDlt/tEiz8GRbHJ/74D2P6uLUctfD6C9WEKooj10lPcoBTFUVSg/JkgTmdrZq6npZs/xag7
MJCA6FCNjYfryZ/6rqNYhL4NDcCsfDF0nbJqGmmw3EZ0jR4a8lnCXAwbOkHCAhlqOmb673vsaNVZ
jVfnNfCTP/sN/agMtbCQmOaYRcYuFNoBTRQTciriROLdCwas/G8JRd9W0m4VOPHiFHFN7DLQqKL4
77AImt83PTwqtlwu2EggU/vcp3NTyucinSeqGcb+7PMGHnvQ78Ze99t3oPtQENas5TvW/s8rG6uP
XaGgxqhaaY0HGNU1bJiG2YwpQ2KX9eo5lELO3YUZRN1Pj21XAAwYcI5HIAOWsHEPsXVVWvadrj+2
z0CmZIoqhI43FQDjv8RFcmebc3Obz0koFPRUgqJiTHxVWAjppXmo7E0PjvAsKSeZZw5KAG3Qc/fO
vEHXI+CQVTp7bcAx7IfZ599B4i6TQ3qxu2Z0CAz3a1XOW2Tg3zAqYyA05LpxYKzFZWAbP+I6mwnv
TS3P4bf0JDGwAcPxk9AXzgE1rUHGjFzE9BfzY4omO01WFN1R1R6PCbwCskDmVNn/RJghjCBW+43B
UGvEnOg2oesdoHYqqtxsLFV2X1L82Hwh4EmiOBAhc9spP02pAWsvu6mcN/7o5O2tTKTlxrjvZgvy
+QMiocK4iBrlmpyLLUR6/nvRJr7NLVwBT/IJClvPOzrB81ZpU3xoM/6fKpB33EUmJKkkhX9haA+3
x9QZ8xnzDPOMv6Qh7UmmMXj4STHMk3bOhXBi98lDVt3QJOOluz9udTo8Q0PU+gApK6/8/SFnOzrN
zWPBrrYJn05+jaM0Q3EhoqCNRa1OXlZoI1F0DpnjVCTD06qIj085+/szq6MYRTTfF37TjHNLmCdD
KdPBMm4mZKtosguIHtEwgGTJtPz07mCygVzJeDW85xnbmGjR9AOrkqArTeESw5joHlXozgcFOIbi
KO7NF6VtsVK+VNw2wJp/OaIbhmUF1avJrPtAAncBqddYa982KeC+vtC4aA8ekG11dyFRoZvx1akd
vZtM5a0UZv/uVTtzBpwKoRI/I6T2FZpb6KhDFjAaTjY3P34FPMSSqZR6x3dgjIGe98vnbg+3oxJc
937WU84epxlf9kZwcUtqoU+h8SpKdiXdUcYYGbujon/W/N3KNyzxHykYsik/SbRmOV2XqUaCPlJ1
MC5gLNlnvFJ+591CaGUCeEhRFJmjCjRMAlOlvtPcU0ybQBZC2AqsYgZfrmvb6KaeAdwZn8LUwDYf
Ck4owhXT51Tkh+EVg/ieKwG0yuajFCl1e6U/Jhlq0rkcfaWU4F/Yehqx0v9U8IfB7MOM1TNn3mYZ
zkUBYQiH/yTGnMsOT5I8sE2ffx6QeC/7fiuYJJw2ZITXddfJVCiJxbnU9gXZVERzPkAJMWr1PO+n
pLbCOsRhH0LorZfN7lxbgdpHUNjtwSxwnTGZMouRJhJ7uyUgf1ZYV6UoWrI4SeElgZPO2n0wK8f6
+fXch1ql8GXkDWCcJee/pyHOfVanlzclr84xnhQqBbkPDcUKrRn/KTe+dH0ly9Swd/0wmD2d9atY
UE4qMyix8x8vOEPAi30cGryQQZx5MeWkOaFVMYumEBZCNHuQzZXb20l93dLE6ShGQiwMaYt5JlQP
6BgTPMMiBPdqVOrHdeqN9UG7wMTytP4RMKTninphHp+PDArW9D03kGmEiD8YnOCXwEuutPgeAaND
PWf+cxJAHwI6KnFddbfndt/uX8kDuBeF7IL3yGBtnEQ1iNYHZbrab+yydf/hZWENSuMMxRMjo2C7
ezE0gUMKY+6nbPMkORXDM63TaetDiaGuMgCAs5uGu2ZWghlpFSpoEphouFK5KudjeiYceOhDa/+o
M/eIIooId7gn4WM3FnBQ6yQ/JHAGuFvloXs/xVolAVy76nncplWLNq2qSPFlyHCRsNcHRJIQeJXX
T0/KjzCFLyGvdg8eKwBPR+Oaz14iOQTlR3fW/HRt/eiHnxfEpf/j3qWjKsb0gNKaOiPCgMFFDR6I
wXSE7vPzQpQ/th7lWq5l7Bp9yn/0KFenFbQzBpVSWBX14EQhcVhCNfaAJ58UD7awEXFWjt/Ojfu0
U9j7d7KonvcU0/fnyAv30+f1zQXaWcilR2br+egBBYCJQldqpjbH02Dhj7JqKoAABxvTtyJ7tv4W
YmyzM3E1Nc2Pn8/byPDycsGh1IBhHaqrOZ1mke/i3OX+YldRNoQgrJK1XP9Pl67z3q4uNZQkCaSA
zKvFxTQUrdBws3z6EeKVBQan6ujNqwrv3bSjlokkcu/gRTfl3IYkaVrdUjkGD4TUdVrh37tVWBUJ
Y9qJbgFRXgLtXFGO6BlLq5mZti4fY0uJ2QURo+kxEeUOR+YeVYeAXTOIcEPhnrOWgCTh660/DUhV
g+gBlLPzluWOEvGe/7/+FwyNJH5z2clLEg52zHlS2x7+sz3tEr22pDn+YXOZ1mOfn3U3wYTrqclT
wEAy712wON+s2gRA7ZRGAyPwDSaW1/vXcZicpphLn77y4WWXjbT+zl8qB6eVPTIDiYTvKRXBS/gw
e75n6FvFJZ1KLzm8iwmX2j9dmKlbHzZQKNdB3rHmE83d3CdMKdkyf1SlXcm/GrTKOvMlQ2HM1k1L
tWBPsg8lmUG6EKifAiLrfI33O34hmqwo4sQwFXmTtEF54XkWJZ4DVAfBF78dOPioBnfHZI9T1/JG
2Uh3X5DI/ONOxl0FPwkHbo0TIxnlOJCiYoDqKyzqlSBYysnl5l7sdZwqmjFvxxdw6j1mqfJJ9DpY
d80mdg4in3Mhdln+Pr0JA2mLo+8iPqrCxvdtG3U36DhlACcRtQoEjIFFfF0gwx+jGhdwSWGhxLH2
vEyr+IeMBzIM4rCDhcL6NPStgpwo5lDFKbiEYS8YqM48n9h74Y62YZM8rH3FpOFFWc9ERY6HzYM/
Exyp3Ll7Sfhjg+YEwdDwsaNW2kdXs39fA0JKk8+rwpTvFEQy6aggXWGSbzWpfF1lflJd7J2zH9eN
HdTY0AWLNZfpnHl+7+OatJRBNKU/YilUhu8HSMkO9NlzkTipSMRxwI7JNtgCTLqBLxfhrLiVCmKH
G3j+Y1Bnd12m8MAjWMkebRi++4BembI0bBMvP91+bk4xJ+XILZC8EsCjFwnv5avHt45bl8fJWPk1
OAsU70YDKiSUPj+OEUctVoJNuyVba+gEqG9wXYhF+HFKPFCRirL+2KkBB/32NeItO+QiqzBw1IEN
3toytU0efsJhav5KxVthNzUE8tiIwltz19H+T2GFmMnWSWPFsS8Ch7pKdU5aUG8nGLrtBG2t1rQu
7a/xAmIKbyVqEtSPzYSaK5wjI51mtyLznRp0Q4lg6apOwLH9p5d7nDia372ii/yZRhBOdMEeoWd1
XDOzOAnEsXFoiGg4jUdkP8wbemKos7UQGsegl5vZgx2HR0l23kOLdnykWktfb/1YoDcG+jpQxvsU
3ryfBJS964jnXZtOULXspNfFLP5Se2If8aDfW8KmZwoUPC8lab39VNHCSiNbMSjVPesGB19tDwEn
+kX2f/GzMAzd0GqGZB4pV5R9WBeIEhuVbyW1XWJ8MNpEhN5yhlta9KR891c0pX/kYMbenq58j1n2
p2X7K9+ZM1uXm8HW45hmOvnpt7q8ML19RvAXHZhQbu1NRaa2QpKeyVXz3BHxqVaZ5n3MRUNkBAAw
YLAPg2Iz20JvGEdWUwFk7f7qir8Cg/vC5E2LcAw/W9sRb1EkhFhbfm5Bu2RdPGoRjpZF+qs/8UGn
8gInDR8oB3AD+GTOli4+FGNsEFuIPVonauGE0iw0vcLuH7CoSMS55A6McgPuNC8te7b82/u59ZRB
/Fxfw4RuaZlPkcWWVIFyuF5Y4C8I+TusEbFBmsaoefw2VpyhWI31ZKOubenoBf8mapf3rpGdc1YB
D3ZqTZ8KGeANioACZTSF0E6yKEFTcF/xzClta/Dmn9bly0d18G2Ed6JGQACK/lQPjzUYWG9hNLSP
WaJmCfkxSL0sOYB8kNr33Hq9Jx1LtIJp91ext5MUwOZntOfdHUC1pAZzPvRt1PYxdCceQXjERPgJ
DASDmGsG22tAwwudOiK4p95F8uBULtQqMve47eJX0DhfGyutvJcrz2Rl+LLthHddnIIOqUfBDKKB
qmfSGzcpAyjhLUStAo3J/aqs6l5YLDCUmlzRcNbjwZhQudMBIIAm5q7wWk4ivm+y1TeNUWPOykc6
bA+UDktxjtnpsTuPrbgAE+Zq01PfogCRzeJR2t+RvMrCQNRbsSQbLCGHyNewSezjMM/UT/BnVc0/
NWD35PkmFc3vrfuyBYKXUBtlarUrI3PUBeQY41HZ/AcXMrUHfJK2qfUEbL/Skj7ZHUwxi15lZIxN
3yw3mrOg8gNqtuTxqighMN+wBASYNJiWOBz4h1jGq7Qq1w/+lFNlpQmUm/GTt4EyAf6r9bkRkq8z
CRVEAZjo3wD4HenudO7j1So5el9azZpKv4vI2ysPqM6mzbk3VsYvhazc46k58oCQRjsp04MUYIF6
tW5bQqDBKLUSGflpipXS/JvRoRJz8QY7EhGDC5G9BhgH8oUi26wMR3Ik8cnlqBEONMkV/vfkaomx
fgTEfgn7WyblYsTo+EZQz+oaOdPkBbayaQIHFff6J0SWmZQeNEOALlxO2lxqRephYDE2d3cqA5wG
akCRyaDsMvd+CI6dMlR/Mc7xnGQgPlxSPNtCJqKTMRcxqqlkSwRbzlZtQQdwWiv6n3ocJ6lexxd7
GeDL2nrwyQdka85WYcPgT+ZOCcHgTY9Rd79uc03k+2GiDWTnjoV7rlsfHTzfhRhnANL9TaZRE4zO
ylcqYfY1dScxRndNCrGdpRMetbLINXINAIkz/AcIRNK29Lu/MBirHekcP08V2cHFvOmoqIDGlenQ
ZYzBUd7rk0GKh8pnapLFpuYCBR1ixEiwrK/WZs0TjG9E11ZAiC6+2mOJLE/hwOOd9WZvb6bYiBJT
yCVTwTLuMonlYPmOZsMOGNo40nSLuJkIzopGDiru++X1j5Ukn0ufL4qcqIPFgU0ejlmJJuOC7wYo
S3B+xh+xE8SdkeXEQuTVkjKDnLahJwE/NuRs6fIFWiepPrG2mW/vnv6BRGcjB1JfnxiC988mWBd9
aaa7j49tOLMNrA1sHUlf624aWzfLWRuT9VI9Lv0lEG9SW+LTqmmJ8m84JJsxp03W6nzuSJiFPsWF
abQrwBaPW2ZUuiGlt6Dv0QYPfVRfYRzn4yff6KY6o5jFdy6iyBgDHr9YcGpVR576SbdrIe+A/yI2
Kw6v6cEgr2BPTw4H5o7WzlWoUzLB8uepxoBCvOeGY0GkCdC5Ktqq/Xi2r4orFUfarBQunXUdo2Ue
wjVfr88u2k88T51pXXRyWb14PLt81FFArduwEy+9sIVzp1eS/CJoqgFUXuxrtOwIeRGDNzhmPAAT
zc4CvANXx1yvAsoXiNAo68STZ7vrBKelT/SST7OzvcnZ7uxfOwCftKn07BDtZ8YRq6fBMbW/kY7x
hfJihJedl16M51FMamsN49BdxlX9Zt1wAnbT97gjXlHNUAll8nrm1tJydo62LlSkPcJhVWCiMfdt
U9eFOD4jh1c5R2/Oej1znCt78Ta3eM6Uce/G2rXF+Rrw9W2s1odXPVITz/p3W91UaxOkCVvEwI+x
bWbYps1VwbjfQMWzu/HRU7uGSHHiqBhTtWnramYaWb9BTc+Y16lGeAYsDGFrDCwKHB8Go7WzQDzN
UyCiyqwwTAv2tmaH5SqK9ERE5cImfj7yHesula608XT7+K0tHj5kv/bWtL5CXKiJsW+EUkQogP7m
eLeIOVoM4Z+fOUfrT8I5ee6JC2uXU9ACSVXoY21SEGv8mse/S1X9/1my7SpDBm0GeNltYzykm6Qh
9fy5oBD31KxWRJvBzXuYKy4hPyawGbdYdcWgYZZjYzxi7QPgRIRKEjU1dBbzMQk4HJh0mTsZNsBZ
SmwqnUugvcyM4ZM5qf0jUP01BD4eFEaAB84dndLsYKQ5w61HxqZbc/LWFP3c6AycOOXyekM5ZTJP
9Ym8JS7j0excCy66YnYfpi+kR4cfGyA1m3s6iGlwYnSwfN7Q67MGKYQ0dONlk7saS7upGpATXxHi
QIje3DMRFbpkBh+myCoK1Z1056p7qLbYWvHEzwpfjjAuBL1sTBZRDv5LzAIfCLCV0HQrgbIQqGZu
Ze+l6Jz0FvM/bv7Kc9dNbsBsauMjWMx4kCD0WZ9l89dz/cckHDgKRJni6ufB6mj8RIy9ayK1sXqS
0AbqWgn/fy/O9/turzzyCpiMH6kQc5NulLOUXKrZGoG+2oZrFVamUahwwF4XZV5ceFUweGVWvBjR
arn5eL5F4oIPhpESEYv9og7fty1rfgAaGh5rmJfyT1j//wDLPFtgKtjUdRTdoaBbkWL0AI5AHufA
pzq1I6XtfUMyL46zXKwCxraRrLOTmw4REE322fFrvC/BTB+GKFcnDgjyjPyWpYJmGcqqtMhhsvNn
MdymhgB9ZnFdZsW2yqpDK7/Ws0PWtyovrVohFtmykGaSC2mvhjvhY7YBGA3KE+igbXsD+QN10KJg
1NyEanq7CQuzGcoxMNpcUhecr9uBBH67uvpCyrEq7My6NVFchaw13f7T4jgHV818itlfmubvU6Y7
Aln0aLXXhTwAzMXrHYt3JuZU2FvTDoi19yrXQiIKRnBfqvwHZL8J24jxBXM1KN9Pj422kr1sYTTh
RDlCiDDnOPlYeG+Bi7Kl0gf50lhs8uKRMoUfy2YJMN0mNEquHQ6o/2HPIsm4eg0mJ3PHIC5mSuNb
U6N9xwRS8qLM/0NwcByJ+WZToOceQ52LXpH6t9EMmBB2i1JDb3teVShivn/2jZpKhQ0rPT81dFJi
MsACf8ITmkfn+843U+uPOlxlkzsJ6aP9ldKz2r8GQy/+UL/Ronvlpr4NDtv2HmCA+DCWXTapaQRx
vXIySuXWatsvLtQ3atyhEsRIzd90aKO5EAfHG8gTLYTW5zuLaKy3AAM8lxgYIHvwx0SoUTBiLk6j
NzMiMTJFAOihvvi+FHWwH1hYdtok539FZCBF+wMcyLmggDA43NLU7JAKU6Z31A96Vck2cGD+sKGz
xMlbLwMUTWBECUr5YzXaCgX3MWawYeZPSt7PNrxjbON2pzRNxYQUXZFTy4pTx/JfJLI7J/fkuPPm
HfluO3E9bY76MQgcnPhJXszLUJ7EqL0MRnh2fZDnAy021J5l4vvQCt7QmGikiEZ6/WiKlgPqAK9w
Y7w+5THS4lqvFcqiVjHiNeoj6b0Rw80BeN+Nds8lgAAmn/yUynRDlkD/APhBGfcppbS67q0DwNsD
wl0DaQ6A8rl5wt58hFJTLJzSS29nLZ/1MyHCGC8pAHeZN/wfsQb83douvrhkyOMKVZRIm/bW2j+K
c0jonnkYItLdC5qo3doCiLq4mcD1oRn/UbdzmLZOgPCAXq7KhHbRKG01O+XZZ7Nf/xObpZaEdCOY
VQ+5wjG2Jjh232ykCrqDEKpRVvkGL+OU3LG9yX24eAQoINyL0cplWgySwpcSDUGvAhmbzZa0Ev+v
9chH0CFQFYMvEmpb57FQn3/aJfnArQnIlJxNBij2tMo2BFQMyrk5B/nrxFe4E4sGNFvvOWf2zzgt
d42+LW/K1PTF3d76l/cBFnLuJK0W5LylvdQsPCFdW8QWk4XZF7gZCvVnJdWZn//r5fUaLyOx4R8P
AM/MObtxDwa9PVcCWk816dts/5ovVlqDNnqmpJYwCw56uBtZDeA2gUT+8ZRS6Haxm1ZdiJsU05gh
iHmwAbbM2xAIh+XCGEx/br0Uv296oI6vpI74PDh+HMdGsdpCD+HEEjKG0+ZouLDCELVIE+QygeZN
lwZLceDXsh5IFblUdq4EewzT7GpJ9ShI5MOtKjk9nUFDK0X4OnmkEKjOPEdsUzoHIlEFdwNnHyRq
B8GhE9w2F2fD4XxBYDJXtGbejwhM/vx+cfU+81cl70KyZqNc8FuvZg3RzD5TEmPCA2G5t4Ncw6HF
k/QdcTXeEwheCHaivtKq05sq9qoNsZvAFzsRr/q4lBUy5IYtXtoyktEbYAo2sBdMnMbtF3r3TlZZ
wSfn475Qhxl9V1Bb+4JM2aL0V7vjxayX2+1BY41SyGTSxw5iqDoBKUptnfn/SiNLFTTkI9zDz5dd
kB5BON2kQza6/7KKeBOPvcoUWrxVJcXv45WkFwlK9200iNaJjWJ0GiXb5c2YQiROw/ZeUYRMyRSo
DiEzV9y3kNZqmbcF58DWju7fAdWC4ZhdzU/Y5UQrPjnIgJmpNOfWOOy3Bpk4m9OjXPyN6jryz1W+
mQ+CZ0d9YAusPtLtl17hA7EgHhv2blqw95bAEOUOp4GLYHIgKPm90ctabMaW6e8tP2pI+LPzb5kc
0WI12AW9RE+7lVt8spvqZutoVbi8MxbGovDd3ymS0/4/C7lLv+uCl14yN7LLOlse/H1SW5cGJ7S7
rsGHVZqm54EsGfUChvFf6iEhRy2xnEizgGz03pMrVvW1NU1CdNTVtOZtXOdT18WYR8JHA0cRUDD0
CHRmscR0EFVsHgdtiPrI3mu0tLWTejX7eeUoDll/njTQRaOSICJORAwqEEQ7ODVb1dodNcZFNJM2
Ws9ZZrWmbihx7JkzJHUwamGjYAWuYWv6ppMQYjD0mvDfNxbYoaFWNFkdirDectypFp6apbmifovg
Wz3qoQVlO54I5Pe/phwNmJjmRH8wvznGp79yUoQP20fNcxY/3wxqsfGIaUEQ1kE1j6Mp/BFvHO06
u16zq9vplU7FrfHdmaRP0uJQm2Pa6UD6vNLhFuRt7Jm/9WK67rGPHvYqmqqRYKaDpa+1yhHNxwuI
R98UuzGFTETU/gUrPMdH4TksOeFBdck8w9shJvoAgBRBWZVfnryMFSHNe/ZMf7w+TX0MLqOBWvhf
NGiczgtnqzRudVrmDxZntboyzilprmUglafi4bf+L8NVW5QCVsPrm2akljq/oKNZwfsLjfdEv0nU
sO8dj9TDyJmbPBU/NXnozIJ2YIx92gkdyd0h/XxbIlWZY+Q3RvkNJ/tdxxvTKvBElYpdtN2aXvrL
N8RYzeXfxzTtwq0SkD+IS6NCHizrOx5wfNt2qq8C7qJfNusq2s6E97C5nVQDFDXT0dnAbTUY5YF4
n+o2/HboI1EBlrukwjp9QRIFChIu6FhSK5f6Ub9vSjL5HrP9eCone05i3jh2hweCEElD1eQwhm2p
HeMdMHDGWEoINSwXsujkn+HptOmoeY5vKQiEGMEuslkm81/kmXXaWXj5A628i4lkHY3j0gQkx62b
2V8RuzV1wQnUV+TLd66ISmehCFkoecMjEH3gRiTH6rgc3SfWOTz2kzdUc3rA2dShxfeO7oWzjG6x
Y6h1LWNlvZflT5ML/q46mqebw4gI07hxMHLLe8NKuZZUL+cDPGXdEV3Fdk3qTSeJz+kQzKf1g/dD
GV0wPqWRlc5nilPlv7RobiOustCUZmjrKAyDDM7j4sVCAJ/idWA5Y+UzSsdPtYJi58iZJxsrrlh/
9Nxi/CPUMBRsBX5/q6C75Pc3z5wfpP4MMRX+WlFbaDgGcxo92LKvY4ePhGsduSFAAwtrL65dFpmo
+QL2RUegzK0liC2R2O8wk/6uZSFPmGJWSihn1QG5u9yhuthdLD31zma6G1KaG/fG8uXmIm0iqBS8
eRsMZc+iy6gh35Dbq4yF346l6q0COZAExNBpiZpkjj+oECBnRxtk2JndRmZfiJ+We///pOMy7zAg
My0aDaFMhqGRUah4UPBV5ZzSquh1nm8y9IVh+KIKqxGmVwxBHKj3N5vHYWU831BTIrey/Ja8QcVS
NChNkyki2bxobjptMhuQAaQ8sv9PuOMejqcVv61MjcRfYL/oBSy6cFrFH6PICwhl3m10LceBgtkw
2QZzbAMHSdnqWvKgECpCN6rwv5WwjKx8/hNRU0Np6GirPEGz/pxruIR0W5rrFb/JCziG38AfEI5t
8VYDrAlBhWqc1cBvPPQRqtMx6u1EUBZ9iMnAWTxlZsNsuv5Jqdj/pifi5nTcVbJ2yjoPGc0KYhXD
Yv4quCODIcglr8S2wgt6qXdj2lPw6kwk5bDT2TY05qI3D0rlaj8O3HL3i8XO5dcUAw44NgApHfmX
7A26tlnfxCjMP6E5LYs09+09HPyVE6daUYI9hIdV+jGB9bImec5gL7tQWIzYKCTT1Wl6bpNGtFrc
hONMOZ/VhhP2lyvlAyGd5htxYzkkLFxmwkFZPwrwbvele6Woj6e9TwdNa5O+Jozt3akmdbZBMMJk
MVo3U/gUctzoXkhRIaBGZk+RfGTpwcJo1qlvgj+E9bDCO6r2pgQqVeSdLIEtldu6rubnQ9esDPNr
Ys8/yMZFywAcJHEBdqJTQabBIvM/O43S7fK56DD19rz/U4oPWHx2PSATeOcKE+l6Rg/zsUJjV2pt
f6WZ1dpjnNF7ztFqFOUkiHohQj76v7oFbjqs4ygTr11pt8omsd4BXddhbQ+1vraceJHaBSN3IZ6b
zZDs2zFJ2drNZZcosoPBTQsbZQeuZ4588llRhQkdh/BfzPY38iwZOd4H+1FBfgZlbh9bgkV5RBhX
/PurC8vdRjEqlt3kdIn0A/YEorBmrAW4xiWS1wdGXs/moWSg7WcQDyd4Ce7zUUaDu1PuR+OU6JYq
jbGcS1RCXGG89GYQqbCWoE6W2P/GrtgStVLuV2JZFlQGr3qnH71xxawRQ9JhwhPEsjR1Rzn08BAm
4jvni0wZf0u0RebaKvZb2l+y0a3DwUKz+VJeNAl8si/BTt3EAi6GQbfzHbsRY4yKUMeyoz519By2
jd7TxXYqhxl40CS9WGS0hSkqyKdI20A+5YeNVLs7nyRq6+Q2p1pYnRSAAYx6uCPbmIbfKNyXmcTn
pJm9lMhhgDtUHKgJhjMyChHHrILA1CmgA3+OtbjiT0oxJNBRw0B3uNC0IhEWgWYsXdnzsdz5OzVr
MGIV6Kn9HY4cQ+SIXqoQVC/+PCKFKAUW25Qn64zNUGTtvaUQYNb81CHbA7eclB0BhVHL3VuYdoi9
1Dz1PYrQNtSFkgt4H8gJAXLONBkFCFjaUAQcXCmuvg2+GyFW1L0L733rz38jDgSC1k6PH8pS/yO3
wROOfX5qOXxE83N0rfWwLFNCNeg31bwBh+uwSdAMi77CrBGKTHcuFnJcFu5OsKo0Ytj/4KBadK/z
aHdBmgSYaJg1vwt880czjbfSOb2DeKdLLEoUrAtuI2QyCfUlxikw1cpQCJ0RneeSY1hSeFhXd0b0
sNdLCpl1H+7wiMgwY1kHOo+qQbzpyvmaHDPTWZi0F9R5S1o3+LuKPQGNnj/dlZOju/rPf0apnphD
NEZEBij99KJsGgdEz6CkcE0FD+vtd6xmYuBq4+o0+sYhso9QW5Ju46qZ1CGZD9rFG0t77TAQWtd9
iC86ArXdxwbEaV9FlsldMNmswsTxsxT9noo13itTzX71cG+98lJDLxo1+SB0AAlTkFYD8K+klV9R
KcvpWfM+R5SHGWeYqwHu/s7YV3D6MBHozC4pYUd8E+eWrPqwicFoDsdE2a4XYGikNrkyyv/7vx05
0QVkmz2D7dO8ztoVcLrKD567JWwrCo018BkiDT7d8qxEWHSy1YLe4Sh/mlwS98x/0E24z91ToSS4
s+VitGlJ92onECuFzF5WfWiGnjFrZZcYxS05sOn0K7Ybiqed462JYjYYHq10x8t8jEevzMXyrlsH
b50jW1Szn1H3BkoAGjN+BzQrYhc/kZPQ6MNn0jcTiuY+CWTqLYd9wHAW4Mgj9TGVuR9vBoj+vazs
xe+0JUKZ/kOnsh8crAZmVIfJqKCZuf4/pFoJEBfxcq+GUfR+ifUG3Zm+EAJyy1BN1RtrLS1YdUPs
IuwMrcxEATFKG972NnaemWmgIorGIF5bzehoJccw3oy0XQLm28EUfFz3AQPcM41yXNqfNtHwTWWe
yE8ExcSySr3fqriB4SzJRgWDypgV5Yf0OT5hCN+P9URwS1yr5Jlh9YAnLlzYSFyk6Kse9h7J5Pxs
REzzW9gXx3HNr2833MMgM1On5YRawo7tyj6ZEUeErOCjsrO0+pn6b7sPCuQD1MxXTyaDFJWa1czX
tn3GBFvShD/I8dBcAbwF9CKys9jsHkmnZGX7m2nYGVmOyk/u38kG1wdKSbssQ3/7V0jtWTmiuBsE
dPGGPQdr83+ZkI0i7+AJenLxpZkWzQGbIvyXMpJDeoOZZfKcxytGaYWv+h6RFKyPii8mHnXO7gB8
MOcRXqyQOhrfAhWdOn6dDsw7v5of4E2wlSnQR1tqG07bgqvjBNTnSUGhRK6V8hItc9U4767CpsbX
L+7HfwSmuRqEqKgmGdJByx7bVZS5Nju0H28EFtvuDctilnZ/DwrQkukUgoY4zS+RiF7c1U+E7cOI
MuvAnfdgJDckFS3/95WPtAOB83KQAzYwkiiNpjGugQeUeR5Fr8OoReczqSkUJFoT+B0BkQzqls/H
AEelVjX7GhBXgHt5vEfo3qpFAAMIlfG68Nn/DerYx2HD9M94+7oQY8UT+kGJsJ9pWjIZl24vzQmb
CYupzJWbXdWQyqUa4kw6OexZYg0P8jv24FMOXVU0Alyra3mD9Ydr9V5LskvRjjyj97+vhv7wkAMk
tL+l58b6ccQ+viA6x0Z5LCw319tFvPrnj29p5EtPyD1pA2TrzCJMrkU2ObfgTZq600Z7QxR2xVWn
5uV/2YlxLKwyfJ0EwXv9FVWvP45dN5xeuqDEG1NLdpGPqh1/FqFBv2br9W0U2u5XPGS2U8FvKo6M
waW2lsUbWp4O4sM37PRsk1Ji/uvLgeDoYjkDO/AbStgM/Z9QFQdmQazLsCDFI066J1zyCA5oUFSR
kbMXVOdFQS1Ms80rOz6CYbkQk93AulWbrFBGm2xsrEwekqnYFcALhE/feY7MqT610MApPxjWG5EF
y/w5zt+JAVtu/FPteuvnxENowJh73GzHU657jnjgTdn5ExOSJ8JSN0T4ejfaeSioo5aUsTp/MBh+
sqxWhK40Tgj3GDAmh580Rh/8QCgZbtLksmxmw8MdPA8m/xA6ee8ocsK/Hvkb30vIxzW0ut4w/4cP
m5NF4QbxSDFSIhiwi237fR2ky4OfGh+5Z6L6PhAOCQNcSc0bTKod6n8FjmzQyoig6OZcPzhvDhVy
ScB8OoGyvQZGdowk2NyjYdvv5JD7hKySO0guUAYEPSjuWdg1GU1dtaDxEDbdkVlYjNE3gZ2Jd5ZY
pxNjWSaiTN/GibtqQaW62etgMtJhh4EXv0I1LaE+v9rOH9B03C77JsMGeE/IWUETeDAy3q+WFJYx
qF9CupJ2WeqM8tKFb8sUAUF4Rha0qLEmgxRqLZ60aFnbzRWfsGfl+JlgEwM19oYogcxk6MsNhrL4
HPvVGVrd60HPYDKMxl9d2ooAUHADPH1CwuSOsA6LJe8GL7gMGG55UONivJi5mokb2CRPy0I/uI/v
F5LWAEtMb05A+DHFSK4or8EFU241fX5sejy+NL6OGwPQpNaOqpygB1j51Y8+S79szNdV1vE2OaQA
AToE/3BdOtoJhEXxDQNv9NVYbmcxIsGUCWWsMVVOCuVkwgFv6UMvHLMhggFrRz4dc1SQELyP7ZQn
6jhCHKIhIfS5n41XHQ8XCKYA43HFlJsgPEOz3/elFZ8wMPnjq7ngNAcuxEtvlhWiDw6mEiqCZP73
sOd0hQNUJ+emkDAHaj20g/1mYe2ecavrRXXluaJcK3Dk4I2H9GfTMmB4ZOo08PTOwAQw11h3e5uc
R3GXWIXhytNHqOTQKyiFf79/qNWRHCKc86zyBJWhiT4CdCZ6WZkGBSRTRwnqKKkJ1A4A2Fcy0CvB
LPVUPhj8coGpivSwRPnNvoVpy+lF2pp05I275byIHoWVxZul3yldHRc4OELvm0yUSzYb/n47/QcE
kd2hgtHNQH0a6mKuMPirzF3MDJ+i8MT9rJo46PCXhC1bUI9+WTUSqlgkxqLryH08xQbx+l5bJp4E
4GFdLOCcS5EldX6IaX7LXmgDGmZvcOF/DVeXYQkBxmJW7NDj/+B26zt/9/DayFOuIWP3TdA6R0sk
W1VU09yPkQBWwfNodpzV3P7Dam0uMHdzpEJ6c5qtlqFLpoqVxOdFSUBmohy+Qqz0rZ6KRyeo+ov7
bR4/8RLHhayLxbG/TR6CwgPLmrSFtAKY8s11kP7DsDWJ+8fMnoxa/4XBjtTg2XxLRao/Cclgtp6G
mt4ZeUy5aQZFl4gVCO3RJPvreQMhjF9c7MJJBJY5A5QKZM2ClfZ6kOIl3zQqecOo0quzfPkwHHFX
X6Movtx4IgB2oRmb4PnIi7vz/7y+IX7YmDYtuZVsDnuf7sdMENrRISrfjCwAQphP+j3vh/lnsNoI
vYbLOkfuqY+KMD9V0GwpbI+kUz2U/CnVNW3Lkj4cPgFFO1bhF3iw/QMrzRxzJtXdCnUdXPSg3sbm
YxcPA6yEeJGafuC87bq9vD1Hjq6o89J8y6Wjs0dCsMxOCiA8IZbKkgDPXic55EUdnV0QsOC3l/xR
28Zap7S3mg15gDlGYjajbkFCjjDrkg5LQYbCkydLpXm0abnjyIaRQZy8mwVHZp9yhtbfFwd9tnu7
tFlsWzxiD9Cw904R+O07Lnjal1dzCgqoZClMS8duLPixezyjrU2DMWSL9yxb5pG1jUMLn7ASXBb6
RMWfDHu8i27Y3MNrTqOESKUbl9ZfoLl/OYqfxBCZL3OQFOeGqal4C1QZxf47xOWiLPpeEmw/4NoW
xgrkkTsNpVF+8QgsDuU2LL1vwdCT24Fl2LiMZP9i6Fn2RZkdYNfrOMQBpyycP8BZ8bhxNFdJ4Eik
sTSZMU9TN7vrP7uM27S2p6M1yAtMVLOy52T05UBp2nW0dCvxdrFg+6Sc5cHKY0/lOVjCOcpIEiBL
rAfhagGNl5rZPvqjU6+C8JxrcLwp+8i8mbJR76sLmI0lbu4U+q/C1o0wQer+WhARtNkCPVg1XpBf
4iTKr+ymsS6pJmn0kj3zjmWfLGi1YQOngunDnees6LEQ9MWX0/s9XnQs1u5QmZ1CrAwfp24l64+G
3zaMaAWXBliHMsIvn76m9LS+gVBDBDqUVkL11K/QifzgFhOF7Y2vwcLQ3BGnVeQZqpiIQfhY0quA
dBG35a+ZYXIHpgDka2YBnW9n8fVVYe4CGipHis//XbdIjP0tLXwQOuL0ECAbizlCQOkI70h1oy7U
7y0yV5G61BGKke71SDE11cJ+er/L4rkpD9zF394xxBdLLUrU3M0MDcirpqw9VGFWXYDTC4LtmEqc
IH1KfpHLHfv8vfYA5ZZh/2oSMtbRKn6uP768Tr9oS0Ri1tNThs4+RaG/pEQljU7HaQSng4Pdo6RN
EDLSHEKU9UtT0cebaiy3s67N5S0wjEUl2mvqke2HIrNeQuHJ5+YeQz9Owz++rRxJCQMFdQzAV4BK
KR2rc8vQhaTklRhntOtPCJx69Ef4LNVDc5HPlllagDRXcRViwOqwlAeGLAHZ2tiQ6InHQ4BXbior
8zFHeK7mcSMnlim6S6aj28g6vabjubGTyDkCD7j5XNFaRqhiX8aX1ERju/ClIPdI98GdwSVhv0hw
OWir6GiUBa/es6HECCs+7HN/T2qO5HaiXSkYsY/+Rglf2EQ95ElezkjqWbroninO08bAI+vXQIHM
S4hp31Jf6ZMitWFNN2ywSUjDTfCleO6ZID6x9FtW6xBVcJ/oFnZTqtb/LiDt2ewzFJA+Irs9yqZU
q2NIwir9hZC/WscFINjjmdaGYDBWakCMS72FSetB1JU+FxTJrd9mu79gy/MxP5qi3Ay9oBa2r9At
mHg+GevCxXfYrC6FlssKLtJUoEXuPoPZlU7taTdGOmIzByA6ZqKdDz6cXukKYYi6tTG7wjJK3Med
KmNJ+2x23XyTDmS3Cae2drXsa1WjztTb+p/BuUBUbZXoH6Oypf/5jM4XRKaQ/krCUrcVhWnx7xM3
dLCEohIM3K3RFYE10i/qI9e/ABLtPqOrk42mJMvGQ0BHmLZ6PmEMVy8pMG98dOz/MFzq8wryW8+U
Pz67zlj9Qwi03adLhfzkTD7/LkmUrGcV/TtzgubPA7U+gmHPmiAxxGjGcTu7tlrxWH0J7yZ6/FFt
lhJCEdBBjFdt7HqEMklni0a7d7uJMTdNaTEoCVy5J8/5S4h4yVI4SlsUe4a1hYFri2DiVMiWmkZD
vjSxokOPPCSscIzxTQ5cge306NlzehIbeev4EFXcXJzLQVED2HaV6QATtUj+2hdXQn5OlLzuQIzU
kWdyB3+P+2m+VkupWMeaU+au+HtL3cOfdfgzlOzmw9q2oQjkMfei/BRW9D+kDfGyGFohFVWFzeWG
gFTG3mWICalp7skBAE06Oh01WuWeRStyt1YEI8doNQMA09VKH5OqOg9T+URWjzg8P+SImPBjCX8Q
nwpi6WA871AxleGBehmgpOY+1xP5ouLIxArtVmDqo3LylFqPbDowKvMqZxSX/okp7SEqmBFSrlx2
eIzpuQNSvyfZLKtxZrR+2SW9Q1DKLHGvGcYi/+L5AnZnsn4i0HNtjLQoia4nTRiUcynoSYdvIPqU
B/jvulPVLVC8gwYhADETcUMy1szK2fBRS6TkB6QcRhGFjlbJyFM6mjkhUhGHgXAOvOgM1BdQonS8
U8Hjig5fMtTAj+B4wms0zoNZLdlVZuV+u78ka77+iTTcWEnc6K0uC8EkpyABZ70Kn1UOdevRzHGS
xBMg3bmMYJslO6rDnfDa6pFsNOO78nqNPaL9jh28GpfYNoNmw6+gTEwj7sX668sdF2GPavITsKCF
4NEW+0oudepe3om793Rr8HsuM2we6PlXrLuJoU4QSxxZCLhGlpoxjJnd39e4NZVm3H0QT0QdOUtY
r79WSUnn4CK7rGIVuMPljNlvpO7CHKCTLQo8KUp2eYqr3J1rEtaTCEttfNQ6Uky9pQgUq3S+e5f7
hKErTa3kuhICSNBL/+2tvigaCl3srLRFjLF41UEDr2TywsNpbBMVEkx3XlzT68TjcrPQfqGmvhYU
Iq6V3R6q3L886in9+xG8kbukc+I+0V/NIX1E887dZLWjMDFDdqlU0npNe2E54BKqyx3R196dYCpP
KpzK/Zxo2ApW5t96lcHxnXqYhA7M5T6NeBdPEvAEZ1KEehdtrgFyx/gsYNNXgj9dwfpU8ycZm9ym
XuRqDAwptxl9wnDYUP7eKK+DU0RjDb4+9Aer9XZGeoD6as+ELPhEv+vJeV3vUOkKu0vAFwvLmjEq
/AzQowFibTfkJvJsMF8+N4wKQxuXZ0sV2FdUF/XACvXuwAmNlX+beC5lKOBtfgsK/UTsmQ2E0kZS
QW45nevPEFEM4552kEdWbA9d5clLtCXvQsyoZncAZ+cQalUlRBnNkV5MBYKjciY+DnJp30W+wbiu
rsABnYMhMzZXm/bnoVKvLU1BpIUCC/OCBDMrRkYlq9rkHCgAs7HfldvLIMZNzXW8MiLGthjOavQF
JapuCHyB/35W/mp6TAU5byMKOLodsh2taOPyU9iHl1QVyVT5lijNnwrwD5tO6A4/NB1Qf4UEwqrO
MSJteAm9szgcO8BrJdHCcwdpdaGxeyelVttPOrienUC003kUqCsmdi9GdRXT0ztVNIBEJ1yARKvt
nzVSsxjdFcbe+xGNOGg5ftzX3EuhZjwr/Wuae0m6VnCZ7QBLr9EuhUXdRdFikWK1nBcLpqce1AO+
sI1CYTrwmMc4eipPSs9iFXOlBv/U6lMBB3qtQiZ1jxE3Sr9vqNMeqTaUNWxZDCtG8RqSJXyTKjep
YYOK2OaEX3B4vc/jKG+SU23s0RfCwFcPPH7pAnA4gGVsuwUS/dkeMcwP/heP3/U7yVNovMmSHBxd
vLt02FN8SLrAWaKhza/3eOQH//Qh30CvrxcrkEGVGxRAuCa/XseklCKj6Adf80KcGbKQv87gH0r0
7PYuRAYMqxFNwQeo5UqcJ80mDF4LBz0bA2Akts6hnyC44qJGzu0SykADGS5Tqtt2++SWrJ8BnsFM
/bNckgwWsr/aAYLggdMgV/R6cByp+sDr5sXebJcy1Wf3A35/JPzKYEWeYARuqJ7nk2C2hUK1xs2D
je/ll+v/fywKae/jYBoH82MzJwNGJhM3krXnKMO+k+OlU4X95ZhN+vJWLUGZaVdty5rXte8BRJCz
VV3cGTjEyK30Y6P5ClR+Ny07JMAYUIN13HvUYh4+b+RI41mJo2nvVztEfFBMQgr1fs2GC6FajpTq
QoJwltw7PICoNvK06q/txZ7aemCgUMNtnrwKwHaCkn1oROahcn0/J7133FGI2g7oiHFio3xcsjGo
b5+EjPI57uAcgENljoYyDolMApTsI6naYxnEisnIxShiU1KBUze57RyHZEv0CP7R6jq38RwZb5MJ
9z1Auuu3KAOQSXEY6DCfa0a15kl/8GpJGjrdvFjmw66bBUSaAx4n8QJ3Fef2Y+K93Sg2E/ooqWvJ
cbVKZ8VN5lAtQzOKyqvSZpnIQE0/Dr8q5uyJJHp35yt+sdzw5hEDvGOH1Fh4I/JS3ZrT/V3BJC/6
tGE4cuNfs3QJiw2LsVfNLDIj3RqpX3lnDrGqtKfyCWkrWAPUCr6yUsGkirx9upbnthShJa+tuXrI
CVGq7hLhvtq9vpl9zCpYnAvyTBFBaOk4V7U5rKLD0NTm79DHqjE66W3aBTrQDmZLOsrSOm1fNqy4
RW9WsU74LdNjH0LvW2074PN7G2jjUQSyKyKI3LYhGaGxa3uKxLoMLDiGwkmAxGeaU/vVGYgE+2OO
LFy5XnfFVolLL5T8FbWSayDCCeX7bng3vp2qJAyrC1G5LZxD+3gReXIOvG9HwZzRCeE/NUxIn5wZ
SYzLCNtfcfwRBCYEZPUpAriChE89RpbYqL3iLPN3wR19lVTusuLujfqPxIYXPxHateidhd+DvbB6
4T3MMBDczE5f2oZ2+MrzNarBhQXhuvwm49MWxov7Qmjo6F/V5eYw7Y+ilmJLwLqhz18Qa0MQ/2z4
5xtzXo6ZOvhmyu0mNB79ijsz8PT6zIjUXrXxHs/d9jlIBnselH1MeM4TYgEI+H8mOyzBKBBDU3sj
HI27ZpKspUhAkOZGFgGH/koDQmrXbiwyHLVo8nHgRhFcdMuAnhRqg/b3bLgtNqRq81PSQDM7U139
aCJ+9617EksnVF81ZgzAS7XUDm1bRv05JlbnW5b5cBA9KB3/Mtvxbs2txXXwNT5HRZ0f9ERyaNfd
f74Oi+fsa2Ruh0GCDg15pt63VYusN85uReYKHS4a4gg01uj2/dOyCo7nkDkn+QiCAYqzREOVMHr1
LyidB9fJmjclhImT6F2u4FA2HKWQijVzynkHFwmaLTiVjobjpj0ypCtAx7wMQzOPQmNBGaeD4hfu
3z0sArVqcg8N/XKXoAzcIEYclHl4hMX4bHamdQuZaTBTPitEyTaPZMjrm4RRKcljbmBKw9yAt/+Q
hkCyeNIC+jETbGGN5k4GHfocM9QFJ4j+g0jd3RNSJCAa606ladTtHMW/SCWRA/L+aCkYrRbFMR5a
q5Jg57eLIwR1r4gdISMVyS79kgcxO/xEk6RJz9ei1Ck0w6Vh+ZkLjU6Qjx3Cmrv/lBZ9Wzbp8Gbq
ssYQgv4UgKWeHGKr36YyuXa41SubVk+nVJ7CBA7kuw0cFfUpRuN/ET9ReziJUYoBKCLBQWCPCVWR
eH7Ei8I44P6clGjx/GOlVnphV5Xxx4VgnJXxU5k6AHPZRoWAx3aEpDHM5EG4wBBG0rK9bMPTD/Bx
f6hgz3qZs4LxJ4IyCMiQ2u1UrRB12MQclEoaRVL42PldqnjLqB9hhd/uCx6+Z3KTTJHXVV/UTorY
s8Vqzdal96d7qclJteO4Ht/R36kpbRq4D6ycr2zxgJbVLse6XAP05waUVxMB1IzmeXu1rIFcg72x
OIIqxKK13rydrp2NaqQi2Kj4a88I22FYKr/jGNlC0e4Qk2Gnd+zcMdjdsPhBcvDkpx62NxYdbnQp
Kv/MpILTjtaLa5tWAm8O3NZiqpOl53zq4/piAmeQN8B3EsbUzbhOHy/enCWAfzo5WvttcZU/QPa9
7lNqirmpn+E0MDuZ7N5A3vqmtjGrscpKPa9KvkUr/brkCGw07KGnFvLK++TySvKSm6ZLV6HrXUWM
QYHCkH0hvqGxhayAsbquIHC+XS0ymltU/RJF2pGfeDoDmIFmnxZOEyAeHpV48tmvQA5GhATAP+pP
k1f9Rfz1JkJovWothWWXLJAFBwcx5ZTBQYLqJblciG/gNTkHN+CJEhiwDFv4N6rznEJBbs8AM1f8
jygH6TlCtSnbkWpdFydZ9lD3LG14qakP2OiKsz3w3FENY2jEgQIjQI8hM3/gVBdJ9NLGC9eJcSoq
DLPUS79V+selJ7S/Dxo6lcH75/3wTj5l1KS8EzXUrShvBr+54d0eT7edeTADb6WIYjchwcljRdtE
3mw2/y9WLjTt3PVyc9y62nMMvhpidnO4ck+AZ/Da2QK55YcnH0dd2XTnWihpauFoG31L32/Ud1yu
+PmlrVthHWbdpoHComv70IFApddWMHnAFu5w6PYBAkGfk6iH2sf9EhjPZgolg1j0KXzArDRI2/IT
1AmCslgnpwOVxM6qpYQdtuS+RRsTFLv2Mre9qH0oLkGvaf27t9E/NNk7UPWTtrJ0L0OPUf2aJ7s1
FGbuO+V3LUq7D1Imt+xaOrUHf80x8EyOyiSvJLqLxftcFpjSdBMdvS0Fp8x+cn/0xgocIejjOwxM
AYqCnWf5jr28Fpn4xpbF+GrZIW2Xf6uLn5f9m6bV98tOKoaN/PF1f5Z/MXCya48dzERQA5EblRGR
tXrabVaMpdQAK4GXl7eSnmElimxKjnci+K2kxllaFaC/9F50WPG2/fvVwmMZO2u9T4Np/sOsxlKC
MGehHOIXq0SNu8C9nqYK8ty9vwloD0fLQIsB+mgc8UM2mWEBaotaGPK0GTJuPBw4mYIaLGE8RKXz
HZfvzgtirLUtmpZCeixK4cczHUT/OBJFLhYbYNttVTprcVMA7LGC7cAjuug1f+p/EG4RMtzb3r2I
UXnSM/e4PPOjt4KSCYivLzL1Pdx9zVFtbFSsxyJXEPtz0EFXGFlnUXwO88EymPE4REPNpSHqfesJ
GzshsgkTmB7ToyuDvyEjc5BTB1Im5xi5ug5CiBMu9hCKhig9WrUeZN1Tv562vpbjg1wOZ1yY/uRX
jaX/sTKaSfGbx8R2VJDGmd0dDEH36/OZaJb5dD6sZQHOI2b2af5D0qNG09qOb8zqFK5/KVmBynw5
+stQFDCDrr84ejRqIJTSPfSpSPfbRy2ey7o6+BjQdGWM05Gn6xMlrQlC+oyRI81SnNukpu0jLznf
zYnUKsA1hbUMYIABFKiXttfX8u6Hj2YVgHQi3OFxCmORaZe7LYggvI+NkTNQw3HEqP52Ho2mYn6C
2H0SlPD3R4UvO25wkSuSxO8n0d6tIKNjqqnZgyEX+ZwN2PyghKQkD9Ae9/NZkOt27ICDLrRcI0+7
t8+ApkLdDoOme5zxxQFXMctNEGqkafgYLfgrxWKO/NZxKue8n8VmNEKRarmlVTrhuk9UHKdJRQSO
nH9ynX4jjQXsYmyKLkw4JHnP2L1x7aC7R0hPyaV8f9AiA5gGpp024TbY2G4ynBICQz5qoK2fTTAp
FGsLyigWD6f0yHLoPORZY64s7zWhJ2Qul7P40UeaPJ654c7srhcjyIHNbg3wBNs9qfjrqBXyRdhc
hYXIfnS5uoJvpCQMxikmg7LqlE8AW8YVn1Ub78W7LPu2Oc3BwTaA+rTTKFu8ncHjT1Hj4Mxz/vfq
0XNkwCbSDoAsTwqW0UfCsqUCpDFx/swQ/Ze2wOkVNjTaKNyc2HnS3sXmXJKrRL+KNTfwm0HoCLon
b5fQpZANzUwjef7XDBW0RIiiiIpYPn/8/wHNr9BSHTDKbzq4qot5d5WtP+WbUD2fvnYHiJFTfPxG
ONyPF5C9sJJDCZxs4dlfBmZfRJNBS7rUW5nVP6QqFSuUhnA3gK/qn6ffL+ExV0W+qKQ/7As4HYSQ
EF20wRREEhHBOaT4DqrnS+pJZa6Lmwj9VHPNvGi0sU90SUhjaArPmvhc6FdA5P7Db1fhqITIbN96
WbQryxdP/iftTpp++6yS5xxLZ1Q/Lu0D6jmxLDk9QOGSveR9reDvJ5CT2tIqwGOfAczQoVyobyA/
grISZMozVZ88RIh2QYUmPQMTc3mOybYY6g2X6BojRtbhhwlDmaY52yQMFR9DnS6PWohxtWnl2t9Y
Fm0XFB75p11MxwyvcJrj+awg0Zr1X6rglHzRRS3I5zfq4BC6z8lSoJ+tcRwQu6jDKj2UZD7n9tkz
N+ZMHEhZB02Q6mXTROKNvELWq9xgml5lfHVCWs8NC0kPq+GZbDi5CqLFksaYWHt2EHZ2vEZdnFs0
M9KksdQPpWwtWeSgyoOe2Agkp3u/zwzhQ/B/LP85PuHRR/y4iDfa1kFUFlkd+EAAmQqsaXElDsNx
SQQI2e98LjEOHofYllM5laMWFvQyxOqVu3thG8hfmujw512kLSTJtCLY4GZrmc8CP1cQ3T6y13co
EvdbLXJD+gIUedSP4aI7N8Luxe1FHg6rzw5wbIFNFYMOHJowkIiQoLfeX8IcyRNzLh90hSBiKBkj
BPKfeFky8cYkc/JWo6MVk7TQ211n57z9YHWDXItGuXrCH9r8oioIqq26guxwSazVG/3ftTaV0vFG
cXxnb86X7gjjtTGFepR8wbkit53iKBvlKHCs1OOZNB8+TrxX1cP+YRlzv2cJbWh04Ua+aNsiZl49
vZnPEPRqt3fj6T3yUkyLeLVTz9Z129sg9uLUe3qVoylrvzno+wZcgkd4aY5WSWQu7+R2zBkdUGSh
pSkKWF975B8zdMPNIuf//zsU2a3hra4zp5jjlTY+AG1hnY+mlIHrtOJQIg1tvwqI8+1eZbMEuiVc
6WIGZPN9n+UP0ieyvNUTFDa4LCu38vTXSU/e0wbUtsgAdfc7bd3JL3RbCUnu4pl8FUhperszbtOj
GW3jgNrrAhiq4a687qoHLD5NMVyzTcHysDJW5sCzjIO+qpJh8/WX1QwBm0F1d9nqakU7jzO9f18G
JfKddKmojzZobuZhcExTamZIK/FLaIQCTOLf/l+aSxgxAFxQOSdhM02Oof3W5vo5FbWIgdZVnTaU
UVfT5hqGbdwF/uEA216tTZWI1W5L+Rn8P885Fno9ta3O69d9ro5rnCBwAoQIrWzsHgX+pgVUisY+
QNoVQtvzkO5+ezFjw4g48jKpn7ub8vBXrE511NpxHMwGtz+ryg1PcPCsZgh3XKVVA7pEgiNQAGWC
mFo5u5+e+B5LOz3lV7R9Q0j8i/23Ia0P0kGqDTAERSMA/jn6iumnfNVBEDzKTH8GPR9IzPesH4Jj
EwBLDS39Kihy740c6c/T7g3E+gJZpuImjBdnRkJvOp4MM2EKiDpR+II60VvyXW+R53uZY4btQaS5
OWndeKFOwhJDFX0MQJsEOTHWSBJsvBhFuxPC20o1ETqhMpxv8baj8iQX/eAVqdPdLKS1FN978RhA
6BWAbGr0NAsHIgOLaBAugJHRJHWBFpV+zDyKjh8nfkRqI06phBWWnNYuQvo2Q9U8Ax7b+Xo5/xQR
nXweUfi8iMouSoWnR42vlGC9mEW395IfJN/VMaFQbmUh6Il8jdNydxhXdSXluLoXxjh44HxIXF+5
ACYJJliibpIAZox4FIFkifrQeq/sOYj8NeI3PkRH2v3ziGgUguNQ5m1gK0pGWaTqLI9P8UQfcKBR
XBbyaM2G3FSCtRtAeVHGhTGpaNhMAwWoNagtUmNu0cLfYJOPIpjlZeTRQy59iZ8Q7UBJEvrFlU1e
3BUXS22eeT7nlzQlRuEPLF2KeoBu0eQXS/i3jNsZMZdgjtsY3GuotP2atKI72VkTtGcBFxdIc97O
/Z4rSyamKZc9W98ZI1ZJ0N231+yTyNquvj7Ejx8r+0XL3CcvRT1Ya+RtyALq/8oycs0BoZmgiAQ4
DpZUZ/iz8KDUWaci8Va9rjEfUQXLw4lHf/ygETbUEkFH0l1+nXIM3DdEah3LvlZnNTb9a8iMn0HN
8+1GHSjjOgRj2PSK5C70REzY0skUpN5sRZd/EP4b1GvRvQBM/4/78pxzUb17xrNEIDz0jT4fi/hy
DdepPuRq6avo3LyxhQLpeHIxQ8mIWw5h+6jzdja/xH50QTtCnZUxA4G1wvZnGMLAd+Q2p/m3kiBc
krii6FqdtFHck2ktjjbiBcmEg4q9v1vqcRwTfj+Ak+B188XPHZ7D7ugouNAHJHas8Jr8BnjcnWGg
uBKItmjJtywjV1O7ynlkl8dyAaYc5YIt/8Jzd7aMPbEyjeg0RoTWAYu8nNbzUnBFy55yl9moSRUe
WwX8rK3gWengf1WWIlOoCXUVSxUOCRYPogpyW6ASESkXVvM14l1fpfy3PydsS1iWZBbZHYtM4a1F
DNNYgoCjra2sBpo8i0Dz6d60EK9VukdZyLdNDqJno6bytCN5pFYaEmkEdDbm7FoclJinC1ZAZ2lz
JvyC+hstjFas8KJW8QNYYz+HStWHOM+JtWl+3YDCxqSCbh6h+kCiDbenNmF1pY4LAnYpFzVU7GHO
0+0vw6hVw2+W7fdXypw7QAQ53jWsiwL0hA7toQDx5S/zp0tAEb40x3yPrCzFfI29ziI0XOKVPRh8
yS/wwVM/RI04Lll2x7A7dMSABF8yqq0fbj3pn7IOGreA8ow/ijiX3KYVoRFdzpi0BJrjiVVZE5SE
SHR2QhoYam8lNNO+Z5mlAJSmQa1Ksz7xoIicGHEnK97Y1MkVT8+XNR2UBUw6GVfSp8DzVXubin5l
GVwPQZUFWp62asiJK5xHjWJyQbbgvjodFrS39EjtHdvCwlvz11fVVD0RlrO4BepLOLmvWEuoLPTP
yosJXrq1yBkqBXKesdgiK6v+LDJPn5CYZM2PQfksevaxjbJEvoDNxtJ0zqp48qD/fTxw+cILS0c+
HbfgguH7sVTaQVId7S1iyfFIZbhUcJ5eWLqzDcXEa1j1uutXni47IJuPnYM64h+RDAkDH21qzW+R
HpmIQ8AvTOHmQnvxSeYvhL8qdq30lajAW8LC1RMPERc4RJv+o1annGkA19UFXxRJr+CwlnrJVANy
Z3LdtDHIfQK/+HKsuNtEzvfQkqmoLSl6iN6lt0WCByYfAw+rBj68+DWFakY+8/fQv1ewlo7BQUvn
KOwkH1vZTrr3beGsUN9f7xFclG8bXQT00I9DrKWLTBLa7lIt9JGLWot4SX0bIJt4s2W8rpa5ZTsx
2U4i8+rrVoB6FuPKNHnjtUL2RPsaYs1LyHi0239lxOOcG2V3tQzXa3l75MNNzn+E3ZTPiVIseSXx
uC0ndMptQl1DkpzSyL6jPSszSGxo9luPgjvDxTQHDgp48e+duWafXcs/E+Oh50ouJBv2QgzJFa+e
TgA0ZrMrsz3CrwEDtoKeRfi9PG0Z7CdUzGXjsehgIxWLT/DhjUs/cM59Far1S0oKhQ/pErINm7QF
chp5EPTyTNvgCRRjmMPUkted/QoymvYQOl+zuOzE2VFLBvxAyotdeNTzmbIzondyb1IcqWrnWZ2F
BE4OsyJSR2xLwN7MtvVCnUeJBDX5dGp/PYk1F7H6kl8RAT5QoapRcJuQdVnY3ezQOpsyr+hTqlSF
G5d+yGueNnCQJhSjNTk9zKvE7+NUXt+gVvyxWjCzcelDJ9Ah07mU2boiDTuYZsXWrFBqyXaY8GGZ
ag/TMGF/Cvl3olcrZnwsi8xtlHJfSp3beSWAVSoTQvN8cHT467659aefImNuBODpMIJMxJ4GM1D6
Y1W2E+++CWFBwZJtFWH1Lg6tH6nItpsCpdoZlIpTea3j/KPEz1KmapP9cYkyhCZH+3u9SygzNqXH
HfE+xAy3/gEtiixdwTeASXuz1VtbATItTS/wPslOB/muuYqOJWxLa9cbxXkX9NrEzA2lCEj/lYHc
cVSU8yH7tTmudvSKPdi/CCmW8xc71g5d1CNKvNRPux7XM2UOcICioSSyOZ3aUmOxz0/xYPvoNGzG
wtMTPVIj/DtV0LPAHHYRe2YcJ7qPInouN14LPYuMyGmEG58MFWNl0/CfnGGMDgXQxu7VHZf2N/c/
QCHf84VgPyKYi478a8Rs49pE5QtRqFhDWV9AZLnnzS/6eabqaANBBV2MLhdTotsvR1FBgaCpQFyY
dbtcwKm+xockGc80lGgoLaAX3zDld2tOxDW5zJ9KA1+/FHPKXnpS6rrQeF6tMkxw5PN6PS/NBPPo
ei29nudt8HXKvPBqdho0OupkI0UsoVR16YEbva/juw3PVnv8+chElfUnrwRn0GPA6I8Ni6UpHnUt
t2VpoJVdQ2Ldkri/ywSWtsPsqDjxc/aMibGuLjI2wTtqXMadavOQqJm0lnm2ybNzuwzVZD+H93RP
DfYP0KMvQPOnwNYqREtDWOB6zwWv/MAmW2Z5+iPW1UmEdpIQTyCqwXvODcrpklRnpUBwV1seZkqm
jFQjgp7oublkNq1XHUYkFsjBq53XiqqzB+yViM2uYbMVCn/33kypFj4oV7hPWjz96jOTUdf26xnf
l5kGs61EZk6yVNbnBjM8rbfMj/2Pln6xTr5F4o+lNaXfghFtLqEYAYM9sryPZjoOKZe1LDepHu1C
M9KnRb/MHUuitEmr6suZY4eA8k8iZ1L/OqM0+fUGWW7GQhFcW5H8tjcsbPXob7pzFdTb3+YaS9Ri
kbCyhRDqV72l5CN0BDKlCRpiK2jJvF7q1d1rW4yjNsyGMitPyBqE30Q0jkfkbUYjWi6mQXQ8nraK
ndZ2le+jJoVqPMB4HO1CafhWFvpJyr5SmCOx6EcAUuK1Ti23iTYdK9XCN03frNF1dQpRnaRqAwNj
4ipqnwSZIJiWOUzrSw8KXgrZYYdk2+XnJS6o9xk+LUMA71JIkOScDG8pNGrgqbIZyXPWUuxGBhwa
DQhw6KoRHgeHKw9WBtASFV8NwYNDDVNIdjnuEbpcEHGnqn/ZDNcfxCnr+jNnWKodc9aAii7GQjS2
R++OyglxRN8i0EAVS/YVZvJNxIUind74KbfZcnPP5bHw+2XLQEKOqarUzyP79bOSlqIcH9kOWZ+C
gma6K5FEI8/XeS1NFJFpnExVyDHDtjcAmbq+aDbAwRfdkT17T6qQ2kqulkKVdLVYubMmz1g0uUXs
i9MoQ23BkWO+QSPF38bArV8a5LhT/PF7vC/tZbjOQOpkazahlz/eZCo8h87ip9/UFIqlEhfaV2v+
IOQ/HAtu2XNrq+haispBUkVlTCNyzY5h9fBQRC8ozr4yeZfVoh6Kj5AtjUHW/FoYjd7gh3uRXEcR
gSzU1TBA14vqYSQYz+Irisl0hkPNufHnidhnlk7LVipl9r06FLOmYo9N8KL7kDiWGY51MkBKA3np
Xx+Xh01sS5HJCtIX8+IOwpI3obsktvf+Bee4vyNL8Xqa+frITjR8ptOk/AMG9V/1DCBWsxPmvoRE
4oni5JFY/3XyUd3JwUfvNapQgl0Rnra7NMgKtGviZHEFg3sf24NExE4cNKqd0/F0MEZPe/+8hAJJ
SXlvw/hwYiPjAhhnvvIG/wKsR73Q1KdOzoNLpTkbAlqssqU/rLLkyLSCovse5ZhDzWWsHk6A8AOO
qt7cLlvsANTlO/Oo1MvRTymwW1jE6y1y5L6DgB49E3ExIroxp5WWdHyf4dWq8h8kgHiMkaH60+DP
ZQllBqXApcK1tvHQgKBvEv925eCgsKaVUFS6bfkINjcD2DmYF9h0bqLuRjuOGcBtJ+Pr91i2Py39
GM/V8aO6klf0iIbxzuch+4P32aSG329odSoH23BgTX0/PhpWuFYsBUH0cXZkY/UZwAzjB2pZKTpL
CnXpGzRhS63yrMz5j9DzAUnZnzUOttXgPhaoixz8KnC6P6JzC0hJQPKehyy0hLm8k9JjwUaltC+7
h+Jlbv5G9CAvUIteo9C89ko+EdvVO+LaBgIls8NIA17Ubk7V0O5Cp23e8hi1MJWGqotQG+iykkzi
aqGtBcIkN/fRCfaYC7cNRhqx8mSqkozw4PuMBX0xSw14IBEmQnbl2kbRudS7r3LL7k38dOZ5cd/O
EuD+bmdLOln9WhHN8pHIRZisl6vzBPdsgS+o/9sSYG2U3/nLb3SXRYFUN8zIqW5wO4BKFpwNMQV+
cUjvW7t2VtnQuxkSuZFpfUlNEnKu2muKOvfRr/0J27/mG4/ezViS4hFAeFEEBgJz+ASGD208/yKV
GsEpqjKIYHdVdSngYRX65EBZ86gV7f4h+DqIfWpTOmaeE0y0HAt5wF6yifT808knUasIzDTU0Tsf
SA8vMJiPcfzAk+UTl73AnC68QFpG9WK/f2tMs3gkKka2zXpVxWJx7uGOdWW7hQ7Rc0pcJeAX6kKW
jOGN5pi8rk2Q543LU2xKhCOVqXlgcoXwKvsjN8T/PFN0Xnp2fFN8tt+2sSiL53pbVPXOgDr+OIhv
zaET67LcOqbKJL9u0e2praRaO8Ldpp84nr2uQKNzp6gpAAynh6PqwaNgpDsWgbJM4s25i9/H5xLD
m5FsHwiAM9USPtazF0sGBR84GWrHQlxLiPXFI7mupOBAuSXlBPca/XP3lhSwKhqKXnBQ6eeljews
sUmrpaFT3VVve4YtOMnF2g4FySwXwa1BxTMxkDkTuEFCzafpTHlc1yhqCH1bvW4qumOR7lpl5d21
2gX9H9RwIT7JqJ3XnUfTOnnD6GQApJMU+W/CZiVd+uVAP4kTwyG7Ob80kw7wMFPH2h1Ry4XHm13M
dgjjv1CbMAZeYMvhYOnzr9QIBt4/IhsM9Xsm/CpgjNOT10HhIFf2KDlLrgLx5/b0x2h631KC1o/3
YYQw/d4yeWhYB9FG02rc8tux+nYW+qQiiMgEmohZ1R37ZICHYt+4mK99qiFGTSrap7YTO7MsMVMe
fnrv0ZAbP3ElEeSNoTYpJVqT23gF4zjqO64gfNIA7HMlAtyHHKRLr/UgdovVgCfzeAk9mr4vQCXS
8QyoAzPyotAnPuOJcWVfYx9DMcdPLRRHyv5O3fGVlhnyszGHrVu1HdE0d3xjfNtOG9yy7NsRHhL4
PFUGNjdjFSjxizpGOrYDGKUw/Ljk2qi1v0vCSxTUL2vQpzno3gnrsWmYr1yozcy+T4LXgl49DwXH
1prz8FFwANZa9c32Nu31DfX7uxSflGqHmumdfgxA8+jAyV49HWSqyGBTelv/ZEesr5oxFM5Xv7ua
HtPDhewZsjWnjsCoA6QuqW6K+Q4Nt2mc6c3AIrmxTsRjLI2zphaQRyZ4EGGqsK97uzncuXLDG+LJ
6YI8qEa4RjmGADE5OiNNIdyC5lUKLbtj1MbCJezND+qDf1qNJ1RV5SjYAMN20OdcZbgbLjB20Via
QTa8Ng8khmURjYjHYIA3JPucxaBXtlEuV9FCtqtCTtyvQi3xGWme5OGngUGGDE7HP84CGRmwOJJ9
unyzKUyOVo7jH7PE9phLi3HEN/NfdiUFv4/VbOPib7X32vvYOPMtbXd2p83ze16ByUNQLExrcpGj
JtO69ZjVKuj4SA+uOdH5VUu2z9lNib63p21ym9uUVkLmOKjy/wTNuZVhmRpxlENUsmZKSbZlNIUY
o/sWBkkgud/Bj8D9ocayxjif1jcpSmIe7Ken1tUhKWyPkbnRniFugsx7A8ScXmK3QJjn5CKbrD9n
II3hlMPjjoEdKlbddu01N4bdrXKmoTn4yLUynKbkwILYpMlVlYr3wV3ZhTEDgfk9oZeKZruEi6Gy
7htxn2B5m20dUhs/wnxYx2h1MZZzlHQbnVD+jQZ749rIhhO4VJGyASHglb9jpv7JqMosFoCqb2Zk
QUXUd/+x24/M9C5LkeeRhygCvpAyEnuURzfJLM9dqOWabTSC+ICoVX805Xnn/r9Mxpaf04ssCfn1
xIO9sAUdSOay2+ubtabzS0wyeXitZvFRXJsFc2IR5DmyH0erpOOp3AXxUtaKbu5sO/20X7GR79zE
UPAEY2GK9n9t4D1hC70Ey0IhOKTKI7OqrxJc2l+Z8GStmUDkp8VuB2U51jM9juf0sGKqXT+kAXoJ
BGx+5Xd+SOHsrDBb1wt6STngSFrxA4kQd57a3cuZ3embgy4ugP4DRUlvL76Sjzho2TQQ+gjUHsNs
D4xz2ef/eLG3yHXsanCx7Dz5kE5AtXTFqE6CqSfC5l8GGTzdJWBX0P+LQYzHOCmCi6a6toOTmtuH
jOvWbQvtU060LBQOAReKn+rkPOeW8z0TYTZ5nRjFhDZGR/raBtQWWvQFHyfx+5vaxAgJZ14pd6GT
ODVLqCnv42lwtr5sH7VTjE4k+JnrYoFq26OLw/PPu8RpbITve7sAMqNfNsb/DhYOmkNBncgm6yj0
S7mxGPZP6RwGGKJjRgEOWdWwcgPLVemZ3CXPkXcKzZkzlZCCqR2w0tSmcSB2DawZl9CZBr3Co1sg
g+Ed4QoTZ5m2QzflZtdrTB323OBqur4byp102og9w0xxJKE+mIgwen2Ed+DoJoqg8BkQ0nGQhIVC
CUIwYZ8/eM00xedTv6yGmd4s1W6eiizvSnC6AE/bkpNIy3F/z2EZqsB39L/Fhl6Z/4UpZXFFYHM1
3bjk6thr+xIaFvYacR39x6Rla1X17/JMGEjk5lTNimR3JPmx9f8tmX8nv5MnqlYcRn4D6tQrwuaR
Xjh0QgzKmkKWM38XxeyXzhwBvRMM4uUUTRaZilXhpRQNjWvy6zjwgHZGhA/MuK8r2q1yXDjEO/N7
1Leb5xo9JGUOlSHGUPbPZgztfICB/6rSnkwd0snPT27q7TwKDaL5PuvOnZRJo/3t7qrL1Irvk6cX
gPt+HsR7GZ4Sey+MldLYfzcJhs7BYICKF3749JfDepxX/bGZbmiXNTJErVYS4C5AZVcNTQjvrCUE
Pgmx2Ly0cPLk5a43vDltgiEZ/PYGaxOXUABj18k3cwFGEHyhOaHKSebrmt488EZif/0kkba78Vt1
xBCJTqMom92Zt5a7o2mcHuv+1QgQPx7eeb75FKmb2XHy9KlDVbQ8aQsruYKcFpDNMglGSRhsYN5A
ph+EqAoiwr8qChk6/YXDOVrIwMLk6gftTJIthIW3q+mCrSv9enc48cKg6BGbpLEoXEzAkdu4wZ/A
yDii81/+HppIWWB87NPtoNYbmme2OH6F23CM+78K2fLgo7ePivcbtWCu59CXVd8o591zLaiuzGYb
YLtQAS2rmbAuL6h/m0zSF+U8YXuqytzp1qkDLkZWVin5h0MtIAd5W1QrhimlYS9q/1LiPLUZ06Oz
gyKkoYSPuj+QMDayBfjDZ5GpXBvMB/DV3Bqh78cUQmtBvDy6g/5agTS+oozTf048+lylVVPd3Q0j
ff2ufhAMgQbgSiwDlmkw39ItaYHMhXUh94G6vuF7l6M5bWnJl2EuHJwhTgIbHA1D6TbXGxP4/0EK
mH0BrEjG/QpV5xbnmmgCEHNRJChuXGanIXdkgSxGXQfO5P6abor/4lgsBC84jKoEYEKNxGF+dAns
jodruEftgIS9xUR2V4CxJQoNdsQJ1G2ICAtAA+pzvd9f0JsSqXXdYLtp8GeFRSVtQInso6RszmO1
Rhj4OPQcFVoVUrR+JSGZlZ6bsM8PcN9Yt5tJAC/HOgDROavNbMRajUV2nX6YsjPJhMd/EAaAswx2
v7/cigfSzYpg6gvwyZNpxcPsir1LQ/5X67qDmAVLpttNfOQvh1vpaXDU2euUyv3A9tcjScbDnHLq
kYsp548qYVaDw3vHhJ359JXJvUwPpwBIoZqDhUbs1jo3d4xqyX2mWs4fAiCLFhP+/RbEgHeWBArH
hVZ9tseJU+JUqedLuz5fH28/6XKEDo68jL2dNGAsGTPuej21QX/zbRPmRk2g599SVR5m+ifbQcXu
kzparERVVzP1MEpgfYPSNSi9JT2Fl5AzP3ZUS2G+XdjMKbuxJSfMX/+/ljWqjUwBgq/d2t+GHP25
U/GrgpEKtvtdiCk1+yE4VjdNLpjy4jgfXFlKP27Ek3cCQm/0ohz1zn1dIEwkQzs5OG1gq2Gr4Y6G
4A3YYpMstWM5u9xdnvXaqgt5a70rHx8feVvDdMFLlvkjyt4+UGaRfn4ixLiMO5SKssd6fMhiC1C3
z9v0QCNMF+AQl9YOo2tBXcidFjqt9PbkutSeU9Okv0Dg+aPitUmS0dBYaJWiFx7djNdgh3k+/pzC
V/SmQZYup1XUyDKybpLUPM7UG9suVHCAuztV2V15zBHhnseV9oh1VRbr9womOqQSIxBZlJex/2tR
wDxiRJZ4T2b79O5dh9eP9XDMAeiCKjybIvM2W7kbvTlG/HhSAiYZHPF8lsuRYnGoHzvQUC9qpyj7
OzSM6NWjiYcZUIJt55TL4rJird9zgkk1ZmFjjo/GjHZlPzhMUCi7N6BEIbAOtndRoK7/1t+Z3xz/
8n8ohhO36h+f0Kp4maNZR2+OOpddrs/hFzaFgCOHL3ajr+ke+Y8N16tJkTYWEEj5ehceWWATMkrL
Y3+gHJBTug53iMql8dPSGO2aE3VjQcscoUWo2R43hcprSh7eOYwmxNLMetBogko/AgjJBQZZrfI1
QVPfc7F3NaHW7p0YFN9xFcuhjMLsjBjFAORX9zyw57P16wVpYJGN8VIDiQK9Pbf0UsrbtcfBInsU
BmMfru6Sprg2gNyZmz4gnYdMqt8tQ8D7PH8h3xziJ7viDU6nRlRhNFvKIo7bueNAceLyv3dtTaOk
W5DWmid4u4ZgLu0gMAUjNIExHV2e4NWdei6ZhEk6OrsILauEB/d8zWDWBIRWYFmtWku3vRi4OoMF
MYyyJG7ZpPXWbCuH4HALo+4eafa9pfot7AS+PMqfm3cHeIS4liyP7OnTrbhNddt2xfjv0/g4FsBQ
AWMz1D37m9tK8domFPW+uMzia6Dk4zG0lydATkQgZU5mlRF13aF3oj5vKR92vHBrsqL328ga4p0p
HaspBxhtM3BFNmxH7L7nhIQMioxV2UH2q2XHftkvpeCaUykxZi/iFBaD+7Oz+WhAl4ULXlyxeMup
qFQ52spaJIgDbFro0LiYL9mY5SmRNvRxO11UGXwWXc6fY5cenT0HsANvR26jeiZElNIiNXf3l2yH
0fxeqjowCPpibMi3WyLvjZEULWA9XQhttdR++TPJ6KDvOgC5doROMlGRKz5/UFRFe4f/Q18jt5mH
XYPgd4V0XdDm95LAvJQUUoYWGk+9mu/3OENOTRpwyvtfohDIp73dgMZ/wMp5yV6ZmSp595ls8iIi
bj9ZvjOwxT2IBT3dx/b8G9uwxsRMLgMjEndBjFHaLv20WbYdvk8yJb/H/0LgksqZLaD75skl2rx4
lO5+3dJBpUp7vKifBiPM8y6McEPMZTc4jsxHkVF2DLvtvTSulTgN+sGOuuTxCM6847qIs862Br/v
1XwS1YU8wwmhjv0iwelgbduz3QpGjNXeMsykF3YiJce6ZuvrQymGpyiVLICnYqiQxrnVInCXod6l
vSE2F12GdRKJmWA1Z8JGP5TafCvBUwaLpoYbLuuTrLjiI/YWJlUEMMHFDYK2lktCgYLzofkWn6QH
7L485t1BLuROwq5jfXX+mj/f35z3sxoUtABZzGU7qw4j/jRuKDo27h5pn8+snSF0plBCL6Nj38ff
A2HyA9UNPflZGLZqioPCBSXzK9NJQ9ogaXMlU05lNr62+JFUwts0V97W9ffPiDiIj9/p7S6Y4NQD
AhJbbY2jaErn6gNfbhxAXPtIW1fNV5tU4lGu9BYNnLjFJkPEoEYRByrQ3dW8zDNYIiagcfSlrvpg
ycy1Rb/eP/Dx7+4ZPkDiLTyiMeZ0et1SuLrqU6W8EogjkVM7xmJVapBl8fVhFNYLhcx6RPFujuHW
ILiypfGC0b5bw8AHB9ZIvVvvi8foayorbiTZtaj2bHJpNIjv+dc4848Q64TwYbyzkeSHLOv7Edca
/ez8ct459TtUhlvnyqenckkHnhYynNKJ8BKg+MsKAPU//29dpQCFcx0vkX9Vs8jK5cVizYgt9+ru
N7FOtMzHD4aiNFiVqWcn+6VIEuT2Qr15mtZh7Fllu/DWFwa8m4DlFovGQ275WGVg9HLDWEIxNXrM
F3qBiTtmUWOwZv5+HJQRAnKbfZpedIiStC0gJ8L6rEkQMPEx+ce+bWV/hxVzS+J5dbYMw+r9IKGP
Eo17VsRpchBU8pAJg0AdFVedEQac4k0lERI+nqkLHd5aSFF0JbPfxJgH5UnRXYapravEoxIQ/06T
L8MpgvHElRrrK3EABqQ5xQD7RtF+pYKcEL2bUIkadjef0ZyRczBjmwhEfmhEQmmop8k/p01M+tRq
Dpxk8JgxhsyCqNt7s57ZkvIbHoHA4TLyWGOe43jPRnpgQHyGp85OcSRQEvlvrl2eXnLjaEJhf90T
264JwxF50uHP002CzIutje2vHYH89qT1t85Rl8yI2PkGC/Zdb3wZ3DDM8C1mIrSfV6kfWBq6orQK
IKSJ9+3TqZgcZGF/hj2apAQOfNaHD8YXShvwVehcxCYNFf2tsnaMfjMggCuB6pYHBpH3+XTxt5uy
krTp+Qx1BY9aAk6lx9j/ck2vpN6lDhsmPIgJetvzs3dNE9shsT/fX77xrzQfj3dgrlCfHVQUGWuM
xzOD9kh5Wfy9olIp8J/1/DUj0lBatP9xHhKbpW/ABMAlLn6WplGpFhCs/HzPpqQdiov2TuItNEWp
Vo3BfRyzFuMWMeuIA/FDcXHPYD+SpP3xeUAcdwMwbHPPGoLZvKSZCFaosKqgu8GEXQCmUGNsoVBb
kcQB1gfSiQFqxziCeUl7w+H+pMNNaSq4Jayt5VVNirE2d/kwPWZhRGiJhy8iaRHiyVl/87tPFujX
fTznUPUrSVhxP6XNqxjZLTHLcXSzluDYgzQKnIF01tIPNMzHCYXpD0H+7GoElh3Bdmu0uug2bl/x
mxCHN7u2L5XtdhsCcGYq5iqvUL3nwzRT2aBPOpuCe1JD2LCSnSAq+LVGTw8MKsfeJG/3uj5jtwZO
FhANgJSAHaXYyaZ9GlzNx/pqQ+8z8ydyPaasKb+kZhbjq6PALjQ1+ujjsQCaFpCFue1cpIe3mSuj
+lS+WUfuEu05Ml/UCkIyAyDiHhwjOOu/2i7cDKvWmZKtTD0sUvGqHGtnLzT0oyHGLjo1o2skED8u
Eq7Xe9/x0ymDmt7F25kkzvoEl/Um6CkHKxTKqI9aHS4e/EEeS2GOwIo5fy/tRlkQ2U2muUu6tMbQ
EOLpqHhUQH9cduG8tO0noVMv0sDQ30ayNNCSw9K1L7PXeIDubNxElx6NceGjrEWcwPT3g6KACoeJ
juoQgpyX+Y6dG+RoxWM0sNWIgOVLcV+5mzKUq5N3cNAaFtexEc5W9qnVmRmxPWpt8wg7I0dXa+bJ
mHZuR5iyvZ2m0ZIzBEIgYAZeNacmoIHhET6i/zyqXWN0RoD9S99Xr8Rqv2UxFYQLKTjG/nwFRFAu
Bxl9mL/ldgTL1FmPjblXd7nPamhG4B2KveiRaQDZpAKvw5cCCsiJhrIvcpGur3pHdWNfFTGIK+IB
mbBEt4230aJ8a4QSCTn3m1NOy6JkoQfLMuNZZVICNfspHjglI2d9l5X1qRd5bvysExEiycofdoXd
YXhGN7RYKXBpp4455MwO3uWPe264BaNo1y93In7rCqSS8UdIpii7ma/5XYZTlZh9vPZlIB3SukK8
yP8EWPx3r3waTuF7e96gN9ybwIE9WFDUOLgarZ9RAit4gvEXVUuT3/b/Zps4KL+TZdnRAuu4iIsd
LKL3hAG1heui6o0LqLkzLONoUJWoFywLoQ9DcmWv8okK80RU82WqcC7F94UUR9M5utbqhMdaZrYB
p9zHnaCAZwQgE6vCnhK29wAW+Jg81ouesiSr8KJ3jXDHID++UBGXLYAEzbMzlA81i685Ou21a77G
toIEuamV8c6R7qbHKQ7Yqs2d3Dgzv/QXUQEpHc66UcaNINz0LQFsk7+RxZGLUDLh9taCU9it3Z6O
xOdZ1Bzvpiw/neVxMSinYYX4xCLujxvn10DCfIlgIZrbBJsQn8V+SCrp/lIdXAzHdGcPm/z+J4sl
ZFNxThGjzLTTfFIq69XfeL+FMzk7QOZXKXURD8EWXyxHuYqEzZLmIWycDAjTgC5KIAHpgmODM3ZB
ORI3lNr9VGmAWO9q+0jXflmvJBhB/S2RbjuC2eXlrukzt0Ia3oj5gQWaa+gO6QzyAMvunp5LHBCy
ws1pXa1ZCewZdubLv9odhtdb+7rIWzQ2cMX1CM+RAcoPEdZ4Fre0fWsOVztG7fKLJc5wTumFX7XI
CE7aac7SyDIrKJqte+3RvFlJg2OsEY+HmQLJnxpoHx4pZtLECC7BchiWVC+Y/vTw4ECh/4PIX0Gc
gCk+3d2fAsOD/rSVqkMLSQ7VofSev8GFJSuza/NhqmVgZGfRxgHLDl1hzLWcy/KEP4dTURdGrIio
9vwX8oJe8WTQN2cIc2CvecedIP4n58aDEbSNJniyKD8VGyFr5l5oRuTqGxH+eAUyfViYjh7yfarI
LNE6fcdXwoNqNma5Ht8IruONYVOba9sKJS6zCIYcPmYCP4wHQJK6AGEiopnRVlNR0UPvIxolHDGh
qmMVsMCWksd9CpwsutYW8WF8KR5V6N4bUYKuTHlw2ZKyjVqmyJxv6ZYr4iBeuJlJh91itvq7rIsK
Nl1h25gZY65MESgpL/sKc/Xwu5JIwHv/q7VCMg1/FDBNgjM9yddcRtuOGEfrusGV9hA1Y7HD4uB2
FD2Ocf2hmWisKBFLfrg1sFx2pGLwXCaGHmjeWScYeBq9u9FaVTdcNchyJzuAciVobxt3J/bDKL5r
GduudZI6rp30rC8Vb07IWno1Wtms4ITuvuIySivUQxADt09wWrAyxbwp8TAuWI6WYDDCRlC1f1f3
fLmPqUYjLocrYXgA19oFIPcKbPzt6LttqmMmbG9XPJRNtdTpVofMtnMBHOP3aG2WvMLoYxX/cCcG
FdL4WnqExjXu57GYqFknjtarbyqH7Hp5mjTbDsq/gYyKzhUixFfCk9769D8PRbPwt5j/JIRn7JEB
3kwiugyU5xHkiABmDfHsE2A1MyKH2wjVb9NpsIr15pt2eaQHcMVhX1ilSq08IFmGZIKEJvbywVVu
bNU93vbvO6BDNWZ8kIDvNpD/uNjlbzX09NfMg0R8xkpWPoSw/TBdBjtZPiUh0FkYDzyWdP4QIlFm
YAdBZon3fLjwcmB2lLV434HgU2SDIkktuRYKoV8A9Vy51K3piIKEPDfcpymis+4MIEkCocFUxGno
AuUI767pUaOXWSzFDVOWaG1jpLL56WgfrRJfS+8XG4vkHfMZHxNf3e2k64d8ZMY37kJjs3luOi+/
O2O6jVTXplBU3+O4uOwLDI8VEpJ/jlOrYKTHPOfkRKOEwHtYCQrf29cLE5D+viEDkTwVdiFVFtXC
srGWC/zZnJvyzIWJz80KxbxNyHsyR1dT6F1IZY23FE9/kpEugtnn9ONkhHKL/OWas0870Hyxpf39
1OibR8wjfYXcIBv2yTJW+KSpxLksaWz1j4re3muACrdF5OZfhDQ4J8du9kzrdi7x1ucZy+MwhJ3V
CfI4BCSsGzN8kRpPCGTz5rm3Fz92T9vp4eNDXKSCuokVMMHFyPFoFpWYBVdrLJx0rXLrA4/MJl72
p6SDqgWuD3g5AYVqKEUpspWNAlp8I2euPCrzL0rnbbwL79JGQQI6lYosW91hHtBGD1I9o8mMDPV4
S9NlHkUH5Yzh5wbzECwriWQQuAozxb0mioUFy+N/SqBA3YYrJj3ZnmIbHRtGhEAuQSri3e7832TP
nlxpZ413EyqJHvE7wbyp2fe8aJ1IdkzX6uctgmExBh+KAswmoJ1EgJkx+O0TKMgebRjv5wwnhQf4
oagLxGxB6aS0YU3sN48zVQfWBCxwdhTuiQ+r8kAZuLmUlaGEvexHmkQrMN6sWq3Gqdcy3plbgMWF
xzkWBgyi0SAqGVf3Po9fFDywUSeXeFkNTuIF0kZ2vCzgOG/4GVCGULildBuW2mZl/OdlxjOzCqjK
kZ2t4dR5WjfXaHijUx+AJF7RNOlAAW3vewvNYBvj5iF9gPLUokByQrnQHWqydu7Wr4s+rS2cxUVS
1Nk6rC+QC9xDD6nh0Kx9MRBVHg9Jih4at/IB0zxgNlVNHt3V7NjJUmtN9ydcim2DNgvJPb3MUnA6
990Z9d70/acOK/7k3gKZEHNH5U2vuZNpkDbhDHsZiaeUY6h2ctYTC/+jennoEbjuf18Mwn8n9gNV
zAab9y2evN7juCoNRuJpYq90ORfgffX+rV8b+It9bBTsSw6VwpSuQljgg69okp+b/EZRbjj5Pvyy
rpllzcEhgQ2rHnfNLJ64sDsQ66QNF/w98sMR2vWvFmkR+axeYN1381wBlktpK4OKDqce7sButhAD
0MYlNqRm0BcbrkFqmZ4KDX6E+jnOjqLjAxybJTmPka0Z/ZnUfKfgbm5Nb3zxrAvCu4nJWfM0kbW6
LAVDWu7JI41MyZQ6XmdC6VoGbAVHKwIgbjIS46K/UmCPwUH2oJ7c3LbtFyLjj3djzVcVMcJmvPSU
CpQpK1zSdzbJFbUxM+Qz1tNIQGwuMyB+xb4Gq3nZGxuwPeKRmse3qIgxSriK155c7+rdZ2k+EhJW
jv7v8YAYixwraYmnVuEzR0B3LB2ZurljxlHYjU11E6YRFtrhCG77AU+ICbpw8yt2+2GVl/oCwN2c
eMmEzrPWuReCiVBS9Qxd35FzkBDDnRCvfGmTJBGymOp+wypKik28k/1OvuJl2DA6bwoLG/SZW9YA
6NVjnZEd2ncoC+4Juglbu8Ycws/LmDFiI/G21TFRG1IDIHz+ZX309FSZQ/vLlTj14NURW1/cIMFp
ZjGVu4zD0rkd/iBfP3IIT/C23Rhk3u+7ODzwrpW/p1nXJZtiYivLOZm/SMhvS8zOaWOz4pAnINKU
b0dhe/QTCecQ8iT1nEzTGu3VK5t+0LT+SBaD4Jvq1/Kc40SQFiA2tQjUoFd2SJwbfv8pMc83pv3E
Gow1KMoR8keebbujM/PBxBsjTnow1bW7vlx7boMzWYSeNTigVxf1JfRThehX8SN5cmI4xb+yanlA
BOe8TvuyBmxU/aMs7lxGoecwog00q4+crIel9aGFOOrRwIvoG+mfQr9ACwdOXBshUlk3zXQdh8HL
JH0fECmMHxUG2PwKfm6XicNfURiK/z0qAsji3hfMXG9QeDrTFhrT5bJ7xOsjyvSHkmxRJiuBq+Qo
NeoJ+dkcp4JxTdcn170KuETsTWK7+I+G0VtA2GNhm2/eEftxPeX3YMZ5mX0manQ6WkyOMM3PB7xr
dvkwoiQrOqG8HxXpPCpkmyMKF0MoKbH/fDamMnriz08vRJ67dn2mGSBYl7BUyaXZgVGulcsWrTR3
WUxfNT39M4Zoc7FHeLs2RdjZZOLCTg3n2w3jefClKp5pElSrE6nuhChDvAmZuX+Alagqh4kzRf7E
NknengxkX36KF7WTMMUl+a4dgCL43QU6cgR0UcPY2VemzbAyPOSrD9FfNFFcXjCKnmdOBbT2S49z
XIZAkoqGrf+URriFZkIJewG/ci0TydHl16btDycY2WGxX4gmrfgC4WIn9NEi1hcXlPwrRkNjwoxT
GM/ocJkjH7IXeoznphhSWegOY4x46+XF+2JgTC2fJsx1G5fq5Up1G2d+A6xMoa69lEQQ9ZKfieCW
F1rEZJIDuE90y4iEkHXMU3aUvHnA8dt85peVQvj8kuqIP32I4+HcLh3ucx3AGe16F6kuK/b/wU46
myS756irWwHCRfM/sR/HjVRRWEsKVe8W0T7u8w5gEZeXtK1AHlUd4ZmQUFAUv1JaUoo1zGdfLUJY
bxyovGqnOAscev32HhEq9IEbhnudpFmZrHjd1LQBlYMC05YEXGhr1CQrgKwK34X4Joa9eMGVpVvH
sodxsDGsOQwUVzj/621fmmS7LfhCqp0QgRlE7d5IE3oO6cM0NGgetx7QIVzAPmvLtpF4qUIyLeei
9U0TrkT/eTzv6jV67IOnfUbTHz227opKKP0rb4aHftFak/BJxdqTo9iks+JTIM7NTrOf1T0SYYm1
v2u/3K3ykjYFKYEd6hkd7PFzIlaAcf1CEjK9cl5cukmP65Wkaeu/No/CLCxpSEcQz1ifUsZoBt8s
S92KaERsRC6e0d5qP/tlaT2cvLgtmOZATDIzIjH6JFiB5QH3e7zTZKE3KW+wQlq7/NJKyHe7LheO
lfnUgX8Km8pKPnEp/00u60wOM2KL70qddGGqDOSbBDYI7hkFDpRjJuXXSNefu7k4WvEeoxPrWw0W
JaXyUcb02ojE1ajhCN9yCvZm+ySQYC75KG1zD2f28nHnkHWgAqwLPFdqstTyc5I35efA6piHCXTa
v7/29+YJK3R5mOoGDc9hVevVxxbEEr8GGWZpuYy+IUVTaBSBCj3QgY23/6qQNvdDpGIMZhf90mQ9
q/03KtJbnKhqJ/ciiwg/jJ4O0BJbVQvnm3GtR5s9E/AP52CRSOHiQ2Ix+6fM9yZoOmmDmQHwO4S0
HQ4bwiKAh9oZ3SELRSdfmsuUyZ9wBOUbhHVVTXkU5PZIap6NbIztiBHRhutdO2SBS8lysuIlkYMg
Sc8evBTnKoljl9ffbM+Q4kYT2ik5JTGfyTbz3Ar5yrMKpkN7ejcIMddYb4wFNxe1lWU0AqMv+9Gp
VY29tMjF0sdOUK0b4u6IyS979ZLdsMD8dp9xMjJIZtjilEeLcygvult59UptiEXbbd0VzkxBYUH/
BX37p2RyLKJWwj/ljVcskyFjPPh0MqwJWX+oI4R21iNEaoUe1P6xyaDXCWE7g/ILwJaVi2JYDiNq
If1pCidhC+jv7OSOUsk1JL9DiwVDn4hhv3ZvB8a7L4nAE//MfOoM3kyp47QNOZYUuSKk+p1cJlsj
zq8J61FCQZud0GvdkNyvPfXbAl9NkmDUxYt16a4LGy7SOD3awOHuyo2noWzKCGhjDls4zt2c1TEd
MBwluC3qOu1imBI6c9iZnL2ZY+B9Hdl4f9JRjakKJALWvo85hP8e7qlKwBUIoNLYT6rObMqp3dVa
EsJZBVv8qcwOAfbWH+rxw9uw9Cf6GjH4uGW5OrRORzhwk7pOwhMCfQF+bWDKG/zVm7CUd6Gw32yI
qNmyLGdHV/xlsdf3xgSHhnuTRHnJJXwJPwovnCHx7Au4JoVm8l4nR0/iRHfZcOPARCVp86Y4Roew
FcW/mFZ1yV1cobkXKygfThJvY0asOC0HhoMzuBAnUP9k6k9dTe+iKJVuc1N3cEXK9C6HEqFjEz8K
0ONIdtTyo9vPwoDWDVndt5RilifQkX4kzY7eGfJTRLwIFhQSeQP+G7W9Fx4OxTfWWh8M1xGVizK7
mbiOWr5Bdd8phB3Grw8ItBgQeCPmCEqFbO1Ht2rqJCGbPtmDTE/VZkDVcwrX0SykQ1tzjStD/qjL
+Ejm0wObOEj9tea92mUsZeFbtRgOoXphDI3EysLAsz+jFfwz5Nj7j1kRxRV4tghoMXuJj+jktqM1
ePG/6QBeDqRzL5yNq72t520AuGGsHIO/rS1+eM4LsDLmMNlV1qxHPlqXgut3e9IVUCBl64SZjRTi
++RkAzkHsPUOyV5fwIjJAfgxd9UXFcmAFRaIbWrex+Kk+B/jEE6UQTO/9ff63SlCpdcaj4MTokEf
cL1+wLvAAL5/PD1GjFjkqKd44wKt7bparqo9kAintU1X2M/CUNlvjmmKzfwA6ATQUBkQykmMHMaz
1Sle83h0RRtbzeoxJiG+vE99BY7dWqWiFBU2q53DuaKt5G5EqqtWkAEHLGXvoqMY8l9VgeXMqyYq
Sx59tAItyDdvF/YCtKQY9TU+P1NUqoWt70NxXXm19Q9CdMz6Z378gVlfHBrYZWJNXfFB0pOS6b4X
IS6ykkepfkUDTxVI29K6TPqkKT54dvdujtte4oSSAYN8OY3lOB2zkW/PD11O/VR+TPOYpFAZDz/g
BeVl9OtXp4jzVWLOv3CYgArp9R9XleZCdo7Zqft6oKm9sp4xzO5zstAkWhHAJiceiCtOZJ2vuAAb
GWjAh8EcCFMI3T8ojoJIh2kbNQ4mzb53AefrxoBwhWAeIM6Azw4hSqTuvRSz2vf4FyXYMlRCxEAa
2jsq8kgMHSeflHOPOdJ8ByRV2USNt1wb6vRpUkowGT25F4A7lvMqagvhrt7bXlqBvOCNwodud5rz
r/Tipz9lO0H1V1g8MidhpxaAS1BUUFnckbDwCfll/GXd4Dzy5pdcj0Dhcp683+j0vJNXU9Obi7XA
rXW4Iiobv5j23bdnzOPJav8/ooUnaNHqrVOzMfXG8FRPfPFYjJNRVlUkLCR6JAQxLixfShUhfFjO
1Z5stbHK+u9f5n/OwAyJ1+SGTeW3xnVqsBDqPS1nBJa+1QmaisRg7cXjF3cmYwiqHGLv9iTaD+vb
m9Mytjyuao41sT/vyQxOe+MDiDPk/gS34u0OxKxLOtuy3DPF1eT3WW45RkeGWVPPpfUXuVUmj2h2
so1IN+2r4ysmslMmvwah7gFqZJXjhyX5nyyCHBNhXpLC8VXtfBHNL4YMngjf2J5+VEr11BB0CXc5
DA9tZmAkRv12IOtxRE79K0rIum3H+WOmRggi10gIDjP7/JBn8mKSaJzdmlpjAoKmPo1fQLI02jzD
qVBut6ZTc/Ran9olkJU4E7NGuDDUKWARg7Dds/BxRKVn3B1Ux1yn6tSGeLuKKq2ORsOuEDuXF8jv
3hvMntQcCf9H1sVf2G946u+EKK/b8IOjwfann1DZca2hU34AQ7a4W3W/33SXcdQI9uZWQZI7cosh
GJbojiUGwobbaC8d0mM0uhvt1i0Nq3I9fI3h7b1RAx3vFl25/OPUP6QP/w8S4aOTA07XI5DYZQvu
YQqFgoAL8svdwo4ioNsIqOk5wgOLbCDvGilkQHMB8CtarQSmes2qWC3TxUR/Rwe/1YqUDJZe+3Nx
EiHFn87zhQX8tGMO6urvKzWiR+WYKDGgcN+gkpO2jIOCVIP507tYXPnx2HsCKCOjWFkZuSnhUz/h
JkkcFBBTUVh1VLollt1RuhSJwPV/Ub2+hUGl/n0V8ZgsvYEEOMy+hNgQevXWeQMX7gGlmcVDCl3J
aPSFrPg/nYcAXwRv6nnZDzaYPWt0GC02if80eViWLJ34u4hEMhCMIzT+v/2auuLlbu8YMddVSbLE
k4shl5gCYV/H7zaXljtaVsccXf+8mOusDbDV2ei4Lb9c8p1fzRYgpdbnbfR1wAEwXVk2V9DaEQb2
B7GNaurCK/wn0YoaeM+cIwmyf2FEaCHDL4eaooly9ynEGUS/zRRfVYj1ehTtt0P+aXCjbKDaVhjX
Gx3ceOrzCMEeEajqNU93R3U7yr43fiVDJu3pySrpfrlyNNE7Z9xsd2Vj3nIVt2e6E5TBh788toC+
ICg0/hwhLMV+DcWzu14CxPfXgOnN/BrWJmdJOkeYlAUqg4J7nC0w7Ezg/GFc6HCJKlF5Xx9KqLEb
1CIbXZovG70hLCDvhyysieRnCVW1VWNxW1u4CoIDw66sGKBtn02Bfm0cVG2lzi+WDOypdjq92jZC
FCXT2Y33B1GKqqxIdkBOe2JW2MKec3ZVjRtrWoN5rlDukhhkrW41Nr3WYjdinDf9vcqmYLyMTRok
OYw7sL/Zj+iFpdH5ep22/MzYF8FXPavDDg/atZt2waN5m3Ou50N7t6AQExOd+dnoWi18GKgNYKZ1
NZ87X1OcQ2+sU1FRvx/9sK/D+wyiglkNMtpHwo7a3qm7ofHmTjBt5LFy8Qow5rSnBhHkV9SJM4Y5
04DkWq1pELZBYFBuS/C0g2hLxnNA5wH40BblSnVfapc/liiumlaCqe4FA1FOrPFC6UDOkZPFk2EA
yNn7izCWNZXt8ZhoEHO1UmGEP/P7s4Rj/wicfF0XYqnibboBxTZODkl/8n7T5XtiJoucq7v6B3xW
yvhbA9SBfyPtmnodIeoQpd/it5I5xtPlBzCHkWfWqbOHlKnrwo0O/jM1TpOzQzrIIc/Aw0o5RgD+
sHAHgPoCbDVaWHB+0Iseh75zPCECizMfgdL8r66DMI3/PW5vco8uuveusL67re8RuNhE/Tt1voUm
wUnjJn9VmX6Ij3U2tSKgXORdkPSlA1fZKKI9ls9QAa1amXbXt4LYniFa7yT4538EmSsgSqPaChu/
OcjPIa7aarynxGfmgzRLqv3Y4Ecqq43DZ3m4WZxjm/nLYO5ItQ78vBboHHttGSrjw+oVksLEEsuj
iZ0SWfsPcX7TN9+Vwyrx4Op71X5oap99jRGCeYsGRBM5FI8mj8lS/FE1ymBCxZp+xQ5wEkav4APk
qRrOROy22xj2f2qbJzXjom6WST+Qut6IURke8CFPfT+O9QWWSpwv2dPEp5uNegoKvfPnnAa/u0xN
tGFFagYPAkwX3iC7p2nEgoQBBSl+ytgQF/ddDOoEB7eLVHYBa2Vv4nPVdQZt8c+N3w7OoT4PGrYv
9nuIsgEEpqiYITqSiYxYzUePA48masweYK2YlSRaPclfk8ZhFa1Sq1rUVzaGaHV9dR9VEMnp1Nws
zO/SxjNM08/urH9RpaR8Q1nw082qR80n2UaYSvK3JsamgnOzNCKabCSeN4uj9ovN0fugUkjRcaeH
J2NyWzEAeXx8QpJRm97s93Liua4LvtlhiX3oQvFp4MSBcpLgovrceAuhQN+02Y8vN4FAlYQ1AmW7
Nzi6DRWAMhtJ2KkDH61SvJVklNHsfvzroQKcT588imUi0+ov4p8TVO/YiXhjDC6bTTzv95ZA6Tvq
nkQ6AMy+SkcKqvnbzg2LChYE26c0QeQt5xYp5KkHAibq+d21bjsvXY772i8m3cfPCZ4rxCw8MpgQ
3CteJrcyqdDiQkpJWy1GUCCqHE1t5QPADEgn403AbztJCbUyZy5PXig+pC8rAfwcyiHJO+0uqxPU
+cwe9wgxJKWzNY6dARhdeiw8nvasORwCixg55UHYHPYU+gG3DZ7pmm5Ge3awLNNlb4iHWu6RpFJ6
4D++7nurDdGnb45s+nPbSzi3IirNAC6lLsvnFeIX3kgrqoadGZXXo8f85Px7kuSrvcXN2dSpCKe2
HO1WqXsqY9On3AMxenytfU6Fe6+gcl2gFwu4vRXr+QVECMZuzpaRbAYpmVrTPPSetAzPG9vVElh7
6ArxbEQbkqiL/4EPqEGz4B11AoFFyA2W58HysSWptG8AO30QkUspREykcxZSzvRpkU/CTfTcVCAg
jBJkLJdrwBxUGXnJXmXpf2hoL0G/4CZigQZd1aJFY1hK+lpoeaEWnrTRo/eBnHPDNkdZgbu58GlK
4AoYMF6QkfhHsbgrvEs0+D1gYP5q1Txxq+R0Ekw6AxbNHDW/gUjC1DPCFKrfoWytmZ9+a7y1TKzy
zidVH5ub5/ay8m1NjlWsRSa+bBLKdzYWvD6jmGnk7sOZ5ixUal1uzjejvkXgn+mEBQFbBqyQ2sOI
3UEDeHaoSNna7VQmVN/8JBjiN1SBaeJXkFTL1qkJHObEWD/gMrni2RuhFZfiAi5fndbykAlUiMHN
J6eEsnDuWfGPmWCFu181NiNNE8C6j+ajjp2gpELdEpPDC5aCLXEt3jLaS3NaXH+r4mZwdCxnqX7+
3YB3CSEKLYplboJdAj9Fj3KxSPGW3XCeXJSQX4P7cgeLp20j+bCM1mW5Rfdp9XNd5BsqABA7zNN/
JZxYr/C83bX6/AANS36Ka07zccwzOxWbyJobdwTpdC7yL0TECaSgvBsO01Bt34DZmvniK8LqP8+g
QyspoX38QKw8uQI4N4oltVClRQtXiwVI4IRnSbnjlML6qQxXqxC/BMRiG3xKmXJ1IEmxzKIuV2o6
nxCNSgFUFEp1LS2Uzs7C1T1ckFquYzKVS5wDZDc4fsaVnbmjQATMvn1WoAgzaAZPcgNfCrLbFY+Q
daSNT85cCBKvgFuOjhuPFkL5q48dx2Pzrv9G5wekCbSRwW+jKwCNvCnko44EoIqpBmJMF8R407I3
ysiXpbEsTPhCCiVTXfPjyOu4jvlyWd6xR/jLoesbHX48IMXvZ1ZL/eMvUzmdqpd1sWOuaXO3Hr1Y
9LfpYMkkT6vHkMdAoqOHZQucRTP41hfryzBM61xu9VzUTeOJJ1DVeGAMe6wpqAvfF27fleEJgm0y
GYbEDluk1z6ljs5uvCwRp0CuEWTrqP0IeHE0Ddl5utWZfO5qpZJfNznBwEUYxb8mvre3YRjZEuga
q+/0k2hBdh241VdV+ZIbU5HVmGNa57lU9cSdV+SKWBhHSqRfIYCfxIOIdtWjHq1i3ZKpdZuZedyw
nZYQKh1Uk4dLL1nbPIc0sBHcJYFAgcjx6P5AbC2FvS56HHtHXVXLah0n2oiQV/LbGQtS0iT6yG4B
MvK5wMSynoeB7WDjbxVVQE5gMqhN7+NJMfYcrdi29qVeHzpUYowd0+rfa8LrW/F2MPttnDZHbKfM
5EoCdOALE+SIOwq5JKOlrmb32C/8ICI8wuln64liFOL3DX4+DV/DwGoZPlHSvvVGrdeY0aphHqXq
9Knn4sfPtdM0fL728tnlc927un+5lzYBff5ffRBmRfjTJ76cM1Ln5DIX600EPSp30sLNcgMayL5e
tfhHmjCWSzSHdYOze6R1643Mrt6ayIp1NL/gczzSUmEL9X/Fpf73c0YP1kaMH961viSvJkTmjmvu
B+qzcI4lIn3AuXV6XYqa+H2DkjUubvm07xuoI19MKdlZbYwatMtU3lqdJfgE/TJT4lteg4P6+p13
P5pXCSgSbaSo3B9UbDiqywNUFGamR2ZFxVZbPjhM9bidEvgsf3sr06QRqq17PpCcVMiLVbx0Ve/l
8TkmCFRWx5fROp1tE1WHO9cik/II5hCZRf4zAh8iFdk7XHyDhz3Suaxr3wnSAKaKId0XqQiu0hob
Lg9tBJ2IrLQU4Jyvy1v2zWATP3eTxHFKiNO9yJCH4b1/vd8buPCAE4g6Dop7/MXeHVcWF2O+XDOW
2IlBP0zEVrZQYQvI/NDMDYl4bPprJjds3Zto4ItiIW9BRAU9HQLpwU3n8rfc7KvZOz30CNLZE8H1
IZ2oJ5vKGwItT9uKoo9aPNNaSNFYnrtLnpIVQ382eDOWqujZFThwPnFMICVzBk8HqYWx6cKqxS7q
/h5YjEvjwaupOZGPgKtYT6GMTR8TW6XV3CTcg5A4qsYKph9hSPesWNBP2rFBnNYkD2/nKnJykFn6
cpgoE5xLHiPBi7vwXyNEYw/q54L0oYyr0wo+ZnIs23RRb+dqnWQnf2ACJR0sEF55GqyKcd5NlN9f
Qo+xPLpp4F4RGSPnJ7TIXJhFTOCczYSnSVLf/AfAzKXPLk/Aa9UV2g5VCvb6HdXQDIFPvsjUTh63
UO5UG9Uo/GdqeI6PTWATAA2Fd1WLSa6BdzQeWJD9WTytoPbS2HMl5pFLCrF0Ol91LMvl5dNzxyif
soNV8UWQ8dX0WJjVyz/z04MOtvAjpk2LLncTQzcArq65mgkEhxqsrgHTdl5yLkTNjTT4zyqCfDuA
S/nPiJm7hPLSQUko/qObXKniRwkilfSPOr1xYsazUkzEcxoftn2FKUYMGtzugvh12AyM8/RtZ+4P
O9Ii3d5OAJgayCDb8Zc6JaHpNwdzme4ZYoEXh/5RuREDW8AbT01GnhswdZawAvS0/BA8k2TvnCpV
04WIYLgXhJCJ7nU5z72+TU1pWfPDRrksShTz/wZnUCUP7yLG4N5Y/cfqxbyWIFxtxuhOlhn0OfJf
b4AN1sBYI/6SQfdEer3aniqPuivDgeiNUmNFauavGyp1SxGGVpp8Z1aWgzAqwbw9zTGskQo/hMil
0scowExMnCTOfXZLR7pXjQlyiSD3hyaEjPD5ugrtPcB1S+Erh6hO+aWp9Aa1VH8e74pUqpI8cFkw
5dEmf2sNnLPbMu1A56XPyzSDvDraREpcuHsrMHI36zLQZOhKkIatWZX2KXNvdDaH30g76XZ8afdR
0JXyyWNV9Ik5Dt3Y867/WyJmPm8Fw/DerqIbeugDs08hDhH5ll1AnQXZPZuCwvz4YZ3BN7uNpuIx
nFf6ViVs7lk6BonHyw7RtwJCCeMkHevn035HyDLdDS2tgD4mbpF157d+Dq5KfpKXY9oldsLGl8Ro
0EY+/UeIT3mJLUkUjri2tfOLywRpHaNiz7sD0yzMJs23xVFPAB/6qvDQzhGwClenoHf6GrqLHRBy
10Y0rDWAcvxsX1XNyNaht9L7xV4zgIWHj8GQatWd3r71CC9+KPAIVrdQmdBHFk2xbiAgTwUS2WGb
evkuqIhoG880Bdp0wDZhuPH6alPNwm3XZDJrkqDjH3LamY+NjDKEZ7VracvHbFWr00brJj47C7TP
se84xbiFUGrSVrbsXOlcQUVrSMdkt8cocfKgvNgmiHtsuYa2MjFC5d1W94i4KvNqXnA9dQrqlrRF
+hNjzJe2cZJwzETpG9gx6mGjDQjGcMRj/oVpSFx72CrOWFuZy6p6MTahfx9f9YYOZZN1LmsRC3pI
NkN8COofUxkG2bgferE+9+uJ1KFaQhZhTLO6hkngluJKgfons297NgbgmiJ1dTTg8ZkuHxRcBFH7
eLJPEAU3sK+d7wp30VI8fM1wK/BgaNLrU+BZN2OMed04tkrTt3/vX4ZS30qJX+csHo8PXsuOFBN+
w1NaC2dDAmMVPxyx/utmbv17OpCTwXt6jij10ziwozYJibn4FfVZIpwPUNrJ+dMalEG/81Q2B3r0
c/zAzUYBSyqfZ+g4YHrOHO/V0U1qRw15ID/5q2MtSjFhrwvKFCltxWeum1i9cJV+cbwCWwRtPavg
pOhzr59eKsaRCJbaE02THAbJwOGrIrrKRv+928IskJRIggjSmnYDlM+vf0MRZ7zOd6jLsjwee3p7
RB311/4+wtzgn6WddnpJXGZvsHpdfSABNpBhZroKo6n33sea8I4vEUyOyxQRpUbirRsCI2eAwq4d
zNfLpkq+bMK787pnFqrZc0TCjFMik5STj4ORT+oCIoA+lA9sSv/z03hf1sr2TGf6kreZYN7bV5X0
SLceJ3hCVRq/INmpg47G4r3ZCrSvGzJ+pPz+CfR5FjGRGCpoMlaEJCF9CpyiPfSbOMBChgaGEwYm
/Tjm9tb1DFhpRT2Wnu4dpmBuCGI75yK9V2AYh+54GbvqBZ3/4TOCSD3oVsQO3za5i1ALmNjYoTS8
Go352rUAkuUtyUCegISAREbXZTHsGZIGPoFpt/EcHW6d659sJJr9av/GQ1LBkeUI37UPIK7MxZKy
1kAxckNx98MMDIhEOwa6y50IOZEr7gmxOOvcRjowqMVTrzUZHx7TsloL7v/9GOC8ODzUhgNTNQ7p
eHkDxRlxcowkOnGeW3x4ARTGLzP1a7mEX1jKYF18DfWyO5DcEx4uMr4oojhupJ/fOtAt+YkZvPmk
AjYsi7LMEiEwauyIts33fe7bcN+/hm9qSPLXPHQIjC4w3nzC3Oi29uqvN4mfy+PvqX0XaowRHid6
X0MiblOIJMFl79cJaoWqioc6D6tlAKeykQGIY/BB3+S4padl3mzSgLvhI1VJvZ82fGyApVUI3tw9
4LOVFimDWkl2GysM3pE2xgfLYTcp3WhbzjUY6JGzapcIERcWhKvfrAYA8YZwkFO/R2YPkXvEoe9c
3QGhn2a67ZfInfEvwWe0UvQnXqHInEenDbm+2pf3SJRRTySeAX2c4MA/hZtmGjnTXw1kFniBvwGe
A859mEPBNwvCK/ftBA09BqacoTLUy9/cGOtDKsGvEb19NykyBQII/7Dg0OgyUouC+zPaQPXEYaBi
6v64FKdXARAoas/X3ndz4/jkiGhEZDRvY03ByjaZkJyLC1MQTyctZ3sWKxlt+sG9pOnWdiNv8YBT
zpvtNYjTRxRIfj5INnlC7asYl5QgPf4a61szLG2aRUpp3zeNvHBdpq9onB+Q+xjvz12HCsC6n+41
GdweEGbtvL0uW3iHY4txC2uPvM/5u5jiFdJ1Njg3/IPnb/N4hqdkmXDRTp+PXIVvFJSI+GVddCqh
/hG9Pd5hxz0SsBpsdEDb9aGuyczro7lbDFF9IsxvjQ0FArUL7X/l/Ynb9lpaaW0UYDm9STp0kyhZ
ip1/mjgrrKbdZIQtd1e1XBkSpKGgwiC3xmtCrx1/j7ZkfwNzRpgw8qx4e1LiXBCTyUgcZvfOelQO
4NISljCqUlpR7BRPHL+W+XMUJW6kdoGoYh8dZsfJnIGJ8pnWeCtIrFwd4kMeUSWMbp6Cu9mcGtm2
dZlHFoV4Lc6X+6iQ1dUcsymZIt0NI+RGaqi+zTie8PNMOA72ac1njPv74ZtzWUhx2Hr6/NMQHyIV
wy/ChEXnfTDJECtKtmsb3A+0cCzP0ygEWnvwld8kdBjsA8UdsURi/kglIOncCpBvHYJ3tkAI0csb
ARBZPYVD7mkxQnGjm82Ppxrd3QrVy/qTYjwl82eXMdvXPjy/i9Kx3+8DZiWPJOB6cIGIhlTrwhf8
7X/cs/p+VhejRiye6VvhoTEkq9tkljssEf28Nc1TvJdyCOH81ZJptg59f+9UXh7zFovhWHnWHO1O
URxD1nwXc+s+0oRvUCvfMhWmi/EMzXjWvhYJPxpMyrCIrcKnIvcwxhoaz7PWHOfAunutUw3jV6dx
PidlQn5fSTew++WuvUBDy6fDqVmS0i6Dl7GUyxbrcMzHMOQPLF5iQABkqChH0d0su9rbSJA3V2Sz
cJ4ycmmbg64ZLjgkkyvboSpf9Y5ZQKuxL9nV/sXSFl0rN88jBg5c+S/XSEI7XWdeFtpuo0j87n1J
+flGLBOg6L+nUml4eaU1isX/cbeAYQydfXyoN3YW8JR7+2bSlXfwVL319Vycv4Y+3U67qP76SDJ7
uJG9y3Op9JtMNuKQQhfNZr9hAdnQ1e76qMK0VLfIXbdPeQoqXaZI3CzOXQiTKAwx5Mho2Ek1pluL
4VKElMmP2hlr0d6eyXUyBp/6LILOs0JHrMvfo5WsWs/jI91jB4v4VK+3xUJZwpsXqczOJZsEU6JY
7uH5kRYGGZ/yuzzopwMctzRNyFhd5InAKFp/Q2kseSYpthKwCRWxw1W4b4OJ78enH6zhSJphMMbw
FKDvBEtDNuplnYM+GhpkUD0sg/JnAFqxTJv26VuJCz4WrOF0qiT4Sntkj7eqlvwWv9bJffSTkexf
UeZxcTkEkqV72MWxfLh2MWfeABFwIF8dpPcZYpODet9pnjl3ZWTEbRamiK5O9KK/qdaEq7sFvDQ5
4uwuIH+u9QWLiNkhfUMUZh1MjbSk1sGlGF+WE7tEZxecvzuYcxq5TaR2bBP1RpYMk0UF/VwuctfY
iEVdT1C/icGBgddOQc/+gAMavXPO/cl93Ba+5DmPZ1j0Bl0SM1mrAAvs596d75EVA1/+4utetl9e
r+yZzW/FcmbBhFdVs4+MJ1tAusT+IaM8mosyBiVaIE+SkSAVN1o9+bq5DD/hcaZHR8xHS8m4XZIS
O8Gc+d0SYjfRTD3f0hTrHScdO6q2fTrvdR42jwjVGbTRnWs7uJWDLjp3F2h/Zcsl4HWZPGuPhyhh
PUaDn1p8zSfd2JE3HWKrtKrUsqeRMLmeHDmIp17LyvKL4Nfhd/20rVNqDzYEcPunTMtc5V8S6sck
dqGzOJJO4e12bNXr3fJ1djV9swXhftspgiWz2j5yglbEbrfh8zKrz+poKg4IxyP9uLXx9Gkiumt3
e9y0UBM0auVnKMsJFmLM8ttBxiYnvDNIF3hiV5e9dKhawGaMEiKfe9YOJYkP5FWzwhU7qhteMJbN
OoNP6sTFpTs6KFQoFjib5Xhg9xINHsMZ9R0dbh6anATGyfDpmTB9AKumQIhegqpkbJoT4EqHBmeX
pUZLbmGiVPi8qkFpwoCoWFMn86QBmzVNp53Zxh2Q8XoTJtORIuatRYv0rGAxJtW+VtlXEew5iSUV
NjGqiopvL+A8Iv0Inqj0NvQ5dLrWb127sbW2VgPVKuGWiuxc49si/309dsRmMYznXi2CbZ1zQOWI
7IhCSXq46pbW9ja5K2TQZR2z3ZECCQ5aIs9i9nJMQzszm13rhrHWYUJ3u8RXipRXm3qoYuh5OLUi
rhHnYHGf1quiuopInEM623/ymhOsqfaL0HJe3Vt+RfLmSmX3NoR1BWS5ejgQTaLxfx3jw4ryE74R
LWq3uIkA/iw+YDQOxKSjrRDNVlUNdVNYKprqMbKXZtQIxqQMz1pokagcafl2M8t3FE5leAtf75Xz
loIb07K/mbwX5G0O02mx/qBzN6HH/x/FGYp9QkP4AhX9L/dnEF54wLOIqgXf53x+Fb723IAtsnH1
7Kad6RkMJ+J9bGAti4xIljfdEtQfFSDS6l3yMRqnEGuWln/FjUjGfkkvwoxX981CfbySMcTVw024
AOYbNsxlbRAq7ejSREvNyKCG62LgNwIDk+1HSXhJLFonMgWWs+2JRjciaIS8kkI8bf8ksGYUON/e
gRx6uQ5mP3f1dLAYWVcAjfm5OP/Csb/ikZAaxCuNWaOhXydLzrOvawECpoZQSMFSePYzwfactpQ6
dEGD1Hri0odo431FHPS8G6IFPLyheF4V6T+gj7u+OZlXIGHo6NpvLn0unBTXSt5/vky0545thWt3
9ijhFk2HXE2a9kH0G+Lr5CdZf3/1mZyuB2io8gJtG7gF4QTjIPsIKRexIkI8ycMwE8cjsr6+8r3f
z+03Mr0Bf5LOPDKzuInF2qyxZSRcaGHbB1yLOFj4hOMY3Fbi8ZHSgbaO1MHks02uBHojoSJrqN45
FobgFqQrN/qTqekHOBy/IjSqrjKmNQv+j2/uqiQ/u55LCpR5/veUXMsYDA2Kda9MW9YXvr0CFAY5
PSm9WzL2NihF9qhYGHoMbqNcroT69ClCe3eALpfOkuLn9wlNl2o3E3AGeGWBweQ2PfdqlQmgvb2E
zP24jsTROnc9KBMxi21Ha6vxtXIzopC+XynzE6ywlGvaJH7LKOMReGyKH8EHB1nS21h/jJVPKNKb
+RTzCG1AoJxb9WNtWHh+L6rrqPirEY7wpfbF3ZddtaFui6QpAXnM9bif5cY4291dafUpm8BVLgkP
lSASk7i7bBhX9kEk912jbfD4PCOS3pzBGzfJG7Zf//0EtGx4f7UMXkwovDagmxCoeqmJCl/qEmGg
6Uafvwe5NKRggySave6EdQoqncpIst3SQuqVDYAiAEGZillXgsuyMrXPJqv+a5AoPp4I0nC/sHtf
Lw4etTwGDtEOSzuAxKuOAsSJzwRWyxkGzbZaOOJy5lLYxIUxr6rG5bz/iXRjc4CHuvsEw7/fRmmU
9c/mZ/bD405cyi9xGoCT2QazCpJtlmYtoAgGkVvEqCqCxSvpu3+aYnejF9ZvUCJKq/IONhKbBLig
GCLSFaJjNYTllA44DVzsuNvFwWUf26ETBs3YDMu4eR9Ct5TlEIpG0V/WN/uwYz3I05kN01FCCAwd
lpnx6shc4TsKTJcePPw/ZdRN9I4xJpag/P/IKRfY5i5BAw8d7bgbQHiNyQgd0ILkmnW9XcQkHve6
aYnbfEGv5ikG5bIadWReU49J9+X3RrG3T4FhWL5nUsIqiMkBST7IBOR+wbC7U/UhLdKZgBoHXliK
AG5uXgZaegFnJK90gKYitVfXy0wJbOszFRiITnUNdDhuJUhtyCd5BhfYEZTmcP39UZLQmtXQ9JHq
Q1UF/PHNwaX0kVZUBw50ZW9roQGqV3seaPMv9fAO5vn6tYFmxp5SBRctNuJBQILtAbtd80hO5z5P
2DrYEsd4PY2p86TL9Vi7z4klXEQgo58U8jj+87ra01ImQB9KOKtwxdr05fPXW/mQNyXNndFalWP+
vuMt0/ROiX2QTV5o9LCnCyEF0AW05N2kzCp0zso3XjsGJ7KyGyb6QRie6vgRdEIGVLiJD+al2kaT
C7191Omh5x5d71I/Wkw7Bp8A6a7N9EE9VIFT6CXxZbEmgM9Fy0W7SSjydOkmPLiWxvU2piHU3oWf
XfqTdSCB5Hati2XqaeunIbg31CfeNiYipWgGASjinxfeTXUx71nDWmSkg5jrAnQVoHurMgOPaPHf
q6sCIJJxphR+7QGrRh8xSvSXFzoAb2mCclBvBTdQ1bC8EbhAJ0DaBGWy5adkhHzDShhsI3Zo6yw3
vntIcpC4JsVbO4ZKiMUHVGYgOoqGro7EbGhLZ6pbyL4yHV395w9TaEFMFXJZMJOF33Wjc7GR7aho
gDRD2wRUgMi4pzGU1m58e38OPw+xnPDOXkkxsgxxrFaa68VnTTGK14io/zrFz5XUh0XXfstCoUi7
BOU+UQJmaPwuMhgxXDl4cFATpBmEzgCwErPwHdG+pED/epVVqgl6LrBSyWZvAZ4eN4jb9L5MR9Ga
TAjF6gQfw5SgnBQV015/10nthRkf2fUM3WZCk134Keo2+6vzyC7TYw035LcmTNfNxyenOi1TFtMD
MHHmQtaHTPv+puGc1qBDkYCvHKWg6JWkXxpuQCDh6vhVIZefBOIu21UumU6P9gB5gBi7Y31K2Zqy
EwG1PgehK+XwT17PeXtGnik+NZEOWIPUmHmCWv/dMoPKWjOtbUqZ0LaZyKdOEQwkP5SnTWWbxEcx
Yh3p1t52j7jbDvT5/oKmIXxuweugPbxN6/tHPnU8Q2eTOwPJXI74SmOzTtscdjAvSqoL7/5Pmo6C
yWZr20kdHuKQGXrdULAEIlk4X6fxl2jox2E6j51zNskqjT4iuiySRNl2KyOYmVBspwoEovkqHB5b
rz22QXnCDQE5Up3u5NU6YtYAExyQcrRLxCITzG7RnPV4W7g5j8tufjna1fuhGERRE+4Vq7MjW8+q
7tol2xnB7Q8vANfKT+Pln1edw2my7e2a7Zbv6VcletPj3tEzfeJCtboCqy8Bp4vKNMvzglllEv2C
pJwv0LQaWtooGmuIEacpXxM8E2aIYzJTKu2761zhESHFWaMIowGv5dzYLWXhba0O4SwYDgfu1E/k
/0ux2BSLYg8/qeqMsBXl+OKHfDkyp1XgiSxrTKZ1Q2VdKc70KsMHRwI2u2sj5a+yrCyXQh0ecNkL
RPNv8qxbTvQ1UZMxIrsw9s653I/M7J9H01dR1tNcFwiO56yIjWbQtob1M5ydUy8ZtBgq3ZPFljhC
OG9dm6saOachuO+BT133OT+l1bqxBXzaZPnrDdj3alEiPYZgMRuenKOhVLXPK4fIGijozTeZyHSe
gzcytiWKqcaaXe8QOGojWIFN4Cv0tRHoFgJSiwR23+OdZz7E1Ky3RK4h/T25cMn0oGLwOqlStzti
cjFzi52djL/Ism3e9j3xrAkowKkcIddF7ClygJB/Qoi5byVeDq3CoQqVMnFGDoDtpEiTEy1YQbiO
cYojqmPVxmbahIVucBsL8DZQnSrqeeq8VwCKhDXsfboa3JPepNcjOmUdSjMr4JBiqspahCY8t8xi
LBCYr8Uh1HEcHLuyqIMGDX5PPmP+vV8n34fbXQCX3bhxN6YpnZsDvJR9g6OQkB1Ik2KFFxvWyBOw
yP/5PVTTFpO19pyeiNKtVp98IFEyyj6paLRTDW7TyXL5gKdr5ZBxSJb/vM895hp78Or4cDJ96U5C
+cyA+UkrxCk9mi9cQ43I2Ayi/p4SktplEp/YqnFdXSd65nvM0K32cBFuDw3yCowIc3NyCmuuvvIm
56UOSuS3m2Dl0CMrb3UNnDGA6tNcXwvrXITJKTstiX9QAU5XXT8ZP93IkGBx90YQxTHP3hO9H76I
YdT+oJAXiMg6ObP1kBJBuBeo2dwBVYAe80zhm6tlY28NYqBUcC8xaZm2a4K0dIf4XLUksW5riAl+
wL3hgZT2hf8KRRnEwvXsbHLKGOmOfteMatZ4IdHdsHJ8kle4O0qPKVKjc27bJ1m71jH5Dv0oec2d
A1XoohtbcbwJDjcaBoKZuuXhP0UMeIoZ/TStHHFur1TaYuBOmH2Ud4FJBvV24BhqFB1llrTKYNFV
OpbdfLrazSE7bEVUtzum6gFyVrpomxP56MZlIGLQhDyqrXRR2rlyTfXxDIaFzE585NNEVgpH+DUX
2C+j+jFSWJbf9ASyIk7evnMLuB7I+S6T6N1johKtiiI49dd8JVLHSKCG/3PU0Cu1mhn8HIxNBZ+R
27fJig3DQcLXbg8lB/xsYX4+hArkUMc0miCwJueuzA7RwVOi7aggxWmqwRRebWvjW412mJbmpP0O
A9OeZTyHzIH7SSN1rM3judZ6JB9Z/T0WtEMrSgpS0tZXtmBYfqMcyvTmc4A0Xm2TONiDKkrmHgLJ
0crwBzhOSpSXW/88Vg2SHUChPP+K/n+C2xamLonGYbHBFYytOchUk74d88LhvK4F/wfKSYyBHfRY
aDdB2kUyJ0fsLsVsC280k7PW4VspJG94IvdlBBmUToUSaUKME6h+z0GnqfLR0KmjXLV62yGUwu69
OwrKL2iYU3zno+kM+PZD33d5+RsHC34r97pgetHFvoLgdK5xQnlTvv4ZCPwqSN9f9ljye1hKghVQ
w5mlFjqKuiVgVSfS+VVugj/mAkRVQG1KDQjPkyo/+VEE8v/TGSjZTZBTNA6nlOBrCFIFWO8O5ShP
WTTuadUI1d9YOYuVuRnzPiToZUhR+ow2k/2olUqZ8PXzbFA6jE0qCp1gxtvdju0Ta5E/Ks0ewDkZ
eg5F+KM7aeX+t5U2VkaXfyN9ITi+l2D8Z9d+76OzMSs+wkmC34ZT/fPTC3ETx/MOpbtJH7zxY84I
2D+UFEgson+0hA34ooTN5U2PEnE6IrDkq2Pp58yWfbTn074ew4AYTox5uAUMQPMQUCOhgxL5Sj93
TUU4eT6MnwusCHb7ukUWEFV3kfZjABT5H9kJ9qhWLTT2FcswYJ+zBy2qIYqLB7MQypHyzxaIlLyr
raFTSd4XD85aemw3z48uDHpiKR48P44o+vZztirhk2rSzguU4pzipxr47tyqqXBW4Eg7A3haYrfv
rsDrSSTZEHOgv2QRvarCUZmuTeUEpOAOHEwr8LFDrl4QtMR2ss2T2z8XExAlT9c6STd1YAZuLLYu
6rmtiJF7u4I8DJEx/LySzZYfV5k1jAXUW14aFWQpEiZ4lnHzKfzPU4pnaLaaxxVbKhBCIOTCFf8I
xoOl7EjZtfqb8A+kqQnuhYSYJEZQ9gYxu0iBzOrsmX/Zipwg81zTBwEJ91DHVWwslNuHk4T0pEik
DXJ5Z2QT5SNe5LDc6Ey4wPjvErcdaQyJ8HAediaZb0WWwzbVr9WyXVU/L6LAMnBvNt/qN+xb3+p0
TcSgZBqk/94IWvoJf6u+rbMv+9U75mAvJnZeq2K7IzDhkVeDd372oxR4S+uIL0BjgIJdrEqPS7Qj
efsNz1/rZCwQZlWl+v5RQnbx7PmpMlTm9hwW2auaiA7tIP9xFJOKgH7lupqPTkKEdCcIs3pbBPE1
ez+cneWcPQd70+9HBU1YVyMJbBu0hUs1JEPPqEDSKw3LY6bI38Vb3e1rlSIoPRxY2DbTYwjV1pTP
ZWjPSwaTN3CTZTGHXjNUfaVUiSjI8v8kW+DCeMEUURHANKKcIyxAriaGEYiOkaX8YNhF35zcJlug
JA5VpmWpiGYTCYFfUfoK9EFN8uMtP+GWdy6TlB5OH5dypU2EPKTd+Sha2/dt2KbadqxwC3YSQLFK
q1DF97Rg6K+4kEnDxI7wcl0oBvMUPDW/60YHsgOQEO5I5uuJf5jQzGs5wW4w3RP+H2vqEZofEOnj
BuFhWxKg076Ycqtskc5ubYDnjo36ggCs0WtNI45cVQxi588XkIrPv8QHb+mCdcwLf4lTcVYrNJ0k
riZWgJVg2VvWjTgWecG+vg/PGL4ZK+pBzDZyGzulDfQF6Dsr+NzkmPl3KJJ3njIDo2k5DkUPA8i1
8TZK89zNZ0KtNfpJfC0kMFFYYHDdlkGNx81Z/7ft3LfpBmI1ppX0hGUEinxpFhVT1SwFCMd38cT4
k8E0Ijcsep4gNXPW3CVtdNX6A+TNSK56LYohpnkvdpBGUPmaqQhpwzcaZg9rZUFm0LO/dudEubOk
HkKJu3wMeEoXqLSI6JvWvEWp7y/UG12ScKSqR3U9Lmew+El8dihl13+f16BMghVIAk5Bh/1xNXIs
pxJlbDIGMb4SRIZXg9ksBrrlXm0XAeL621bNIuclDsnQ8VjRSGMMtTAp/xyXwirbqptSOIcRhyzO
BauA+JdsvKFH0x8pAdibDMSQ7mBBGJFGDob/K5owP+jC0VWdON3heW+cD+jYfrfbNoJeTAnFVp5x
seZhaK+mQ2PQMPLOcJz9UF26gQC79g9DIdnht004BZod0Iqa4gXV4gLU7xTtikY4qKgGneJqaguA
3YewifpdI3imkKKPsODVMsbfhkJKLy18mDj5fGtCN+b16kjVrPeEMALgd4HaO0DAaAASl1WBdAyJ
mf5N0Ft7dKpv957PvSYhrLnuAI/6l6D3NnKnNgb3aZ+0OfIsTU6p/WtTZN+HHuy+veSO1wyYMIwQ
fxn6sylb29GLixY37d6HhlnOTCDtHTBphROCauI4eKHEJhvQclQiDr1z+H+zfyStsrUu/rETtag7
bx38KIJu8npx8dsFXwbT3rW1mmUkfpnqEJj0Epi256p4DdZvzFvWZ1FPxI1xFu47crS4REhepInc
pebjaAyL+gINZm34dlnvEKzYqLt7myMMobDpm2WXN87lVOn4BI1Tgteoo7QcqSxWpXV59PkXJjgy
GWW1geHWTrkXqUy7/Wk6DfBq++pD67A3MRjq6YZg9Q1jP96okEiah98V8CYEbqkXhoJ3+EDVuToc
NJ9Yt7DkIp5ueIK5i1KqOYcDIuiJBlNfc+xT/hwvB0c7cP6eYaqo11GGoF4VZGjDK7/EetrTYBcY
ly+d7zlPU2BEToOCjfuO4AQqvyDbj6AGNWrHbldKoerJJJ1xXmZPeuOJPOk2R4mXoxajR2tWMR8L
ZqX90AVkywf4oEKH/KmdMiAJgW79KQZMEauDVo7LgH0EABrQUoYbXUdauzmNx0B3MSogeIcof3n3
4BSplZltHlazaA4yx8HXXXL9lS+t/I3Nl/B5gIBYd0sbbESsDmyAAsdxzkX/CuEuRBsUrnBa1vIj
yOIwHtbrEyh1EKRviRdwu44kL2MXYQlHfW8S6TI7r0ht3Fz3953UM/8AE1rwfwOU14F7xD1Dt5Ty
D1abBDzybt8nuxLOnE0LyDFvtUd1qiBQoOkDrflZDnuFQMS0X+tgeO6TknS0lMGWpnZ6GjSwF+Vi
/jfGRt0v4zMOg0vkJyOVoJPlY04sZRIRD70npBDnxCfL/86Tr5EsQM8OWGZJm+mlKmKvfL3DAvl6
Y3x1DQ/XVWNUhu/0MfKUHGfqnn3tWLRKc9NVnXkvlyNvh/XZONQ7lQcLaF1V4/iKPFKJ31aOayps
Eq5XpfUFwNm/9lLFRp2/vf0yUh46zjxntZr87jhwWIZMJAskOV+kISwtq2nxFedCjscF+yXw44W8
ibU65UbMJjWPjN8fxZPeDXmX3NYKfdZ0d0v4Ii6ly1ikN1aDArrhYjoGMdQ92j9vjFd4ottQ1LF6
5DtQkP6wOy/dP64Q/jZS/eJWWfkh6gjLb8vWJ5FtCKfWqxNHnkmFxTCVbdi5rULyOaDk+yWqlapg
E5gTIy24SwAIwGLdxJ7qEElFCC7ww0c3xuMtPmHSHTTmIiPsbQSD8t1YAb+9YzzYUg9Fl2lodMNh
FqYkp1lVM65Rj1B9rjJyFdIdlR4XmOpSiGMHX27PsGyIfJj0dhIzDgvf/S6f8CrRnVLScM4TTvzC
xKRpSVOiQIcXDW/VpgUE2cj8g5jrZPxrGFkrTaqw1FnhtrHyewBRGFiV4k6JJ/4lwQeJANuS1UNf
E+RkvqVV3Y7B4j62Cmw4/JK6GmYABlo+VPWVfPX0Ugg42YYmanqtUTy9xRjyQZhT97dlZsK1bext
DtjgcmTIBM8tcihPeyQSdlxlN51H0+jNhYv71vyS/9l+C7z1zVyguZkQR2DaDJXQ5MNK1rYFFF5T
j0XAumR3efwaVsziP/x/YVRusivHqkarvHuuW2mbW8BOxeS9FP72gZgCm374GLE3cKAjVW9g3WrE
SsQDUvYKKe4RVPsFtDeZ68GTZDz72cgjsIOMfk//IHTg4wYfjCtFC2xaX5tNGF60mrVo7KfBOFZz
NHuk2ZaGfCKGlW8eJo7lVMqupC1zgytyWRmZS18aeiNhcD/GIUHYZzr2ve0mktUGq3AGetJFwzco
C35Cyz16l9nMsCFbjxWcoN4gZYt1ppeRR8NJpe47E+mPl5eoNm5RJ2kfqz6OhnhI1G14PUtdM+7w
MfsTcwDHWdGDJ/XmilyLUvGAHEKMvDFFMj0rMsLQXvuD47JraqRciQGSs9Ycfv09UjUJ1syqwdlR
HR4eOkRog/opSrT/Mb8EW58pQuaVQBRe9Z2XQimnXQb8N/JtOlqz23XD8oc84dVO5R+3xbaaS0sb
QKCcKLXPi9/x42EwFgOJOYG6sZytt/WPkaocwK6Q/cO9/df/u1MvInO1P38WtSagQTl9+3OmpsC8
LV4zqpqJnkGWhipWVigCFosTEy7yrld0KaqyJLYsgiek9eceRgjSj59SsmeCMZCUDnAdjWqICZ1M
oINfBqT9T3LxnpaFyWycnlXs5bVKsVsGjfnhRmQGDgD8ekI8dP1xWeoJ6mNmqNCgPdwBNmyky3JK
e+m9NFV0A5lSsOhnpFtN7tSoMvpUmSb5ymKZWakZzk8gGgiTpu6+/pcEX3DFORfIQna/FPnIfSgW
O+RNvT4CKcR0qMZCOocXNTxMu8O+sBpMmWOTj9srbAYSjB1X8ryDR/+ymTCh2E2oM1GArOHBlylG
Yv7cUJXR+1RsbBX0grujzkF2QBShLOCkNE/yJMzkx0krN1eaaRrObx/9SG8cRDQU43KCwmEW+gzS
hSpRLAPFeNldLn8Rf5h3Dn9D05P/iwP+HCzjNJyop5bf3LKxIHjyL4QOqlsUp0cNUcFqHMErHAWR
OS7/kbFyTnIADd/RyvPAVJATz28q1kAkfXTt/pzHEcwT4BwgASAlDESVGJrDNyL0Rhnpb2A5PJWb
e4lEwhpwQcFrWZVkiBRn1NgxOlxDsE+d4Nyg/rDpVNNO4RfuY9vEYFfN6kCYZFswF4ricx8lxhVO
BNLKfEV1Lf5V/WdkvrFgSQoQl8U98+NAe+n4un0VTfYQcNRRR6vsSW7+i3x71beW7Mu2N/X2ef2C
Dv0Ahb1XO7k3Hbq317/3VT3Eks+ctiFK+TuIDbboAktBPpnEWb7X9Qo527r6uqorwR5P5J/rgFce
uTc/fgg9DM/DpvhtDh5fq/GIOvoqD0jnK1aV9fPjJ1n02xYJO7HqCewbiD9HOl2+F9v9MDu8d9Q6
MxVQK/dV65X+tPIzDW/t4i8DiT+YKDtw7eVzym0NO8IFKJMqoItSzW7eSBQqNBo+P2uW0Xvm/6K0
59xnXKVakanTNRswJ4s1evXW51Gb7s9/UtabS+TXBOgHt1OLQlEDP5ahTSgB2C+c/QXiz/aGXNRD
Hdj4B3z6wAOc095NEZJZzgvqArEZiF+x+8hW1kccGFPhJRTs+cI+fJ6BRdjgY7XRoTG1TaOUFKkS
jP0gnNYFCwi7zGZFdU0DL2NhA7HHd+2XuDMNCETcJIuIf7O87gJIyzApw/pCgSdVLxzixbTp2mHf
LqKed+G47ImC7Rpr8ZyyFWFi0AuGcba2i44//FiDuNJ6UcEbwXkwGXzfwbg2ZSVnGMPbCJK7e14U
Piaxj3Rw+pqUDNjaEujYb58Ppf+JqPwv6ejhnwUbUDVBLH5ww5Vj3a7UdxxGY7krjauCAz0ZNKU5
hUQNRqI2HGT4B5Ejv3w03pdqw7NcVmeu/OZyO39BkgENPivWivjE1Pp7y8tjlx/UNthzhOiha7T/
YBnVQ4ej7qu+q8slfROO1YtNwLy1zT2lrFUdanZItJFPIFqnFeHIXrQmHrAol7OTHG3+C2nKkUgu
hIAbXoveNby04qMKaqyrphJhS//5pq03x7cB6b6tZdinkcBUKUqlF1cwfGaZq4nylstGFrKWNQ2R
8pypb0yZ3tNea0VesT2f+rUZq3qTPjMsI8LnF3xktu+n9wEJ8C0VX1O0fbD/jOBN/jtT6WZ6MQVa
5uxLEAWNqzdsInR6wmaltE3KD4Ne1J4XkNlLWlq5JQqIZOjje3VUjx0rOPfwvbKmoDVR8KhIkssS
i+ZDZMtqf2YaG+q7BKQ3ftTSvbz0ncI6IDljHyIGClOKossshx7WOidq6BiD+quORziP0NXPOC3/
+GxfthKHyxdLyD8LqD2BdQn9tcRtVkyQ4bEpaiu8crdzCki/PN0RrzPYN5n4UEp7ljhjZFl60Nki
04vF0WGq+aDsii0zl3eI+3H/0pmpe/vhYLT5XFXTJKVlY1dgrnImGIxd0nRSv879+bXC9kOUIdjq
oVLa7i09QXvO0OCL4P1uk4BnQ/cu/h988sj/VaqtzZCJ5ekqFDH1ULtadXducj+5h7vWbKoDIjV4
MRYQGrI90+Zpb0uRCK1kiQ4OYU1hGKQbGfgrly2tG51uk8JYywgm0viKRxelbeyrXkQrWKHwsLm8
QM9IXUPRUpsm2MUhU1GwB/XbXAePhRc5+W8XrlzTpPdqLablE3nqo8IPteC3qhAhUVgn9dtODl94
FvMiWi1aDd3uFkJhG77592HiKIsSGpD7oRS/IscrPC5A/UYa+MdLmipCxVE5y3I0s8whGcaMCH+x
v2WrohfEr58R0N97CujT8+AiIap+Y6pXcnE2Lyi09sH4Xw2di4XzxNAYI9zUjJKD+RoJi7wV6dUf
tGgAoyPk8ONpPBU8/dn/ukkc60ToLLK8Ww1RPSDXN2UXvHPnsRfGFidN8j61wdJcfvzYI5S23+qk
U1P9ERRClQeU5uF3k2xwMLXNbFbsBXKm8SmhIhWxV/cgOI7eT7iJHWZxUhqYRcJkpMIVKVmRwW1O
dCaeUrUf8k6NVGFnWbFxlsi0APBUu5lDFfWGIivFD59e/QXAh/BCIEvkZA6wtsEtW6HkhwVDWzkt
BOMG95AMu0YPFT/eILhxDb9B8P3OEXWtQgFF2mNDX5B/6p+B49GmSp/rAEBQjMIe2KZv1kAO3u2n
n+wYjo85Cafm4tHmPrns4c0JlWLoeUm4Z0+GvYDyD2scxzzGQfrsg03+9GJ/DtqX5dBglfEmWXo9
Djg9VUCBOSvFQ9q8XXRgogaeVPosEmTfubNTxFVTNKy8XX2q9+6JgKlH2XQEAwEnOZqvwlMIi2/4
5yaoQYFw7lkg4TPcyZX6cshrGLVbiT7eyNyVrI7QdOp4QKoyNxBfN2yhmt0m0hppje/5oPxSD+zC
ul6Jpdb4KilPIBtAOW6mxL0xz1t4Zryi/7aSOUawdhue9cXBqSifu7AsffN/YPKm0NP11kWi66SX
5NuOgrd60qWlGlj6/HiNZPeKXovDJCa8bD6NHorJawOj48+FuItQHA7Oyd9X9LA0+jYowuHsZAce
p6bQ+SWyR7/ac7HmWZ4vV/TSh3C9KLZOlnqX4NeBANN0kWoCrqRZ7qcptFDzCeT4ZrdKl3QoybwD
JU0sNF6T4xh+Mj7wj+KjoNTsNaYLC2Ffh9yyntUU524Mnh6nJJHPSTJm0K0LotTlj9RCnh9Wy7WX
KIwR8TEMiWEn0KA4x55BtzV8oXDfFGloubfj4uLEnwLg5keX0ohl6bpMVOOiF5mbROiayVCsRmn0
zHARFbscm3ZbOlx46Oochn9guWadFnBONJQBB9yG5P3rtGVjWeVs3jF7wtp9rDMDlcAYy+NHuiUg
45w/JK8Ukjq9y79AGD4abTR9g68n3sDs3fbN7GOAW0X0/CrqT1K+5TotJe12VP07oQxYejj85sEN
zT9DMxq41HY47pKfZ/u6iizMXHnYa1ZHyYDPKLe6ickpgAYlv9NsSR8yL7/F+SGYQg5u1btA3Nr3
xNVK8Z8D+InFFJBg3lEpSGS7nmYgDfU6SFOR2WGPUvqqA3+0u2yMs5qqvOkIZgd8WQlulk8+6SYA
HdWhshKkuePBW0IhHXK39VF5Z5eqGWHRIUH2SGrDg7cSYfq9aVUHI5JhlEjGY/mz25KLOn06Fboq
QhguNfgZSp3mmXILT+A2xoWcTIo+6G9CCb6yjO/JSPqgew8zLCFEKmpA1w2cn+RTKIvBR9mxXwGh
42vsVChPMXD+eMhAjmDKiAyahnffYlEt6Sp6xDhmBtWjS1fnkiobZkCtPkhRvoZahSDCbBDPftMy
vlZWdPmGKeHQElSxvm5ja7A2SuckBozx4WL4Oqiub3fCaKqk+UCLjP+9Sy805B7rGlepEIRgy6q8
l/SUSUhJaer6vCBGLvVYOQAPID++Wt2sP6wPzXa8gQ1bBSZn4WCrJGvdIfdnROdLJ09KcEA1ziMz
Oe22zl45py7SI0N/F3pSrTsZaowytBYym/ygwRuLFIh6hYiQYi9ISzAK9cGcUl4Xqn3GH6iB2fpl
L8qawSr9KBlXf96R4IeW9YYv6IIXTQOM9zFAsLqOQFZ7rCDBjp0IIjHYIxJkcHTG54t24y9bM9S6
GT4E1HTVJtLqS3GC1MImo+VKNk0eYfnNtmA6I0VEnbZz/pYbnDybT0fxbj8oSrvzdQXJtEtmyfQA
9gVneMqKC5LXSban7ydYZX8B9TNX2IbA+yJ2d18i8/TuRrMbRAMCXjyUW2gw7ZiYPpsG4mXBbi1V
85VUj2IVArnWOfcOmrCfhIuRtH/PAMZGBeg2diSubc82LVY1pubYmrq7SHZh1eqfIpBdA61BxvpF
1357PjUSJwKzc3XAJgK0+KpzD3gqqWu1f8JmmDiKuiXqlXLSdgRyoJIBhtsiqmp5G/jmlruZkUah
mzGBHc2zqxEKX4G3NXNPVJ79fTrxCSXs75oTnOFdroH5Co4qNm6ZeuVcn1Gw7H6qc/4quzVT4fai
PSsgSQwEoMO9tiYlHYZUHWAbJ+aM8KvCnDrv+x4SAwG3meUpQx0uij7OpButMKQuFdrR33kKv2wf
QH7sqGXLfsY0YfdNmQb+A+fqVZTDK+O19r2TOroLWQfLXNZlmoJLCKW+M2hJXHQlAru8JybJMCk+
HdpnmIDAmgLIJBsiii7TI4SU+OQ1b6LCYh2MG5uL72FCCPRGdhS97MXVS7t23rJ4A91lL+QEab/D
8OK/mbtcqwe23TDOUETSNj+JbM7CM1BHCORwwRuXKiywzhD+iBm1x8OQIfReWsZtcXjQ6BAjMYyd
42juAyHqVkpX4bLA5JRCI0pmKkajN/a5MNlahpfWcc6lGNsYMQtJT7/UCvSccpE/JZQFZrydZSWQ
PXyyeAMKFat+gdMcR7phXIoTzajIsAEe5KeQUulBJC4116Z23Tt5P7afojlz7nbePUa6lsmIz/Ls
lKientUTB3Q4WinYzUAvU1V7pb6ERqUbugdcSjO8PL/9eG7tAa2zGCzsqnM8Jloq7H6hVV3GzrCJ
vzXPn6xGy77nfGsQ4MkimfLOeM8+9Z4QSTIxMsIx8wZ0qdjBhaIPl4Lqb6T0MJh2AGR0wB848DdG
WQ5wcDxZ6VzGRu9RNutY506vuGmsylOBmAR03OZ5y/h41fV75464jRkBEYRMRxxppjt/MjP1C+95
q3F76qOfNDzWrd84Up0r2nKC8dcNczRF18YV63I2ggOC0h1jea1z4sx7HR3FaPcyxlM6xWE+dIxC
hEDiT+i/7eDscX8F77HfC28hAdhuVfAoGKh1bQbC8wCiQ/9YVQA81zx7ZqGyzEKvHtK+BQ3QZL5v
bBo7CwFQJ0lCIilUt0rxOzHhXX9WyJlcNsEbTwRFXRa9gM06RArpBHf0vemBKhgGG3GAzGSpkFtZ
VKOqtpp78r+lxKBjopl7aLuxCIo3xbWsQzyiAKc9V8KEfCzvyicwXwRoC4WybMaqWK+qz3sk4jDY
Uo53yyV3ewU0fck7GUKZo4iNJRq0V4x1gB7+FH2ARRZQD5oadr4KoikmW1kVW43I0+gxmjCaLJGn
oMnaMDr1DSDX4lVsaSwsbHgWtJNpFnO/vjFHlELI5GzyYA5Y4dBQzSsbggo+7BnsbEbLbA+FPBs1
hU61FXAH+wMY3TX/KgonmCXvgODUtl4y4oY34irci6lq7NEJduhf6PkwiwuOuavEUp4wP0UnbxqP
DEvEi31hod/y1WsXi+GoBJXoGmqwpXjOjayBAs5/VRw4rx6GIf26VOSqrxrRbMxb1acaKXqbrOG2
7K0eH3bShzTTWubfhEgUh+NqBSWRfTY2F78r+gC2mtqEFNCT/W7Cxipk3GHWyvSAhopROag2pf/A
E6ReleWnB2/hl8FVc3ULRV2Nl0KoM8eIlI1yEC3WdOEHyZXpD0bahw707/1OvMT/YlJZ94pH9oF7
vPE3JwKONToDa0+g0Z3AM3ewDgSC5/xbr9bMbezv2WSZUdPoOGukIa9bTUp9IOxOZko5xjXhRS0l
trVZpLlVD/h17Cjb8bCm/rE+9Kemu8Ynxb5VigiX3sPCPbfc3VYAmHCGNwV0GxLAf/7t/Z7I9Kri
on2KMig7I48yl386kZtjYqzFjA3gB1LQPG2J9zn2gIJ+wUK0Jsi+cOJnTzARNTqRPN7MuUW3naEA
o/9Qc9II5OOPb3eQK41sXaJDly92kyTCU4cbEtsjZaZjuj5CgP5FR++QwWhroc8d0jsOpGmM5Bg6
EG/GQ/jM38FM+5Jf9PEfThTQ5tOfKMsAbE2OULWElF7FwrEq9CC88GFk182zkUsm1O0S3ud+F3x8
DPEfiNx8IfTjy62J12T6VdlXLgPVQ1UOEr+0Is/h9vJhhs+JXqlgd4p7gk+vsB0CWPduHykgqYIy
NXo70lpd3j7h4tMXmpfHbCKtGa3zE2oCPCqnfJMWr0WbEHynJsRcrMJA4is+mJCylicCij7kAO9A
IhgC1wlGDDgp3VYsEIV2FdY8Ws6sDr5REqjlb80XhH67kjicILrajp5NTnTEEy0DG8movloKMKJV
IzKSrPJ9T4IwgeLtNwGAgjq9rQiJwRs4EWbbCXj4pRJ5jFcYZ0f89KxxpHNTqrrDc4xx9A55tnDS
/rTcDtYlhoe6l4rIqc/zqgpBKPq3zi3ctX8f3KRShnSvxDwAQ8kVJeTtxTDOwuD63Ro2iZ3ToH7y
CmifbDpkRwXyZUXNqKDzlxnxHpEZjHmsK7s/egVn4qC5/MPlG9rO1QcWFf1+VTZFzQVZgXXXHhYL
0eKQEiXiEWRigh1zMYT17af1BhHPvLjDddYy34x7LJ3cPcY7LKhryLzaIBQbtDc2J4kaKScMJN0h
b0uzaryXKYodc1IYEaVH/Lp3/ppiRd6R4y5qiJz3xzCIFjm3xq9LfdDbv3WoQY5NOaZIseSp30K0
le6qQfqYIFoAnQJkuVWpy9JjnElQPjzYuJtX46q50+8YmV+a8tPD2LpiQDUlVB/Sj5Kh5suy7MJF
d7SVWKwWlFV/rRvX5PqxJVOvw6CN5uH1BvBEEjUU9OEQtgH25tOQ4uryfRXRqgkEhGQsoZLlycD+
okshRepvaIISV42tPL/FHz/yunPvcRxAvZ9/a4IQ+eMPaJH3qD0kIvInSj1MohQNS7oWVi/CTXCa
zm//6aJdQt78dOsjgGuNcSRIRgsLrJ9QsuKkfU3bdjXsMwLetCrEVcJ3VZApTFucY2Ek3k8XOIYo
Y9Smm9DqhH/IH/+OvryQG0aC1FBmPdFK1ULpNjxK8GmDFAjK6YRdpx5vC4nvGumleifMzaUp70Ee
wrOclbHokxcljZ209GcndIS1F2FpqTJzVozYsxpTDt8LnIE5cfkYzC86nVilNhawy0v8YThrJGBh
SQJTr4sYxuKTATJzTGQelNzJLxs6oKfamunwRC/vB4LKUVwu2QsGNVXM1DQgg5rLz/QJ1F2/ed3c
d+DJ6TW8kle3bHH9fjopCO6PolLU2yhh2PQ/IHKTmOLM4x9qgq4BQiadnZxcB8rPd/wIJlk5ie01
emtFcaJ/0YqwTWa4pBHVtfGi69R2/9TEsG/LymiEH28sNnET9o924tpD85sFUZhP3E8XA6KTYtWb
ICvO+vtPP+zEd7Pspy5kk/BEXNrCanBhVFGeFg4UFHJsBgeA2AZ+kgt7p4HrbcIqipKc18fQ83ir
Kk7SnazRzoSPn6Rvd9IDcx42XZ9/+WyUjPippRq55jszkF0heElAa1eWd2UdCQoW+jnMNXm2WxfI
ZKhMuE30ajftn8vFtkpMn+CkAzPv7AIfvHIiZtdOET/qkeP72f8bjIJO+JwkprQ92GfVG09ZnosA
oqkc8Td4xGj6bjQJzyi+fP9iUgW333erFiJvf2PPpsNz89oQiVVc88M8yjfH6zZO6cpuLc/aG8eF
EhFMvKtr7KB0DtmjL9ouiExhr+vRQXvXngZp82SPfnULcaZRA0LSO/oKJnxrsrv66/2Gc4hdymZH
Qjg/P22uS8J/iPz6W2FXaNZdLWXQ4CVJDjxExeVVQOk9MnY7n9a7Tz+IVIE4FNWsc2TesmTSrpHU
ufPqEX8xVdBxYO/cDT5XGMJteFxErUw7iDwmvVMJ90M/JlHoEyYkNK+N0tCFUOzhBZk/hPIN6Qfo
OGzdICQEjL/wUQokNHMtHaXSsLYb1fJ7MOk9DdzDuA4VbVrF0Yyo3phsIgfost5YCILLedxrKE/O
nhIBwXJ0x3SWcmiZJZitHfQy8WqyKFRYV9oMJG4QVxV9oKNE+ctQMHDjIX33TH/iArxZFT5NDbW0
k//pbDaWE9cp6zk7o644G++1CQui387nDX4sQvLC2WzHSU10s4c5snEwGui+bzoRBesPgelKY/uD
A9Fb4tLSMV7ZcfS4l9H2w5m7cMxN5Zz6+p7Zt67HBvWpmjAyAYuactyCdhLp2LVKrLv/GD0aRJEM
kLZpUykMbffgPqojGbfhdHDvC9U27UcMxkEt4T087ix+hpHtBWSHWcBckGmLdkUPH/mP+mrX/6Ok
xgWqKpCZp0P5VsjyitsOdjdYmtYt8j1111mC5U77OWa4JvCvrxPA7D0LuUulgU0RwmrgftSGgl14
1lThCGYshrm5BFo3AdpYbl234BlRiUePL/tPFqRacxY6tK5Y5piUYX6J3WonEED8xx9bKmDrXoE6
CPAgqhtJK9ktV9xFqvBH7OuasSIU7TtLUKhlOdJ6KieMHojQb4nEaGn0CPUmFlO8hwvRE90kuAcg
6ISbkqJAMTe+hxb+TDbwx88yhkb9IMxFLFlFpXOyzy3t4E7+MFFf38qgmaciKrh6rbCHPQzzJuKE
mQ6Og0JTbYYuFdq7BiFwF6pUKJ0EgmsYkGw7win6+gimrK01uL8Rz1wA7/ZDge2Rf58B7QAOOtgp
pVXgEyc7ztbNOzg/y7/89CzRmHfYoZRn9Nkwa+RwfMwrv/YZrUwegz66aaKUIaSgfzVmEViubKad
t8fWmtgKrihZUYAP1w3UvVS5+jBhzR1FmDDAyS0CmaOkKSyzQnh0rx7Hu9ygzyfhnP/Me8dh9QUW
LBQgIdmqIKx57xmxGz9bbQRmXL6vhd69mnG0ggMEWkT8BEfWMyNvm585P9Rv3J4ZeqOUNAS3f49V
uBtbv/Q0whGzn1zEL8ThPbUun3qHSyWTn8BZhjtO/yvYM9ghkLV+ZSx7lYu13CTSeBeu9ImzaN8Y
FFy+Ub8N+S7Jooa1U527KkBq4gGBU1VBavmmILeedo0wWI58CsKNP5rJXhvu7jMtor1Hd7kIgy2p
jp/43xOFjKJ6Xs98a/PBP/42ozFb3ky2HCxPWerh/WEsRkErE1w0GZzY8wTVBApM6H98V8ClQxqt
CePOAuO8CKh9Rdzb8iieAt8cmBwdvI+I09zIP7j+yvJ2RSYJG5+v9hMCFef8B5vy6+ZoYJYvEJzh
QnhYox/8FeSCaT/N4KdoeOdQIc3THaktA3HbVklmGWhFWTPjGRybAlPVE8haTUQNb3sOSPLG1BC7
AxLAApuuWrB7iFQdjbCpENb8ISzqNLI+EVEUgSgRz0b6fCOfGUR1nBfpWK1L6B/1mM5n6GUZpcfm
8TWhQy49OAyxqrk2Kvidw6uQelTiWcNC6uhuznCppUib1FyHxlC2bzahAPppGtMYme8NDLWn2+cz
vBGU3Fr946z1qVltjR4vBd/aCCWzHFsuzepavvx9paqDBKjl3+DtzYbxu9GqgzF1MCUBA2ZHL1x4
QPN5z7ztvwJemKeqhGFyLg6aX4Yt+wiYU/un7xeHo8Q0z1gSMBYiUDlEScL5n/dfvySscaFbz4Hd
LvmeGGtEd7lHyqZGEL6uuiVN9/uT6Dr0OfzHnAEvCkWVWuFv8yypLydGOCgGBT2pWD+7L8n/QJnr
JqDCSiUf4cK0vZXiOURsyqrXVT7i6rt6loiikNn/zVgqJSTUYqsIYDglRAHGowRkHuoWQhTWYTlV
LhQtnWYXD4Qge+wL+yyQrzNv4fn04t6BTRUxZOXqw9B5KhrXXQJEQBhCC232mWqXGRyAtoZqkCqF
dq09u3haHBmgJ1ss7Fr2vSUqilY/9pG+4/f0FJjV4B2OD7UfrRxQ/01UtqsmAv1LhlXJ80jD5YZ+
UwI7WadHaW21vLuwXuYs38TtFVS6tOYikjMk11gFD52lE4oJhTCCu4y5vTZPZnSNyJPGKSv60E2q
13psaWpXmrXnpyY7+sKom7nCAC8B1ifB9LLrRNE/Asl1/GJbnk8rTTbyaIDrdIW1towUDr1Lz95O
oDE8+q7DSu/VcDYhvkr3joooIgck2U7lrnosUuzQ01HkI6rRrhABk+kQBuio/1u/tGoyQo1iaj0J
M/f1D50vTG99rTxbg5hQlcfJLj1MtpXSKMQZUdsHowoJDsupDChLt6ikeF0ptADijNrG5S6UC/Jy
WtrofsjWWc1+RN/P/50BBzBkwbZRTFPDBLOjQodSn2wukTF3P3nvwP2kCCcv45ccuc9cq51IIQuf
bk31lhICNP8v60we3i92mCEZUDxAPco4hdwPQrDwyWAQmmOHGkBdbO+tSnUOSl4JqEFQXoEVqnj3
99ePWMCsm+t1crWnccc2kP3Qsgvk+W/hJGWiz1rDD0bjleb2L9N73TSLwsFnRonB9nhb9gwldADH
heMVhm/5bspRvajfwUbOq6YRM5/DaEGZhqn/lYR1PlhfaIXQrNoht1MlSHMgtyyKfEKjea3VHtxq
RM3InaDc/RElFVXiNMmpODx/W5DREV3Fn+DXFde1F+cVJiqUx/1hVdVdc6jswP45nAbqGRmCDvId
axwKnTC6sGV4Wcy9MU4foMRwDKOSncpyStuax8FBlmlrBF8kz6Hl03Nw5j7QB70BBSQgSGR+SCIZ
nX3rX/jaVJ4PsvoRdaZSXjIftTT08HVymzPqQck363wsrQ7Ntqa7UB9Ip35NecK3Pd8oKnqt5oz0
wcZhuOHL5E1ZDwxVSMRYK6WbyADRBBz8K3Y7QsmbZM3guLRnLLCVOZwJ7qbOYnIqCBBV9JQHKfiH
3f/gha+tH+TTPLpIw2P0yepedUz5GUO/6F+qS7MCwgTxbckOjFhG2HgFJWD3ZvVf01DOleIguyWm
Ri+aZFpCnr3ZERKYcgTTkmOGESb2tY9MrCYc++HCyuAZadN03PxC8wg8LwXOBOtzccW0wIGyic6T
D4FosCciwUsz7nkCSh49+mlKTsK4F1s7LgJ2nqVP2mcrOHIreo297Pd9A49UrkyEbS7zzNHYm6pm
BfFNj0Y9avPVIrr+AhntZVazd3VB0/J/+7Z4/k40vQOC9TqY9bq3c0SG+JXBfR6uim5M69GK3S7O
eIg1quWYiU+H5MB6Qedsif+jajMf1r61x8+Tt1HvqoR4E9cDZ7zlptpAtmqwEpj12qZcaj1uwlvc
RHC0C5128S1qj1AxeU1qFOkmfzpq1bsjaYcf2QWFPYUyJ4fouTquD74xUQyffJWU3KGRYFcsDcpx
7l83V1oH40DOuXoadO4at3cIcK9W1FBMW/IvuY1UmtesyE9d3QwR0clFp2DTWU6SIcGSWfW1RjrF
glEJdJCaLg29GE5vFNAAHpAKavDD58v6/0rTUCvv4NzaUwzn9VitvmStNYbG1DJpsq+mqU+ojfOu
Vge2653ZXLc6DNNrGMoNz0l0Y2n9jWiEEQrJVLW8cq4y7hFEp0BN+SEyYqsm0jXdIKJZ7kV+yWuL
OX1ZHuT070pdwaFeKgwv582pb7NiJEDzA6O3C4mF6Qfs3BndKY8SW5aEDaEpWwel99OnxZIPZrmS
tm4uKQDCv+v4F8VxP0GdI6XW7yZcjrhnjmm8lHr1ikyF03JtvoxnM8wTIAos/mrg8B7mgzm5zO5U
MyzVtAZ0bLTOQnvKi+h3OxWLa7CtcCbeNbBhYEsWN0ZE54ycns5kINfyUOrZQOKYlCMTJXhp6C+d
c5T/BQYxCLPUsFYT096+Aj7WlN7o+itzT6DWFAxq7WpMP8Awsl39PmCYat5XKiKnlh0Bu8ljgDDg
keGO+/YFpbQC78R5WRPLi5JO74B9PU0cEHi53j01kdRK1PCqZaT//A1wIZBSg3ENzRI0E4lhGb/4
nJLiPIHrablAl4Kru9epwjf7wkKVD91dyhdX0Iq19endcO2F0dvAJFfDg2h+l/qpvIJlbu+Us0pg
kc18nlkzRpFqfwTyXRKZIAW0VBB5yDy0T39g09lLQ8d312PWFrNyF51/eRRajXeiR23HSy+bhbZ4
H8qbxMAlvHWaJ1WPrGKoPTqDcvqCEtcP103P490Ed8S81iTWMOGrAfjhUwkkuyYccKlufcc2Y6LV
a/nU1b3KTsCOfMw4RHL1NLbHqTWGcwus6THw8cewpy13UDHqx4pMCvZKuD/FOT3h2TlE+L3ypF+w
JFn0LQ3OlH+m5l2nDSAYdE6veANxrYVI4TLXV/1WcfyMbONU7ufZIRsdoqBAxSjv7RUs3oJHawB4
6aAEzS4JysGs/2347rhJw9wvKCHHmuQconTZh08NS+OvLe2/nHkJ51cGVkyQAbJDp6a1XiC8ZpOy
oXZcevB+pMSGe4vMRn4t0tiU7SASnROi7rzo7V2k4UbJTIqBfmHa9W91Ldkh6v3LQdr9NFbcBKVa
09TRI92+KU1hF0EKezA6D+TYbim7e5APl+05htk6i+vowybgFyA4+J0Fx5Wi33JOcP4oJ8MV7hmh
wGLN6b2HLh2LB8bS1AIah45rjRro/L7yivYAfD8uIbshSzQcmZXiyMBdcXVrW1WOTre9tTqFeLOx
MkGsULsqgCbpI9TQuT7BFMtOQRWx48bWMIE0hv5d+rjFRVJFkIPgtzLB8zPaztI42Ta1veog8y1U
Gt1G/22wK4e1GpV09zlU/kjMakzfIv+09UmeDHDmbXzrs7VBd4VV8FBhyhUWJ+wdGzd9Mwbc2wmX
3Y8CqE4IH/ymBZs3nYPpwT20C32OJ6REWHcOWq2nkCfFH8jzoGdTz6SC/VcbxpU35uef8lyaBFVK
9xCqoC3MNgDRU5bdNqdIGE8oc7vTuRB7vLx6wBKlUa0So/1kLvekrS4Z5cmvLEBtxp1GHKczG5lm
pGgW/WmtVE+K9kOI8pAeDQSbVHrJpfRmII9Dn8mUgJFegpzDHQtczhsnXBywEcsZBl0LycQrbMaL
1eCaHUOTcQthxjTsPRdQkvN2OBl7GeO3GzMouaJKx+axKgLmrfeHcA1g6YKUC+0i4NQLmZzAKIAf
r8MEWDYEPTpHvSSp5heP9+Z63/5DgT74wGrWHj+rfhKpIAjgteO7fXbNrFg9/2e0zCtT1DB8aCsj
0MH0NdZjoHpBxS7kYIye6W+AoqgG5fLuRW9IQVUfHwNIuJLofk+MXciZrHmxF3MbCL831h3BFX30
TTupjdAmuzyXUzOBq+KrkLaeusPEU7P7nHPg7y+Mw/CQqNUiKycN7YyBgvi9YInS6GbqhBtjdu3/
J4pBXj8QKsfO6vyNGRmWAEZY9fZHdqftfafJxvjyJrHCufuKjgNXuchKbjJjKMrUnQ96MKmLjxi/
oDhkfe7rhhGu3j23hnHXBeg1IWYEAM2ANIIbwQGFrvZ+SsnRxKH45kimZ/ySuODb+JqLaWXCU/9M
gWc0GhZ2JkCoAPPbse+MIpxL6W6ILgAhG39b1wwpDy2pIrSpMo2YSuRftl/K3m+5wVeiXW356zCf
Ln+3DRzhas9/6DWBqbgg7MEBRw0RMMpGKKiFfIqeAP20gYxfTm7t/qZV02ev3D4iLh/jNl8WTubN
ULGGZqC4EmeMct8wnnP8OBIQRzF8U46qQgy3hIHK64PoR6nxBaFvGDr7DHPF++9SkM4XOte9PchX
A+ewe5DOIU85eG6qflZMwLrLUgrztko7zDcCsfRi80fTIcgKHVi2FjeGBEpZpvf7b4pTjGcQ/oPl
v2jVlTUsn2hjNOmgFrhOFsXErnt/PJxo1dx6Tbq9r++Wx/HUKfuTle07b2PiBDqyyEg1/ZBVqyCC
Iq2sThm5pZ1juGUOSqdgGjYiq53YhbIEid/LvOqK4zCGoKvjQHvJimdxQXoSkLCeGRDqBU3UHqIl
h6Rsfx1EeFWDc8gONDkIPT/+BQKhR3Mvt8PXYMxoVSwbpys0+kJPjSlJyciSXpK2X9PhizaoNKgu
gdmnjDsqQwZWQxY8TMFGxj1pSPazEHZZFRNmxhVjaTy5xVA8xZCdEKWX/RjAcqQYnD6GCrT5gs6l
3we33ZPUVHAJLzFL6hMiqbnuvXR9hSCOSzh/91lxzmwDKbozu/jzvnJI8nHfqilqt+BUlQGLs8iX
SH7164xufHmCfyxN9qUW/fekVxz2GUIRjwf9bzZfgQ7bF+dfOGXZ8u4r/d7B5jTq0d8Wz2YCREHL
hNhJnBlWgsmh8QWfnHiZgOPmyHbdi/KRnlbl+yW4dzNP8+mlxm70WuSpgTyfnnKvWOeQlF6CJ6iz
AOxkPBY/Hqk3UrNreS7qfhkIxcE1w0TGg0bVMWX8ogzZeZ/KLedZipLDeKQ4arABRZ2GjCMaswFr
GxQl5miUwombPP/saO/8Q4MesxuthTA29GdSstEcaMLYSfaCMy+eBr55NxcvEZZO1CeIGJ1oRF21
uMD2AEUMNxLO952hwaPXwGpkKjDgNY6ZBbvvr+XKp0adD5zcVvOdnD22JYG86bPyNX9y0GDJ6A5n
ib2XG0tMHaTm6xDq40ZA+7RzFUF7aStQvQgNWbKHs3h1vIRR+LFmLUFGnRrYXFqwFWcdSKK1A577
rBT9eb++o1TdVfBucNcpUsTFk8i0dptDw8mUDYHNJIiuf5wceFcyQf5GFtLKvpS2DK35EahsabhE
hc0/qa140BYeofejxoA86Z52LUocUhkMpt8OH34/8HFjubhbYlFoHlDkOdyw3fK+kr71Fud7Uk3m
N6+tIYFHAehJcGgN2GtWDWhdcr8eTqcrNzzL0qFEBPOQW67qYt0qv5KVqfl7SLDEdkx9sdVZundI
neltAhhdUlTzHyQmkWqQ0A069WBuO9VLhIYpvswvtSvbeS+4C2f07mGnthSLT0DpldqAlo7rUH8W
mjKqfwiX3OBGCqtzz4grF9Pdn1kt3OG7+2cqcy4amx5EWvt6BYjGNKq31hRIPfGe2QHdOSM+wdep
hjyF/poCgXkIq5UPsu0XrLMIWqkv9NXj3Gkf1/Wdz+ceiJuwVsMIDM3hMCtMVKjs+vusuXoKHBrP
HaZw4+2AF2RTX3O1Ka9KuiDoyuE1vcdxP8qFD9vzeXsq4udhWfadqIBjRCqmv8Luy9EaF3ZYvel2
+ZOqxk5CMYgK9KhpZu3NujgENImTELVCURARgLJYuKdY9vvjbyp+46vtmZHRpqOOHg/6m/2CXveF
cpnRhjT5H/nkoEcSS6xblS5J9kP1SUhVAfvW6dqocQUCWSI+l+phlIKs1YmzicdM8ahOaMlfJDQ1
UKN80KGalk/fLKJu3ufIQCSzoobkFmQLi/PNhzrxs4BieAC7wv8rJaGjFULI7aPF6GS1IORLs4Nn
EILNkB+QpR0PT0GQVYXYXaJwryAlbH0V4p1o9J2z2nTHmlHcBRo65f5snw88yn5MwF2d9JLogs1Z
pvhvwj2H3OknAWJDVP4nxs6ad7/Ry5TkN9wDO5LPrsU+dDzWOvCH5Zwn6Wn3Jv8aI8Ts2x/B1uHJ
UK0u/vBX5gxQZZQSQvXH4JOuEiC4F5trUGu6RoiFe+T+aBjrclJGmLSjJHMXb1xTKkJEvI7zyAG7
qUrv+1s/fIoILVMbuM3k+Pc5z5kw71n3IdO2m2xcaTVpEljCBLQWqv9UY6cszpuxyBIog9uQArkB
Y1GMsAvKhUnncMTMRbL8Y2qrrqTMzK10cnvERWnHRd9+TdWMn+L6YzPV3nEX8xeDlTZqo/nQTszW
haTzbgBRKrcWFMyu6Nf9fwk6wRL0Tl4L/w6k34r7ud+XAkmJZ3FJq02vUeuCB/Yf/9gEqYHjmUSA
NQjTsLjAeutPoD59/O1kCuIKSTgn+1Eez+chGRemBoDLs33QRSn0p/DRYAA+nlQSjvzjYjfyohix
PfkbyYzt9UznztUleMxvz26EtV8T+kXId6Kbkus6HyOyAU2IzP+88xFq4x5bWmfjY+qvNd1oEIAp
puynRs5U3Y8ly1M42OKRB4Y12f2sxOwacXo2WKkjVCT/YximyJGvs8gmu1KVf8lu2p3anfwf3V2T
5nLDq4pz3CpTZYskE9Mj07ERdknEboC8UGDZPFFulLrKTV/QeGbAJuYfdd+LD63ntspwzxgozMLd
ZpaENexrJ1nlKsLX8l+ABv4b2CbpFIOHDWLP1CBYJDfp4XwGnpATvW1m1LIpXAy0zl4aOEmcK2Z1
NGBcxLvjVtN7qTX9WRtWnlhYIA4B9LhApD3hpspBWU8m6Uk85it1iGkD97b3LkMa1jSN4n5c6RCf
nuA0isnC21ylDiUh+mjbUfmoLJcX0/AtlCBlCGmXvQ8ohG+Ee9FG5lleTTxo6A018PBP9UN2Phyw
umHmnx+kggsZj3i0tQunczYaWdsarbbV3IZumQYvgj6GtTL/atYp7J4jNfbcLNFWM2GHeUR49mKU
tbfE7hRC7HxMlg3hH9okwZYfvgSzYcCULAnDdhHLdu9ZdDjwF+fUq7N2pO7MYmTJVHnQ5xdyydqk
uV4IOby8A9GrEiXJp16g1GaaklTb2A33IdeXlq3ZO5xb9NyFR5Zr1w1lsjfN7c4zZC7bdbOI/WkQ
S6MPnfG41WD/y7r2NfonoTHhA08i321A3cY35czIsZTizN0gQPBGgvaB5MIbQz6I67Om/MC3V+IS
1GtXBnArcaFnGZHbv7nH2h1aMGJTwKkSaA6GVbqvyduvlDnQJVXc3fzc1MUW6IsTbu0I1MWFKajR
Eg2SbRH1H+yxljQlgnP+pSo4p6GdnqC2Og4bNz62UnneJZ9A0B5iQLl6ISVllg2SKppL1ZchHVkM
6FGahbFvX34fsxHYZYbiU3DTIdSDGVGfODC7jTP5A2bu2VxWEkpIQ3x6EFnvgIHeWn7PXgdF8t0U
XR9hZg6cEz3VGbxnIYMtteRKuUcNC3fKlbpfsjuyOYHhwbxU05mq4rA76Jprx3p5i4DYZes5C9cP
3WTXRAFaTTgT/0t7NzUatPTqObBMGOHulU3u3HXyU1IUoWJzcXb2YjeN/Y4Q+7ffLqaLunx/EmMo
kiySN2yT/CNkgup1htidLjcXNLQ6UWgdU6Mgbvo8qEP8/83phMBanIsTFiFIfWuJuC/txS75zLM6
cUl9pYZ/BLhIyUSl/lHZ7YADvfLL0vU2aU5H6KQ76FS+vqKfDZIyBdDJjXrQF+hpLABEP7JJNLLy
9jA/BdaA3kWGMJpvyVMwzhAuXPY/uEfeJOc2TNtIJC9JCXhV57Np+8hG1i60vkvKJ+aVBJZtrOpB
4SLJzjCXjRUkzFy9kO35mArN/7rQU4ZU2KNce/odipUMMxQsGnmhRt9xRaqnjq04H/uyofhBuse+
2Dvydn6qlvCp2umpKKg1+bN7rbC3igiGxFNnIegpJcQHNVdVPKD7eCz7c2GIpAQk7svso1iDz9GA
7yv+D72J99cFQVryYw9OAtKAJ1YNI0JBl+5UfdBBNNQdidjN8eU8PGjDI0hyTUuoxijj2yP7egom
DVyOjUhvPzLKWSm1Bb+fbZPT2icSiYU8B/gKacaoVev84bMEd7EEje8meF60EjPhs7/Uemm8PWw0
6gT1+Cj46HHHYjmggjIb4W1q+2YSfda6pIVDc+vgngcazbLm+LNIDhPBb4t+r3V0BmlclJGA+GMD
vhrKn6RMprOX6rLsVKAyUASleUW3AaSwUzB3iVJ9KHdkRn7QCqgfg/9e0Jf2vfobpm3P+bYX8wuz
Hrdcx+h9GlgLOvFJ7tIsG08xF6D3KSYDtk3qcX7wb7E2TD1EehXlo6uS07LX/QCXuBcgIk4290Z3
8xnvpi1hdPjfocO/JvdghQY1h36iQgIQ9MXY9EmM7LxdVa1lonWrexybipklVBa+bqHKNvv314+s
6yRLbDk0oYcy452yj5OOPBTxlu0yK8pk8VOz+xhzal1F8eA5AO3GbnCIhJM1YwA5i4CTLv4t0c2d
Iaw3wL+nniRNQdZWo3JWe07UufQ9CSWeaopsw+blFG3Y6EMCsxggQWppByu3jFpurN2Iqi2pLEw2
W0b3bZs+WBmJ6s4G7RWYnTijfbEzYBd5DyrsODesazLiuS8FyCbT6m1bwfSc8x0l8lNqnsPmfKGt
H/i91b6W9gkPI+wsyUEBXKu58ywp/nq0HU5TiuzQklvCeZX19ZpQJ2GcrbLwfSu3TuaGgIqIagG6
XJPKxPd71OYEWaFNZ6fdqNDD0roQlnC0GezYb+mcOZY9dXA/fguIHDvcNy+WZlPm+VCqIPETG0Sk
JPxIT6XMn26z6IouRGe4mgI3gsPMlpDQCw92hQkxhYw1mg5YhILXYn2fPRVxN6BzaUPhbLQ+TqJ2
qR6q+KWpiLLXb3ocxMabYFRCNj4DxP2f78VjyvTQpsjULX6v3Dl7v0HJ+NB0UWcVFIwX3X1XVf52
Rg+XzNTa3GFAakXMp4Rdvx1CcOwMDwWa2nWXrTDkPqSwcdRG7osHypetDfT2skVXoYxsfBjikQd5
PvYe3vaHxtVgZQIMw2XuPZl0OWDS2NGbLxbFCIYtMp6hzifIZo99AE1JuErPnVxQ0cXzAd5l7lIl
Q5nbeVchejdr2ffpLqDpl/bHm2wELAdGZX4Lwd2gOf9BggXdb4zk3tBzORRb8eslly0udveukalM
RAd4YQDKEybXBME1zrfA3G1KAR0/Y+WBjHc6P/ANwjwivRbY4+A/zI9HIpTsgEDLFT43eFVG4mps
WvW4bcxxt4Ojnj/eBgMPDwyyI+OoqOxeEdyMjJ9EOZ6gLnSUzkF299LE4Mj8Wj0umc0JFtPLK932
DxLOZa5GgLNi67Qw1vR36n5JMzYw30F8si5IXzP7FMV9cUD15oyX3UFwhOHtS0JrZnLZbzZCN02r
goG+1zUx26GdfhLierfUS/Jj7DYKggmYPlKQV03kXlEi+dcLsA0xFa+6YVx4DYAFNBGzI3Lge8xf
73uN293FNMmVH0fxz9s0U+fvfD8tBN4M+towGylqMZ45by7u6sFcsq4FQxvvH+Ct7BO9SBB/VICl
iFvqeMn5vpSzR8Jgy9vEerwgJXgBBVNR1UkFoWzH5/YdbIqYYJZAKDPhihclkLtniPu+ARWloOxl
UoiHb3/kvsqBdd2pgULcr4VJNtKJ3/Fx8+80GrWJ2F6B9W/DQEt6apacByKCOB+ANYYOHjPmJjcQ
Flt5aMJeZS+Auzqjtr1RCkvYnFzczB5JQE3njnt+U0bS5Lgqo9cSE7vLBCbrOR2u4480Wb5RZf4/
fQiGpZYr3KBiGbKcOh+/jkz6vH+Chv9zTVoNNR3arHB5hvzOmPeyuBc41Vw5pETuOIdQKx7QzvKL
Q+TbkmCqhANPM/47wve1KWTAw1YTii1QJ75tjfXVXsM8wVUVomcOlpJgQRuDtJoHxAtHpbq+qM03
hCMOYbjtg/FMTXU9RCvRsAd/ES6t+rWIJwwXyzuWm/zIOoaVvXQ3jXsppDHT/I/sbW0BZ0NEzQyL
S5Sz0co78DlPgrYL+28uVqgIMx2Ap1y/tynmwVyhgVGX4sOmZKEW3P8x3T/dtR9tV590ZdUth2tg
jRzH4I+4IjmsX1jU/ofDMxShVpHggvzhW7k9Q/fu2AnQr/fPS0lBtu5A6QZ9R7/5MKmKbNFdIg0A
KnKhy60o60rcYh6/BWptzdvx2Cvdag/UidnQsqkZhaUxphLYrwae3OwcHXaCTAWR3a2wiiGap0I+
MActYLn7sc+FLmxxlX0e4g5Rezl+LKZC/HUyixA9/3kKYyZt2MC0sAWL9LZ2ncy2gMaUtYsRwEKa
+y526EvIGXuaQxflwE6J8MD62QiV0ML+vybY9tfgG7Rj0MbYzZamAFnqfjQDXXjZj7BVdModV+UE
x1j5bZBfZqPthLd92wNUYxHanrozbEvxSaunM0h547VcKmPkp+U0bLVudIv+8cAtWx9C3JAjjM8E
m/rXg+CnRSd8UNMKw8Qpkziv+t0YIMuBKpZyd7qhwjiwFOMwcc/Oy1+Zfg+NCdKZV3vU0yeR3rMZ
7F9mABOayrjTgnwspHLKy6IM2hTt8DbC08tkRsFbeDoJFRkPqEB9FDX7ssVbcxr/J8+fod/4SdOI
Xu55H95UMOO4jExkciumLtxNkzR4aCwuqFa/8sg2euenCfTbtn4upQJLMO4wfMv7KbQumZHSfea2
hVfEnqSg4bWNPEup5BJw+n7pcMklmuZbU8u8gZ39GJf4CEQVbxZ8ZPFmeX/5qHhyhDGT+/MozKye
cGZMkL7wp3AMfXEmJIuPvC8JvSgrhS+yIMwWWB1xKVWa0deLKPDvXMSoFVcSCiOQhI77Z7rddZ6L
Y0uaypkql5tnq+32G+tdcb4Vg64UsFxShw6RGXHt6vzrDbZJUSNdtJWRJCdMuTXUx3vAuqYcU1vx
fhns5J0J05Ug3jK5eQ90/ehz7dW9JcUM9WbfGpt3tUR21treVCX5A7g/U0qxkhTz/kEwxGcYQc/P
AEvSlUfOsxHiIlVeiUR5vVRUEzzNvALT39I3JbQnPn9Oy335u7nsQFKWucs9H4wEKua60t1Q58TX
MewW/E0vWtb0vXJ4M/FqMcrHMOX+YFeuXGmLCb57MPHj+RzqYOozD0aInaBrWb7QZfO6ZF2ToLzr
29rY+sJLGMqAqXKeydvgnU3YfAUSeePwiHiltNnPMAUe4cn0gPRr1Qet9+2JQhcFe1z4Sm2W+DNb
gIf5i9bwxHfMy3EJUwfUC7H1sJ7Rw7+ib/UrI/fyvLdsDWMzSZhtaol1BpV1bs0fa7hThNc82MF0
eq2s7gb31POFN6tMgv7v5rZuU86WcW8AZGGU9eYxJFlhhqjofu2vuNP1G+g2gnMy1YGFFOyCC7/S
iWyxUPuF1RU49Szn0NGkdsUH4lar61jxX3Iwp2uOUIjK7MUex1gtN71wHLiVOoxbjTbaBovsinI3
DE+swVPF5WXhK+/mAlTTVoHHeyM2+6boXA0ZiirxD7JUtg8cnQ68QeW1AKU9Ut/SUoB32UqQlD2T
4Rgucem9Tnpj4TWDqIQGpsfI7OblMT3t0WNY6g+kAbSgWDXr3m38k+j5iMy924GNWsw/fzyUNmTR
npaGCojuTI1VMku1K/BLMbxdBmVAO6W75l9JVR8eO6VPZwDoaKGLgbbUZSbRiNrfXwlPfSgFfts5
m2WcVAjM8HIo/nNQzrm6Eg5PQyoSbkb1az4jb7DFqXFbWjdhyYvTkKMIns7qQLuCc4qGnFxTVDV9
vXnptDi+gDZRmkBJhaNbDD0B3V2tRWO+BvAzHtC/Ca4O27MxMSh2tPDby+JvpTVyMFAK+0jpGknx
DfhQfnpInufcezDFXndoMNjp+h9pPE8Y7exwGXDF/IBD1sR3hEU+DByZCBkNeGGTDuLNP6lHgrwA
jnNo2MOnXHDPunTbHnZIPa3IXuY0Y2GSfI+Jq8QLqGcMUYiQ//2MA4K8uW5FRvqq/qcCyoKAONDK
7DLQWrggHeKCeEGzXLMXAl6VsLtDm5eSy7cGn/oGVQJQcY2YPA4QykuOWrkS56F89MSwgM91zAbp
tqbXqT/hdEbK93x8VeV+lc6yH4vTZ5hk3k8zc1a+TE2TwGwJV3s0+EINFEXx3gcnXtOaXOTy0oOI
v2M/qwjp8Y+Ms2/v0W0PgaykE/l3nB7Tl9vlMcgLST9mOAF+9xtdwTsuRUqr3T4JSGqPhSM/+Dfd
OivCwXXl5G4xhYob/WKso4/mY4xC15JeDUqsldL87TgbkEFHnm3WvEuNMcvJgZnCTap2jLy8DroS
8Xmcz67DxsBunqjHdWQIc9yZbCxqnDoomiG5Z4sUJHSBBJUw7Rb+I3shgdiWFVrho53yF5Wcu9yN
Qw69v4k7DNTwODEQrCt3AY8vygnqZLBGsKd6mwXioi3BKWfyL7VcHP+qprZnT5rFYx8JbKieQJBI
2n+eRttFbncFzFN4q90dyBwTFn+OwRTuIdzvsV60D6P2tEw/pfyoK52mN82dVEiSNxKkSzrxP7qQ
zUa5x6weTs6N3/RNqXev9f+nIzVTuCvgs8WgEPb4dtvcOu/SUzHxtWJ9TZpMh/FWSag073rFJl+C
B5GHpSW1bi4HPCQr1SvjkFmAqdE5bW+03BMwC1NM0TUl7GiewSpk5j2v19nbaep/zWAsye9YTeE9
YstuanF1z8gc94JePriyrI1r0UPoRFD/tOCtOXm/Z1VKULIlkb5aAc3SLwnFfeFpPZ0fN7/prRYe
tonfxJuqzvZUpbxV3PlOhnE64c5HLhu7crspYIYdinwkXGqQrAe6APSWtocJe0fw+LkV085onIs/
d+vBCZ4zbahkwWeNmH/yeUHjoVrhIFjqPZXMMNkAHXMguKY3sloXLYTxYzEHrX5ecNimkrBMrJbo
SYGFqlGtozBHnQs5tp9vCK8vOxHPeEs6weYTYMglpJKfqPbMjK5BxZYnXbF4r6+90AfAfzSJvh+N
mmyZXMMgbmiQmFKebWuHN6ZIIsURgAK4zg0/bU5od2zvYcbMWpK2feHONmVlODPfI9DZ6nqGjlP6
nnf6JLeVdV//IOvYDb5NtE21QzjmTuOul3pJll8P6u+HI9l/wrQ8lkBrQxL/OVjgPFo6w6x+35AQ
1WbdPqHUpSHr7i7vqMK6XEjfJqK77wC8T2td8w0+yBGusyRJkzgis59yWW80n/Pb+rAOBzJ4+0/+
qgDnHQpaSjL4bxUS3A/q2HNcI4Yn0djDT8RloQHmGcZ3WStZIEhpb8N9q9Rf3Nsw1cC5tqG7lqRN
wCoonM5ZFdIXeFR34X2P4zA7Xdmrkicn+DysBAfoEgrkE3at5wO+JgXxzgmL2/rHMuJrSqjYGM2v
V5e5QyCT635HktUZ3Wt4dGusKehaqLk741nKxJrnUn+WFyv1qXP6Jn4XOwR9FUEPjE12NBM7fSWX
lWmXM9bwu94dhws2C0fDzmXNA+rmpeoeEiMuik8LIeOINujtwo8SNmBY9LWu5fNeHgp7pf1YO28v
uOJpVt8QxvAnjpBZT/dv3rg4SN5hfJ07WABcWJxVIi+QqEvqck24DirHWMKYSGBnd3v+r65duSDN
aqsKPlBboC09MM/bN0qmOFgYLkqo5D3BNwXYi/g1XVCvfFLKk3bsWvnFay+eED+cXCbU37pmdFZx
wgsKRjpTgAkBWe1lmol7Zo3CVSDMzl0NjJsOuJZUx4PP2fMkzUr78cjJmHRuxmsXlDp+i4pZP0kf
YXkRhcWYtUCIjEe98VvUDNvz52gZ9+YeSTavwryOUn5o4sSMpIYsn+NWfq9S8L25T+1w4o+IfDg+
rBudDydIktPsrjKVSPcJpfb+y0kAbnantxAPQXCqeAdgUB8NWya5WjHxJWv8xXs0pIUhofcHapPW
5uvvuipZDLAKIBACy/eCp1hVLe2f7wMqLvJY4kELXXs9JQ/9pVbwJx4FGRDZMEcpx+l8xYHCFsL5
QRcj0WlupbHxyrNHCZ7rFbiec1eJ+EK14iCvEJKHwQrDKxKFAuX9zQR1bR+7SVKt6KIDaWuc2k3q
Z3FXCQSMUjAYTD5Bjgik4WwKeAGcigOUrOfBP3Sr9UIQyOfasMWEO2ONZ755hZrelHqen5ThKJll
USBSxAyuqkrmbQA2UDemkiyJpx4MsVkIzzEqUeUyFnWOdrfSTF5WwVAC4sIEsYWUDcz167VgC3pa
KXWb7ZjpBM2oWWF3y7FFTwvotIuIwXKB5dRjkh1qZE+MAhbWooOtHi/U8Nd4o5yAhg9/cKtYBLbH
rGs7tus34H4jlGeUBQS7Z1h6poWgM7lsGz/9uNSkYLWz12EbnOCkiymia7mlewDVpVkE5BHRuX6q
7/LSmURs7osZBu9bsuA5FTVVbmGtMx6/qSD5qqW8B83zk88l6WqfyFqf30Ba8dylL5vvseefwdoh
Zdj7/EQhm3qNKnWaGzecNM1QlaoZFsuiq+5R6kdtKX1+51YhvGq6lX/gFaX/1J1cBTNBJ6D5a65q
R2e/nY4fKn9PlPNr9F1n27sLKge5oHkY27pjhGk6zxEEDstg3hA4+MhBU5r9IpmJpxRuWf0P0Ymz
UNHL0ruFGrioMBASvkxd2rVHQM0WvkVYZo8j5+fTbgJkCQd2l1pSVjwNkf4bLYZWAVjhVjnsf9JM
pTEh+mS6/oXIPIsVkTGgEq0552Blmfx+tSlut3C1MYduqY9oQ2BzFnfLHg4Zkb57R3H2jBGf9UNW
ADR0vWxIfXZqTlX/z92fxIO/MVafV8kSih3SW5FAj7PqkEPx2hTuovN/ssO4sJ+KwGE18QN1KUFF
08+VahKWCEi7DDRui3EZOXZ9eAWu7skMmCVVHylQiqm3V4hl3vkUe3F4GjCpsDju/vSGKO/i0FDe
Gg9GXx/L1SrigZq3OR+0FyY8UsVcCeb7bAPQ3R9OTlSLuVtQhdugZLjCAhP9ryyFKMvE97S/GhaQ
Xic6x+GfvYFxaXICimTkh+drzdhLnq7WkL8yWBaKyAa+x6K+n4t4DBXxJgpzSfxIDBGrO3s+fljk
HLOVA+tGr4Fvwq2chTpzYGSHaAfZ2Xcxf4rCOEB46SXtkBn7XgKSlxEPP8oxgkovvIqxUZxhJ1tZ
9Ie8odQYdvOxPqFZld+Zcqr/JWpgsvZ99ERheYFWwUEsM60MJmm5G/EBgZifR8Nh1raSCspAAHPk
EC2Lf90DhzXye+iMASvgBFJgQIJ1NyWU+ZBXFI7zUuZqSHYy32p49KjDgyC90CW72NtraSdfy8BB
RMBgkna86HARsJ9dBxWVf2WDc2oYyrFzXuv2wRI0HOt4M5mPRW1fgLYRvcgWwPWqfNlUdeoFtpgh
5CliRNSvb1nU/DIQuSuD4jFPO4i1mhWDCiL9yyPbFixht7vWFiKmSbAh+CvMPRee4VMgHt7mHLu5
njuSi8dPLhCL6mqgu9nl0367y8FdF3rylFsk6kG3lli0bsoK1wHUtb1B1Cct5G6d/JLGf/ntySrf
zcKpzcWot9iy24HcgHM+c0zdrXvhS/N2tw9wK9KyPCSgtXXT0SC+q+Ylt521wCvdeULzPHRYDKpk
BZS0lks9c4LRNkI6rdLkQyJcgI2u1o8LNlJ910URcKFpe1irq0+wNnBxt+5tBvoCIcu6zKuG66xg
GKk6ap14i6paXg/ckoDRFRGk0DVg8gzYq/DoZrthWre0NuQpR3SkeeEvwK/MvC86TMf2sKt7bQuU
oiqCIR3hsHdToggrb41is6/AjWlQH0H4p43QkfA5j+sXBqj9XK0bPTj8u+ehFLokk6slYaVlwH+a
iKH0Y9Xik6m3VAUldb8IeNmiFZ9BHsndKRWg0z/v++mE5tZGh94SO1TaJb4mLlM9XUX/KRj+YUHy
rCG3HGBQbr0rUFhPdCwkFlnzeXpAH6jolwZ1lJ54X7X6Bq9ZJcmxjEL0T2nrmtyUWLJgI08mc99g
42M+n7JF+wGlEr8Wlw1J7QD0yWyzNaXttxh9t2kizUAnikjR90uLjZqzKeUhmaZxzPLrpiFq//0g
58VP/iS6OwKNU4gCW68r/KgJC7c/yoVAW367d78XVpVIZnk3YfSDYKbrnbvz9+JU4mphyOCfUeTT
D7Lu+4w0ZIT4FW64kSXSb6+JYb0VuYeXUiwW94/UnMTeUnXey7qzsneBNyr1IeMt8MvSirw42u2v
MclfoAoEJKVzgsiSxcwJtrjb9/PV6mEs637fk+xDe1rZgyIpE+5MYHFgDOOtGPoidInodix/Y5EH
NeXO073zBfXyFyQeSNmM6KZY2tp+zMr9YbQxC1vuE2FHCjcVuQivhQhk7HH3BJgdYMXWrgFh59v+
iRVeDogSsCE+tL5eP32Eqltf6UuRbFVW4pY8JkED9cA/Npdak5fEp0bmto9wCBYAg4ucrmX/nDfJ
0c1M3UnpQnCYHJN6vrdfyVtOc9vQQMmU0AN0BiixbTVCBwblrcw/2mNq1ioYMl9gPdrYdCUGA2j8
SrgGhr4Epwv+bRP+4rrsXVh7txAOfYSV2sxELd84E1BMD1ZvAlxoBBhlpLvhG2S0MIPxWJf93I4E
1GsSXaOKmCM75xDqUb4MvLFrBSxtO/Rq/D4GrvgcZOeGKIaaTZ4cZQlinqkYo+xkAcGN/f/2x0zW
JYNQCSPRvO2TToadjqhh06uXo4oAKZr3UMTSe1MP7NbVZ43EyxV8vlRuxaPVkFDc7LR1HQ7YdN8W
Y/TP/FyyEUtDsmdr8fKQFx1B7XyLzX6pweqUwonWw79DkKr/2lct8HFCdDbb3vx2RFc9tFdFzsd+
apcq0hTYer8DhQI6tKl6HqmyA6yB4d3WOFql0NpXcVGv8K0EYApcwohP6kDvsMRVVHDamgOPHlgP
qsb7ih21T9AdbAkdSEWFN9tQiyNam3vi7fyCdjFhT7EzfouUTk/vATsy0HYSjNb+uT5fax825EEK
wdRxb595HM1z1UmKMYsIRxF2tMXhaCIlv0We3Zu3YwK+jv5sEEClhVyfxNUrsri8BbZ5+KLzXPUt
WywdIhbj0QMc9AAA7GZjo6X1+AnJar4SGAqmM1y+1V00VpkS+1DfnP1V+/9y6u2ShoMS32tcRu3w
sNEIKocr/A2esvqclexFuHpSo/ZACaS4Kum+/nL878QhrYqP3/DsyL3yGQAhWlTo6Ff6FHkS1Jqm
gLaf0TR891tjO0ilLfHEiSIPkS73bPP+02yN9aPap701/wkX+jRQG8YJ5U15IRmqUOL4WXoTD00S
YtYW2/nSyC3/OH4Z716J20Eotg6MLys4zwgJOfXmV8udlC3Ztmv/P583GHPjzjzkpvuwHD2BRatD
yGAsZIo62cnaMs2z16VllNlTTGITIAcadEa6H4+e48AfaZl9mFGrRluV1Mi5Kb6J+0QuwSFuNQKS
xJNftiEknh2rIcT/QslJ5wp+49EKqBqM+PVXttKiCtjWfjZuI2kN6oru5ZZVj9hh0xFFhDdHEAtW
Hsvr06xCVcDOC1TznJVZdgQEh5mihhOTe14Wnp7jTpPMf19VPGCFB0vk/fbbIf3MefgVU3+EQwCs
pPt6pqlVy1VzFgLe+YdkRFa5MFI06ECykQqPH4lwAVcnAK86HvH0CbA4nY2wisFjZpzeLpIo7OHj
IUrrz8FcbEYPQjPC1/AyJNKJk1GE2/XI5054lVk9o/hbmtF/DZl1ytNwA1jtmsQzMJchd/6pA6XS
Fh8/H7I3Bku3TS+SSrnptyudG67TWd5+dVmopq6GNJENaQ0QbykxRyfMCMn8OcDQZE7i703CN3p8
hBx75Wffy+P+SGJ7I1xxNfWn+RBZzVOViv3Ajkcj9DjkF3+rEL1lHyZBmRLbWDzvuPxpg8976j+z
Qc3KmMl6FkWx8JvbZ8pJX7Tfp6Xout1h039UwxSfp9WwHAEkvfJ4dYf8J4ov60gIVPcn4TEzmHZ2
BA9jWIAT8rhweY4fg8h+wWC1NKDXiOCGj1NzcTEuW/l8n7xv3T7rJ8rQ+v68dw4hlRdnIVNNLHOi
hxD1OXkP8nHoixAUSW6MI9UENejBj2caqzWUJj/FXJvOy3BQuZ3shmycfnxTmRHTYpdv5Bp6Y9ld
8PJ8lcjyeXhmIXvy1emfCNCVc7UsX1JMGasXhDiReOwK813rUueTNkPh5q1kaucdkooWG83dFSt2
FAeuz8YMGz0a0bQXPag9oZkjWtjOfOPZNH4xD2gRGwKsyhxmtIRHdwj7YW3p7xHP3DslRnlBeQUC
8cvSVls7iczyIwR7/anNHaMG3Cr5mpT+5O6aOsQprTg3GPHIjWMBmA4Iix8yld6oEAEolyiiJuJG
/jfL2PmIFOCae5qrJ5TLNmgmefvXdJoQMDY0BfaY4OTusqYy39LdSlNCryyUU4O9QjMnkoSua9Zb
qzCXCMaTHWi2liqgibYAd73UxLSUkG5+iKsWk/MhvuCZuNtMuDgWZkeH9K+mJzY3DlzLEdwpaRJj
Vxy9lR0KVjY787PCmP22yOFFawnhrCg16lz5IG36Hzx+pUT26DMeVCwyLECeJiCGv4mZJM8E3eMX
OT9SjIgzVbJXe5tmzjkxu1f0U46mlaX7J8r//HDwJAvPIQXMsNNXK92J4glNk52JHSMGndk3s/ON
+/HlXP1EwAnPaLjjJpH1lZ5JRkECwouG1vTMekCr0c3eIs7mItocEIzVYkhZRacta1dgFla/PsyE
MWQ9/c2RfZLTVuGVDa3UZ04Q2Rm/9rPOMxA5yiw15O4EEVP8/F6iYqAs3d0s3ZjlTs+FNQz1YvR7
WTSPRksqeGWfMw01+RAON6LT4aDa7sWEVN2hHfRQJWULBBglIJSdGBM8OhVvA0nM2bLTIrmpTb7F
V8BDBD0N44NfaHxv4Nxz62XuQHuy6e6IxUMbAkJNjQgc+EmThPv+vhUBJzAlcxWffRtX3np2ALRG
RGzyoU4WTF1nZPofoPdlwEZPjVGfeNEKF5r5VSGF2LyxKJ1UZ+9N6vJ/QmbqZemV89m4t+DJxIXN
/Iov2znMsnlsYAM8BFm79uv+n3du7eKFVQ9sOw5PmgQfxq85CKkLuh1b1VQ/+F2l2bzQJLQaDTrs
tZfSntd1xeIKUCldyfvHAiUF2wVVgGkLimLzIiovHIPzMHoE+2OGVjF30q9OkZtHgz7IDAJ6IH+n
VNnoQInceDI007Lla8SPGbwzKwl67pK5ajRI2LMy7NS+nHI5bjAKfiXgDuIz7j1GP3l2IUysSQFD
iEFazeZC3SFVSlkmscxRyD6IPnws7di+Sbw1rTW9o4MYwHp4u1FnV9ykgY/eXzOcwj9ZH2QrRGfk
v35XWJW4ZwcwZv2fp4CW9wr4SW1uct8t8GLJT7o1ciA7aUZV4GKa3InRsII11xoftXB9AIVcjTp3
bnuST/UZqWpOrRSa+JFIjX+BhPdEZn4gyHdAU9ZWXCM2WinwliDDb6KgWTxRdvJXd/Rlxa4O9ZBR
ZVOodi0MsR72mthsUlREpm6QBICHmox+8AO4+plNNnu3Ifqg+bky7wwFxVw6Tim6Q92I5t2oy0Qs
iuSh0RgeAtaDjRQjoXwhzYWYkGvu/mkZ1F3rEHfo/wcGoZE/gSkYIbLppN2hlM1fU3F7yEsDzUjV
XaeukIXpA3NK5zqjz3nzxGkgSK1MI53qmjbr0I0R5jI7tBilfeqzpO0QoOHRO+colaiX356iiJMR
3wo11VhEsXwbJMzjs8BiGjnWG+Owzs+4HQrCM5hT+X7Iz5m4irYRVlt1gwxril2WFgd8ixCI76Ge
L0L855h/ADIZJ0E5q2dn0dJr+MtkeZqau62WPXsY0w7Nh21+//PuJF1XXQPDidtN9mCpJBrMY6jm
busYZVrgqXMalJE+zAxJdAcWy6Edf2prXCyMWbQhtb8xtRbYGmcF3HTz7FkfqfVx0nUkWskrVriu
m9RKoGQMQTilqvwxgrl7VKaeSwRaFSGyQSUAoJ2SMz6AfnRTFrRZs5/1SRHrCiReNRwtTfSkCBu7
rnkVTpMGOunWx1FRxnGH/kthcoYkbKq23sZx7sIN2k1zW7XfGxrqxutPWi9XLVzWIu7+ockdBKqX
AsVF3IfKdNvMxUi/pUg48nVMPQR42i1ddfke6GYkzDx2SiYmM/oTaqUWEVdoSxhKPYrqzrgJvfOm
G2PPMm23Rb+HcBBhkWTpXoeZ4iF9TxzImNYLndV5aL3ElyzCqQ5st1C481S1NJjyr7EZAylFx6MC
K1i9j00LwqvyvYxMulYclU1EWqqIUxoCGxrpqpWwyrpmUdsbwUE9V9SxKcQD38QcupjqGy1uqRo/
PLVhrkf7sTsX8c4rNWQmCWURN7sKXByS5ZXU422G1c9u7CODeksjFyGsPYHgLO4HcTkJl0lDjLLO
sPPO4syrGJQyQziNvdr00g07WDel3JcfUb4SnURRyhCLhpyQuEeAZonNOGGf77N6iQnnpt9GT5M2
Su/S5j/wC2QPUMX1iHefdxeSEaLuaMOXHQww/Fs5JgwPOM0E2RgN9m13n3QmFQ1ebM0Vat/k4WYh
CtmqdoYE6iMdKy924fCsSB6sCgCHR/sC0+FpPDnUH1TFGsGP/tfUcAiZbqHd/eB2Xy7tJdCqr84r
LMjaS/gcszaN1SoNWDyYSWzXyYMGVRgNmvqMH7+MYjsIsAhBBGJfWBnUCTENlGVXMznoJh9yiLBp
oKdxBgpz6ddjZb2IZ+YXPjh3l2A78R6re4vM9YkvaiJushi87Rat/0V9OQTyYzp1EtAZOvjPKxRD
pGmmpbqr7iONVinCqaZWITaROM+KkYfGooi/9/X8MaFCHyrSIxxigDULCQ546Zlghg02g7TmysnP
bfBErbKTOO6wwU/Yu/oh1qFFzGPzRRAZaHwQ6W88BMGMSi5ynEdxt7VkWueUQ2NrECUiwa14LREM
DYZk8ercm1MnvD3RIF9zmQxCaH1r2UjpOD8xbjGzZ8cojcOiwCyIKO2Kny31Hk4OQbeaTSOWaDLJ
IjJPmBLPKYDE40YMxAS+WTO1OYu4ICunhNtfLmZyeQLzKkgOQTmn8yifx9tCgOeDbyEBbB1ulY/k
TAeJ6I6WNsrqI7eK9MadlUitYcgYAuIz1xhYLpmhWYgmlmxaVIO5LTcGIL0kjHotK4cBEAbNDfJU
AVthPq90SutEZM4ce9YXO3O6gv59pD8Ua5qSZx2Asmq3+ncDnpHZ4E5lpqQkw+5fba8cGRPIzKSA
Ry6sZON7Ag8SgMZodD1R/pVNFvhbu6ju0pgHHTkezEaeb7mGtjv+hsxeJ+5+ajIgRiWTV/tW5QVp
2E3k10CeC/x/l56D/h9AM9PKyq7ctiAwzyGYcTEvaJm4EIuP0xQIij1D3XnKiR5Zy9fibKeVbkZs
H+zlLhI8WR6sbPcaTv6kk2L0Qx1SiRZo8ft/7ycKNYwUp6rkoP2Cokkc0XaUYBCb81n2ri1lhutz
fGUeRvCb5aZyjU/agp6fkSH2rSca53e05m4oZB28m8qospi29EyR8ov9C96pV+REXwxGitTGIGjd
se2tC8MFT1OOUWYCHasY4A4SVNfs9qkokoetXjex+xREZeAHxx8oDg1jJ+VfnrklS8WXv1Ko04ho
rB7P534hP808r7u5oTZNAvQZEWIGvcxvnD+oj6yj+TLnJatWkdF8GLz7vCP0Y5IG4TRTO3gjqFoT
4Vtt/tVIid8jKXa6jbDw9GT9EJI7qmkvcHxeUl6ju0u7D+Vm2GZZ3c3duMKSgB4nfIvH+hb/i0b0
NvVeIlYzCVswFLev1Z1R8BC7Pw2lljfdKvg/yHQl0Tb+qFitap+k7c+6WAIx4tSKy+J3bheEGaGf
8B2JqZ5+RP8VUBgeg4XSg7uWEdn0CdkN4K4g2gEzHeZED58MKgWSvSg4PR4DD7Pk0cPLTgYOyjwx
MXAdGFBFwqbITFtH3vxQBo6tMANhzG0QpuzxNpyeJNy/Xc/cYu28G4QfH1qQOnT2R0uuR4mJZB1c
U35xiY1PRiq3nbnR7FkgNqd0iKmLYMw4i4sWlzYY7H5AXaogeG3l8LQ+PN8OFHSNHSGxbAz6ThLJ
TW+rAOL3LHUW3oziNHiLh4Mk01SUzig4ET543o8ayoZYRqJnmJ3tet0dWwrCKv/npRjgLLSxYBN6
z5m8KSjwkIp9wlVtzoQL+S/GSDMTo2ZRJ8wgp+aq1fIDkHy5nGlD4s+EBt/BH7nRHDC3ySMbp1y5
W0xoQwUkQ3wu7lRzqOgi9DRKDL3D9jlzH8hkLgxr/kEHXIfJucYxNVWTRzunNoiXEaxWZphRMzRE
mucIX+yczwsEmHQU66K1E4zAuufQent8EVbVsHhQgoJ0kKTMTOtsp5Bdbl2pOQNqReyWuVsELso2
H5NCkf2wWzI/RDXYEMbCxynnHgUC3dvqIBPTF861n9xnlCIUJV/UcB7VKcFYmvMROH3G7+Rwr5Zk
e1gf20HHD+LdunDH9tBA+XQ85noFj2cr92R+UeglXihdFJHWlXCwD7gpWNnwy++0JGDaEcHuqM2F
/COTCZzCxGcQSEuSa2pP5ErwLZ/iDlHgw+ugTWt8HHa6cqbxoT4/sM9QTCu4d06+MAwjUthIx6Co
b40Lhag5sR9XytkMMxFKr026fsoIKAM0LgFqTed2DRSnJ3hvtIcvbL1ikIIjPNTL1AP6oGW6Bd92
if0fo627+y0Hc0B/xMIBENEEmDbK/aE30zPk5GW10fap/DXt+KnBK9aULKVRae90WoQXodgr4+v8
LEryeE1lxpwEi/FhLYSnEWtMX8tCGIAqNhhTz6kKDoPvv1F9Fh2Q3TeOIUMcM9N7Rll284+NCd2G
UT57YIYLlmsvaicZImTbj5e+mS544THQ5M2qog2Ki1+Bgb94B7j4SdWOvLbjgxpwVRyGPy6IsBhF
1qgELvGIXtrtFgdWHLTdTFZYlB7ET7RwYkGJS6vVzMCCjJQe/0+syewfYW1Fxahg6i5y9tk9yJ/j
+EhQrAHIgQLrHAgqjk5yS3JO0pkhzhuGlEPy6Hm/vzvi2YT1DsfHs8o/6LieBAN8LSkww/JWmGJB
urR3MKK2ntRP5ZPtWZ9+KwnQ0+T+ClSqK9/oWEy5B4oqZH4ZsGf5Y3ygoKSOZ1LiPp1ZHziqCu1V
0ddAUOJqiG6Gblrhi/iexM+NL8dM/sGYSDCsBp4aOpaQ//+jozoUJ9TUHK/XE+2jcbgnHYWbq4JF
3OV8uisQJOpYAlPrgj4tqtHNY9cOULqQPY/yEicPhVk0CZbFlAK7gouIUnXSdp/eiQVtm/sY40jW
qWprps8icBU1dbCD27ZH78b4ms4rWyRy93AkmqBAZJnKdBALif6P8KosCK3coOMxLjLYK7MzATOy
F+u6jHTgDIdGDV4yalzRK5ueJ4/6yF19xUqWaVSJhFxwVjzSbmp/Ee1It36qGNlner5waxDhe8f8
ZpAgq7aQCCm4w2YlEOZUMY4VelR793HwvhMORTXx3euICr/np+xq2B+aOaByEC9p2331km/qMOBw
4EOH+3RToL+Re6OBi46rGQgs2IGJWpKIYOlP0jp7zWxdiOqMyhQ99HxsOPynGE6AvfA2uJjfY5rY
c1Cp5H0OfY5+RiLdwAaxbMOVSoeJHSOoAhB+1NxPzNI3xPtEAS8nrt7O3GQW0O5+PkMzEhHCb+qZ
A78NEIHvYNEdnRgdCAFylaL80fsJjhpskfxTqywtRwA2iqZg/jSF9Sq3TeDIhSAD+SD2lehggMEh
BdVC6J5INZLHjsvCQNMmh8osYGqIEQgJngTvzWlbBRbMnbB27M6En+/MqyDOpxu+i7Nb/Byuj35Y
dGYnKfAwhaPiStDP7lANI5mUSJ6EzlwFK0n+MBJZZw0KqIMQA9+n+qnwz9WzF10Fg0DF5K5r3HuW
hQp91X+Rgs4eAkGrwPfdzjToYQDgDfoBsij0WYxt6P1T+1jmzZ3tR5+/p0gP5EvreWgk5XazBvI6
4K/n6AC31HVELp4kxtuIafqUOc3x8xUUhPPVLHBsUQ2jdxC756kCBSUsrfH8sSSGY8A1lH6zxljo
ftLbhvHBbXyfPnICmdekMhgJW2WC6mxvhDXbFrKZxFkGJD6ywTxZSX1G4N49I/ONLVJL8uL9Eoi/
rSALuoBEH1EmDOhKBxjnhj0QZSfBYmQTgVgw2GcrjzhsnljwwaYjAuEEW4Z6yFO1HbcZhM25ARku
utWniZE5IBa27phgytQ5X4iAVa+1OqLjKD4Ki1ioqOorT/7WHJZzfafgsV2318/3iMo7tyoEE1Ow
eH8+HwdfJURAwwx47Oqx55mjmNF5IHvxWbSUWKt025hkg/v07duKUvz4QiZr+MhYsAeL2Yhx3oBR
2x9cbxwTkTzK0i/iuPX8gh/wwGdXjpot04al8un0fQl7ZuydpXHkNjIJGkeLwDzTTDNVJ+m6K5aY
M6ZFJs/0Mr+As2IIxJfMyJG/taZQTAYQvhaWo1d162uowdxeGRCJETCVlNjOVtPVHfOXpjyU4q9q
AF7bmUK/fOTTWhdv9ZkYAHsqMDUaam5BreskqBpPnUTrLI+lGxytw6yG5eg3q1I7o0obMHO9Gk3e
UPPq/be+/98Ue9Ft6cVZj2RwsGfubMitWdoRSsiSJfnp5e4pQj9y4ySYJvieLmrfoZOz78tbE2gK
jSNzQ4QecMvAxcpZnWdnyJJYl6nZp2MIIljDdZ69PLHJwRs1hFkqkTrZASJDXVQzXocjw5v8eYhi
tBJF3ii4/D3oiVKoSWkq26roQEnvN0rTxhCqtU2k96G2U2zGJ4vHE3wQPkDRD6CMKd4Ro6kiIBfh
Xc1B3SzDvSUV+IHspypVFGUS4zkoKfYdyAO+PIOT0m47QdGXcF4U8FKBfC4r+Sjjc/ZNplGHUjw8
YQQQHRJOgJh3bh0qZvHAyVO5vSwfw/nI4XrJdlhMPT3J/Mm2wsT3YVefV4Iog8Enqb0oTE/oDs9+
zJ5ofKQlk1Av/iC8CjQtlzj0Py++KTyXRxnVykgJS6g8Y1TDUcR3ejkYzOKJmZ/CLi9vfTlLq8mG
2PbuiTA9kWTcqEOR5iAZ6oMyH28CKgMhiUa0hcfSX74hfo8GYjk1ITIAo9o4tizvfNS6zilkWoD/
RXDfXb4Llzeh/WANJiqqmkRNbE1MER30/pXPCla4wTEO9QkVbihRreRd+D4EXK4Mv90IP6AZEvzu
g4cF5nA6xFIa7fGiV2NB4uWKGxjKuBBZAl2oYSkAuApoSl2314kvvMKJCcSwyeFB6+0zJ3OIgo7h
DQJr9wh8LeEyi1btdZeQclnjI/LOGPKzJi0DncL8HqBm4/uaqxSRA0E+LWXyFhJ8rCxh8HkDsGDB
l0D9KjftNou6Q7dN98TFw+tp8uD83i7wDkohfN4Cr1bSaT7U++GmN8UaLib4AIS1BZglQwxKHRud
675uwCZCbp+wjL3P3qkOWEVcIVDJxHyBfxi5/l1AnJNrN64s+yC8CTYaCCUuTmjVTvHpYHjpUMUk
5EI2wpp9fb1F10zYTt3fnvOklpm9BeDCDrBler08UtIeMxNUCBN8Edx2aXDM6cbLWUrlMJV6YWLQ
nChCe78ZlBewcG1e89Pu4UFRoXaCoPWT/6rcq7lrLvrvfCyJsqbuSxDiGzdqReSQnXqeuO2bwSpN
R0Sg6ntauwZsB5RZb8qXROW7oVD/OiB+6iRnXaYbmowm+yu0n3kXkg0u7hUErgt3Q3Q+n35IHGmD
KKpbVQ8RrwBkRV2jX02T7vqTOrxhetdLY8kALTkmb5P8EK3B9TQvURyPr8PWVLAw3YvmayqAUojv
mV2JICtwQjJvb9Gu+J05T90FYR7ASCzpBrsOyUk7iqsTgA8zNefaZ6qbHMKHHCfPY+1GeTmymj5Y
BR6j2BycujbzbnF6RSc0ukQQ/Gk7cy5qEGEraihP7kZfbglesVP051BCvXVkPousGyXvZRb6S79N
fFu+HmzQTpTObXPtaDc2LkGonFXraBv5ZS4vmtbFbDKczo9cjox/tklAdzFaJ72BQaGtcE5QYZdg
/ZT8CDqsZcgxQJOxuOdtFydOXhcn97HTAltYBQzyV1HodTP68prSOYyERJnzsgo0ojMoEYBhFr3P
qLMYCuNRiosWtKugv5qX071p/0aTCulMVi5isogWUBkYKjJhwHJWm3o/CT9wNJPm29WUXgXoG7i8
ll4vZRrzn6+8+SDJ+M/mN9Uv6Hpd35KwSsQBgprBAut0UkYnLIIDMc76ChFJfAbyji6RTaTe57sP
FT26rwqJtysiFyhdFaAWdj5dkMTIorlPOYhlxq9TLAR6d1OMRkQeqzWe5rJUnUyM9FBzrvT2j/Al
BqQEnuBn21fk/jV1ZHKoP4CRuZu/DW0mG+o7sGgFM0RT9tp2UKKnly5OEjOPZhaa41T9qWol27qj
MmpB7XuSUqUWCInWJrD20zQ8kd+rpGnXSCSxAKGxIKFRYQ5UZfTKvaG/uArWgkA0ylQGYnieLDdT
eEOb4mpy08+R0aYNIfGO5gz8tmtK1V7mp2bs3Nlfl9QnB1AY0lwHixyBGgGGNuWVlFyl274md5lP
/tLwI01vHmAvu5LYCYgYZpUNsE/LLHEqrD/qEfjm5H6gYDc5mu7T+OeQAGSqC5exXZc0EFgzkcrm
A3FyAgy8zBZ2RLzQF7nnMwn2caUc/PjZTaX5kQqBiMd6qPlhAkv7l0oKzOyBVFubmRjk92fb8Pkj
G+PO5XLx2PkCQA3/FoyD8yfEDynCdqYj5Tq9+0OfVskF1JZMvrpsCZzqbGssSNuH2u21sWnAMICD
fh47bistkzRhhtQPV4BfCixSSIxHuWaJTcSqHQR8zPkVgscEwzUkUVMtsS/wHtN/2RGNeReMJIIO
miXDdq+uGf+OJhFku02o2KvH15lwP/1Lc/pVICpmArbOuJNzbX2LVitBt0QhSFLp+nKDOjGUK2Se
eK69bIdGRjmzgFt+3MrEmrQyr2KhLqUW8bMxktQpPWn6uJ1M0qXGEc5QSkIFiF9ErP74ndx+7h2b
uz+HTUCnrwQpCIgDmzir9aUs1gDrLBJ1L9GSvObDr7hpJkjpqChhh5zAcP7MbBHKWJ414MveEuIA
qpKewsUlpvhJbZShSexmHbLrXJj4zcs9BCJKDrl3WrEaNr+zoGI6qYWfrGdjV6yOOaBt+xjXEO+j
6RyWvAPFQCGPN13BY5NqVD7DtVdwTlKDUx0hD/Tuxp0YnLiNo7lqMDdA8UskLCgehUVFgK/XP9O2
QkyeZgeG/ZaC1af/DNlBRxNNGz/e7a8lBoXy4juOPQXokMR/Bhar/AhyOggpNQYhjJPVsfNoMPUS
KVFnoztZ+XOVVaRhzKhMG0KU19e20BUwxwuPsFkD1tA+8N8n4lEWFp0Ew/hD1eVR5eOY66poOK+8
D1pWxQ2GjZuKA6D2JLeEfzVH3HnE4ouK1VMJRiuP7+XCfwJvKQedY/EnTSOBEfwgAlZH1H6mziOB
C82Y7LolHJL9rOWwoOA2V27itBouMYYSLzVktmJVmKIIhubG54kP/iPLso8fGkM3bIpYnFMjiWdh
dZxCAN6MU/NJ0Tnm0oD/iLnJ9yGS52BRGv8a9rrn/fkjONa9RY6v2s+Ack6RmJpbQHadya81lhvc
QiBtqh5qpdmtTTvsIytjHZHC2cxP85xXShURscsKl2Mkwwnoe/em7cc7YJ73gCmWGP6cpBp0+aXW
Xf0pdtBTN9CwKtB/jiIAaB6KjxcdDqnxuFUOXS+TS4R3VFRKUAnfd5AhSKSu+wFd92c+k3jaFMdK
8jS5/eRyyqvzheo64yvL2Z5YGuChW+vqnY1ZQMWac7SWoNgc32vlZ/6IDgdgJPFjkVSgED7ZHG/b
Ub5NlhNtJVxvXXvQZAc0mP7yJmE4bbvymA3n+q0b8LObvtGBkC1x3QuShxQEN+MtyIVLiPOU26vI
oXJZNt28pg+lWmcSHnlLzIgSwe8vYSENaevyleEQvip+nMNG8H3z+DtVktyOsJ9d2snu5MkGYVFD
e3bszhzQGqb7zgmeAfpwCKQbUxyLec1xToJR/p2s/g/0NX9rme2FXVdAwONsg8bSqsGavFwoMHYi
tOWi6FferlpZgec1BHdP9hC0cQJXvjGNbPZhFGQ8melGZaX7s00zBv7kKrlDJoj0BOvdS0wHoqFU
3wPL4LqLA9zgG6fYbna7TX3Ebhciv+ZEA32gS3RQdCEheDzykSTkxwb0boKFwF05Uh+fLY6Q1Kfu
z7+qowDe9ZCcY1iEKn0iiwWDxJLQv9yniMFx1uV4RC36Fu5q1eJPIvRfRWBV6Mul8QPYSIEnW3yj
9U7d+wikvgoC1jyne494G57tYSgURKM1eI4MYa5QeqeWrMp6EtZi3BVH1N9W5elJGPp7Ei0++tKr
FXQ/9Z0AIejWbXCgGSwhHMk0oAM/wiO/9xo25lsLR8xDx4AOvTfzque9ubP5OcCm6OEVrqu0uFtH
BOY+LSVPEsKlj9IqNBaByMy6qnlXM2y3Yc3WQzVpTsYpIACb/xVGF/R4mJjKuipJ8x0hxs5sn0KR
JrnbFnDrDABBe3cFgoN1clMdpeNVB9aU0/a/sYI4NfZUP09drnZgeWlIDTVDrMvbO3wdlzTT2ZkH
e9ZH2GKdbNFmgrTpwxmX6LwwESOIcOb0fNyC7Hazwd28nDUY+6/sTzTU9pXK7Z94gSW3nT0nye4o
y7Ob2rtiW0mk5nn+gdbTU0TB7mGSwBxPLkUJaJHa2fZOtxmepdWM6XSPunRL3RQBH091QX47uRUY
Zu/SdKZuh5sjf9NNnQ3KPA4dOBzP8VPLmuMXS/TZp1ZDGiBaAT0wGkfRsTUks0uB88w241oTDBX3
KJm3OUF384NX4NAqJ7KWMvhsHiUyF2Cb6GK6jv69Ma/q+LUI5a+WhOUM79Szbv6v83HWucCgAZ8T
aapkQ3NomxDgwuWqrY84KJA3qU2duL77iAdH54BWccUxx18o1XX1+7OEaULv2hcRUsZLy+2dr5ZT
rQNPCt137+oxEjpD4W+AWwQvNI1GUU0IIG5zh3oCCBqP9wlttQWYzwMb8xI3GIGZbgAE1ohUv3vz
rNMD2thvRqMgfZyyvwmrt5GvsaVkZWlWkXaGJriC4Zb9XB5srt+E89kP5mDBmXTAhROkrssqUO/9
aGd++mqMH87uyPruWSng5Ov92W6GhF/TOVD/Hp46wY37+XzpVCNbMjUhCgnhzsnygvh6vc13Iqzc
qhDDs9nhVhDgqlLRSyzrO9hPbAS1n2nKEWgMwI/MBTOgOa9ixHRwkJusIztzYHPNNB1D66txZxNd
cY460ryL+SIX5jSTw53vChiPPxSvBmSyyoLX9kPYYgzCSBjM0NkRYpa7RhlJ2giCIeYGqn+CKcZs
5e8FbvW4mz2pB13rbxZALtoJ2XB3f0qyWj3HyRvGbGjeGLfGfUkqZThItXgYcLchnZRuXRi+BsH0
jYlevEDhRKMDjk8fzWO8g7bd5g6UKbsQjAoUyg/4ZnkEp417+YyCtxTWNk43sGlkO93smhhKHZsn
5Pkek8gW9s1/MdGadVsk/L9/NpzXlX55E3/lCbpc1HT2ajVDIaR5C4xCH44wHg2JxVSgmOvzCVxG
9sgfXF7xWaLUAkJ3aX+uAzgTCS9DEptkjAC+yMnqEVbGwr0KD5DqaDGCodXNqymSkfbBNG9ApJUn
TRw/UBm0TAo4CGACPaBflfK+vXdnub4xOT+DLc3d0P85iBzRhXJHQP9S/iSIK+5Y6JcFv1xsxvUH
J52WwKBg9TSjMvgpS+07AISkNi9mCLYXLlP7PnydTqsUUcV3l/QMsZLnbGhqxyV5dfph12s0h8I+
CeABP4m/cjDm6Ai90qnmDK0bZRI80J/qH86uEedd8YV66QntiuRXoe/kIHo6oKhLIXqlgZ64zVGd
WVRrR351jE2Y1cYiWQay8c9kv0nEjdowu6SVnsSH8TzSo6u+r5N5xoNSNFdcJaM0TrTpjfXcyfTv
5Et46yOScXf0Zws88qDPWWiItrzno+RCTt96YCdjqvKM1GAnFH8OcRW3OLWNf3oMMJwJ3ousAXWq
mPAI/Q8E4/VYGf2BZOzJrU0zO84SqlJk7FhdWxhuDN+l7qX4zKp3X3qIURNJUY2kcT0KkAwmYx8C
wrYBxtPnzNmXqhfLt12DM48aRu3rCN+HR7pWu339Qz3ptnGli4rP8+2QdDiyj60SDgycD8Q1nXJv
BUVoI4MWt6wdr9gzdc6aKK4PohigOiWhDn+s8jKqr+3aqexz7q51FIV1wUGKYwBL22m34plOVEtm
4zFonwuCiHItwR8Q4BRB1K929IDCBtulzKFEuOBrW0fH+uN/460+fFNcbxhb0xJTyCsqUqT4cTJH
N6qSYyFQaCX0s0Ca4r4+1zssn34cK2dFNa74G7uwXDGOb/MvpF4XiIC4lLKQLiN4OffJjP4BnmiA
kJpIlyoqbNW5p2Sa93FX7s+CGQWKfuJ5vJDQpksAbwURvjJwZbznWp5Cxt6F2dU3iyWmxJY5bT8h
g4Og2cxYB22D/A/skYPcUXavlSGZQR7yEJwCJwgsakvw9qkHPJLs5dOm+DUkxRYSIm02MEwvpZvO
oeo9UDCXW8vOHz8gQFf46bzUq4DHPpm9ow51ftlaK9hZQViAmZkzRKHrlMyGK53Di7VjPbwYgg77
iR2uM+9obVTJK6LPePkL61dLDRiMUqnQ4x8URs2lQH+BHTGFNvEgpk0QhJu2/L0xo/ZjsrzeGJnD
vIj/ETsgM/IpcEtUbz3cG1d4/1pipJCqobchzsAkfFQ6+LuSlr1rdS94h6amgMM62vcMBhJnufq+
GhWJKKcqO+lLv3q84Kno5JmP+/evtfBZr9MF4ciDBuyjBgMUmbbJ0pMhSvIWbeEK0FjzTp0jrCYu
bM87ZEWoKMy1xIs769UHQ5hSXRO6zVOs1bW686V6BTPSdHGYPaaJ9fAkvjM2t382JM65DxQIBCbj
32lCAKjN31ERBSSlvTS0HgPQGM2DFNZDoG74Qipx3F5aoVOdAvBca02lzyBcGkVAK5Gzng2yClPr
dopxVAv/HY26FN1k64RL6O7PQVOfY3XUWp/ECUDeLTdgeyC08FXiQ/DHREmi65RXP5g7q7H9PBYl
uAitWfcv4S4q1UwTG+cLFcLxegWCOgFlttNvGAR+RFov+vpiyko/2JoaLBKcyA2O9waB4JGK6fDN
C7x6VsnNV4Re8aBGDWj0u2gV9DDMgvU/Op87SLE0lIMfg5N/6fijHpP6ZgR0gT2E189SrZEK5fef
Z3e3le5toXOogKYpkLmdSVw6PXlmzPPwEiGyZjEmx8O5R4PlC3loSkkzHB4W/rZ6K9sHf3m41HdF
jvY1oRtUn2R5rHdNryz8GZ4bHb5Y5AD9doAsgDC7sgBcyh9IOCspBAy17HeDFdw1mCEZg70DDtvG
YQOiD4NyE/cg+Qi+WYArw/u6j/fpVeJM+RzmsSoOa5zWfIh8+9DhbIyL+u5DtF1chxXYSyJpR4vp
sKZjj96fZrKl4SlylCGZi6r0AEludRY4CwVxUI9/NNNmVaEERtbGRkN2vu8+x4x53qxrCAYBs98l
qXdrMpPBPQP1QA21JbOJXUIP9MMZtE3b+g8reg9j+krQjmpp1IjU9AJKoUiD/JREv/43brNWt17s
YmW085GGjxpcFoE4NT3XaG/EvvU/f73cX/wJkWQS4VKSS9Oq6XL/nB/z2YXh5HoGM64GuxwYkJ3J
fhDb3NH1C3EdUgML6TxXVkmhA5QLJI20zSykIOS4oXjzIRGlUo3rpauuoss54i2a1nxpmp3oHIOa
yXLovChnST9UiL+OGcHZtOcuSuuoEWihOaV41RVBbojgSIGxTl8804K/KC+bnJFpiYsTuTOC9ZaC
vGjrWCwSHme0adNniIMO0jzfiWCvu/zOesFlqXH3BWmngJzSjzWrAV85+OVrX5+4s7hLhRh1oB9T
y2v6AiYrPpLhhCWlB27aCSdjyJJnq+ZLsJXPlHduwquodA8yD4WGXmAe0ftB3zYFRyL1hjoCF+Lw
JVKfKoim+hgbQDbCTelNKERPKydQ97JU3wGCCs1J5vYz2c+F0xV8PfAa2g/pLYJiBbBX+fGtuIz8
84txTo3g6tgp/hr2xHR2OWHwUIiGkFBGH6oT/oZ1HdaD+fv262Nn8yp9KfhVfN0rbFSpQlk+GROv
iTs4SRpKYNZQXufMvgKFN/qSV80iRXgasfo9Cp8fglPzns4rmCoiNLDQP6o9NUf1oZfYw0A8RwVm
ClxiCX6OQCWc/c0k1RhTs7NLfgw4pLLHRaxUvKZ1lBFkks0mijDi2nDlrNqRjWHE/WEnYezK2OVV
Vyfk/WVvye2UMJ6InPvuo3zrYC+apVmZ56qbJhPqPWW/ijlVU7eyh3/3usRGUa6/4X8M0pyQ3EnV
2IOI0+rDD2+3Fg62tB8ken6A4qNJE0/ZU5AwU1JazbnbBUikdEMbj8JSmlA3KHcHKBzkxlo6kPfg
Tkg/ZHfLJnLVzkoEdKVyAVzPZbcls1hzmoeMj6r8mVR11CrUJ+byORB9Vj6VD4NJ3fGtuWW4Exu1
BOWlsyZYGvydrq0j9w5klFjNSq02MB7yYqKC0Y2sFyljhQXKi85kiVRKYjwlcG6OTH6Pf/RXChIB
7ZQBjhS7RraEk+aGUTwvaEMXji0DviVNT1tilfSGXqdUPAdyoDyyYOwH1+qJ6jqQ+38bzMmQkAQV
kS2bgkdbvA7l32saq4BREKOx6vX8JYc3l0pbyFN1OvY8rYYB+4fi9Il7/K9HrV+cpbDpWqkrzIBY
nIa7/n4OajJ74GR/8CTED4+1aQdjCK9OCvOtwhWyHIFTMjs/He/+1OZVJJG6oLxs7HBTq70FxsD9
1aY4In4z6i8la42DoQ2R60z5fnOujfFjO0eEn3lRqVonU7u4qM7aSH664CgNWeaF84rrjC/pa8g/
q3w5/wQUYNdbW2xkTnm8tWNzxJp/p2g/h1pqK7LQSLYCp4yHqSFZKXnZGYGkSC1JZH8S30zzOr27
yO0zN5xx50Btuiej6MEkccHgwt6s9WEPm25KIYhOZ6gEnq1kB9da9I1pR054p23m7t7TaYOLYkSR
onArYFd8v5vyLKRDtk1zuYTwMLpmw1C/69jybLSHnXeVczP1By1HfKNuUGKDzaBZmLLPowTzpYH2
be4zKZ+oxB3bLKq8dJ16EzFtk0Xt0CoPYYBniLf8sqg0iBE/EpR/c2sL1CBZFp1WI/TzQeSL06jB
lRH+lNd+cEMYD8hbpnobKbxnckBicy74mZaSgS+FQxCE2ssJy2Ug1fIryPM20WfSCab+r71ZpVOT
KW5ZOH8V3qwVPR6xT6hlU0dVe8rDgPTJA3rDHq7BelhcQVi9fYazTjSD+r8Z/0U0VSO3NpNMnoyV
g5LLMXEyiKAcmoPZr6I9hKqstGjgRwJimwalJqlWTnvBOLK/uE0Juu5driPjnzk9+Ki8+GoxLkt9
gEre1LKtq1hD5lwfmDzAfX0Clhiu+9nPRlB7tEPgH2YdDBiGLeIEq9kcd+t3SAqa0TKXZtJ7ZrnW
y7r1OwgORKTVq8s4EDaAjnGy4eFPd2eqAVoSNzQjHuWnCxNBFPQiQrVj0unLYI4cpFnFHWU13VGL
MLymgpoxobrxIqk/CVAsXc7DM9EPEcwgTFLXkNXZpe3OejAMhvQU2BFxFj9xF5XQq25S5SG6p1tx
4494Ca0ewIQp54nyAJJNjo7gbFl60XWC1DlqkfA3UAZNYcQx8Mg6bYqWr0o0VGUZy85/nDzaWO87
efYkhC4MrWhr1HIM9DAQ/PzCfrVyeecYcBStS016bjvthP2f1T80258aqrmoYMw6o1UHMzKXCWd+
O681wheRCU7L5vSzPEeId+TPVV8zKffJlNV+SKOB5hOR0ZfCpf8hR7GZ8LI3gK2An+vFkWErnpKW
gLXXX9+cieQ+Cqv+BsJx/sCZyFSaSCYvcAMx9mu4yLqHNg6TLDuP5zNPsTifvQjYOlCzNL1Eulmh
S3QV4M6m3Bvuc2IJXKrvHaW9B7JXMy+iM7PI9gUTLfMzzFhE+6/TJyVLMKBq9yGCv/9/b4mR8GhH
NAhnpwWd6jTVtNdgCxnOyVn9mbedOJHGbsiXCcoJ9m36JcYl8VdsWGmmuV5npoXa9DbL+bnicyV4
j8NxhgSDZHP7kkFYei+vZr86aF2Mk+6cpjjsL+8gCt47xdJMMf5VeDJpx5L7i5x9808uEFO62A4I
65mZy/24P5rt99jhwA4Wiefec580pwyEfhQp8slNajLlhZzCB8c4YLVuQLXKMkkC490t5m88Rapw
6z+ZNget8R1NC5FOkl3EA0ujqrcsUPqIL4Ipt8XKRErNjld0ivGpcsDpuJdETXHLHxqfNUv9F81s
RQrJk1rOLCb+1c7VZf9eLa4bJ8WlC+3aU+H+SNzIu+oJKSWnvJqUky7i3yegyVKZ0iX0LK8LHI46
4YQZ2ftuTVKzQtc+qVw2KO821I9IINrEd5TFcZVOquYYhgOkbBibH5D9G//69eNZrx6pbhbaLT3U
hUHfU/90beg1u1cVqQTGBC3t12n/Bhrku7Jmxg1dXZWp3+alO/uz+fmadDKzgow4Z17lBQt6s2Y6
A3JGisvxvDMhBWFkJ6mx1MFn8UDrK+HxhY6pvK6wM0Vid4r0BctxFGYTbE8LJdzv4tAzoXyEPrln
gF74p43MRSsUqGVD4ehVAYv/rUC3+EvkgJC9PucCZgzmJOiaNZp/bBH0pYE1ESQSd5RigSsE05yL
xDlcEYyOHPee8pAswP+mMKnu6rWkoNYuB9yTD9xRyuOaSv6mwNNZ0MCnuKCfM5/MKmWATGDm+5sy
k3GRTbYEK+xhN9g/ZRAuxHv7BJryqMxhrghkjUv1GO5s8Wub8aKHfmNCRdCypx+cFwaD/3fg+EKb
KIOZqna6XCzCvKGyiijsFKwrf8pODmWVXk+T+L4xlB+x7DUGKMI78j7XaESfDJiFhwjoa+waulig
xvCL6Qvhk9GCydcttFmy/eERlmDHcGjr46y9F0H0c75VqdJk7As5CAFLnKGDDaPA41DiT4qGDJcI
sa9ElMyqpUVEF4nSQCPgq7zUikoqwuZ11vJ6CFOQcvqQA0MKXRXaRsO7u1zyQ9QYcFFNe0A3+4dw
jZftTHUh2hAP3TtAKXBZ9ff/G+A72hSfXLGkfs4/BWzNEg+aWJmAGHGT4MSg15r0A5/27uNcCrci
AFd8o6FCVeVo9CBPEHcrxi5lN4xVKoDOGogKzHoE2ER8pxbHCdFlexYud5xfxxP8CXrSzN0Nx3Yi
3euITGjjZSGAS9zJval9Da/WKNJqo0Pyngqi0pb0r0Y3suSvFy0d7LtMoD0zr3PwJ31NrxbEYAF5
Mokpm06hfGWzBsypeqOryE9AGNDnPce4iRo9Da4dlpA8pUIgfOB/6NVlJ2wHVALukIbxR17hmQ/Y
v/vh15HEHaM68LkHWQ7FA9YjznwoQgeDHTSwsTY0CPo715WbG5wLOYW56LEOD6frpBTQamfogFdS
Tj+5XVUZPZBQdUT1zzoGdOPecgZtgJoudELbpkczAttlv8QYgtd0lyXyLTd3dwQTcz8NYZTO0C2O
Joi1CpFloGx/9oEbIinjSwS5h/Jj5uMpHZn3jcn5pjzYgX6DAYh8qDMz8KVW+TzS3mRJYfswaFRT
wQ5abuCLrrkDfyyt6y9iZOKLkCMWQv0w8aWXYkqI778Ru7ZNUExTbsvH6ayi+aNyjshAAmkL9epL
ZdyiW9EbdIxS0p2IcxlQLKQbuohDbg/8euo6BHP3zkBacyT94PYUb9L7eEJyi2VbUfnK5KZ4cBww
VYkg5RpMxDC3+sWxxkANvlf6lZOxj4twe15Y6qGhIBz+fKen5ml3JjqMTWpyX2OEe4R4L0njPj2K
wS8fykBK9aF2gZI6xZPG760+XAhx8RRMWrrFhHcqSqjqalvS/0CVidy6LdtVyTE4wnax1m7eF1Sg
RUDFT3Ey+7zbwXtgL8M2IiqLWAV+aH5RGuM+T4U3BnlzObd2dKAV7/Y4no5fl51BBVi88Vi9pnVi
e7IaUbdeQXOiq7rFYxOgs/K2p7xqz0C8jyhis4duRUC7iawz1wjPmm7mFM+0mJBRgKwUSYpC9gw/
XyOdZp+Ju0QAqFfo00oJSnmSP7si7CjDynAyc/ERdDJ4J1t1gLhs8gWUF69rpqxGA/qIRqBnWam+
O6bw2R4I9FLAp+a9zhfP231Lp4Saz40KncQsUb08t68pdpFFK3JDBxsqNCH1siqNK265eD7JKlD3
opLAVWYm8CwhRp5Hz9gvQIfe6q8IAxIXM354V6dsuoIJde6aTPZXibWo7/BHfEjffvd1xbqPclXn
Jd7FrGzOEJi7npksnPfspz1AmDnyzhU/vQKPn4EO6qxI4KGfX8VORHc341uZeiWrjeVqsMPtoUnv
96fZ9ADlOfo6vY1W7MtxyI/p6If9HrK0lbfAXet0Wagtemzw/cJU5qtHkq808Z2E0p7kFZWMcv/V
zvYAS1GjZeIGAGLkovfn/UxLzMuCJiiwz6CIljI6jBohrvqd4x0KYmLWcBNQZ6OXd4KWXlzUztrf
zezjmeTzfeFgxyKFs07txwUBavZ0gz7N4aGhi6PuGr0kcut/dvNdaysWEkrMjD/oU5wTdmXXGa+y
AGTyg04TYKsQFTBiTDvfrbuJjU+tR3jCYXJP2OSZvlXWDqEIgjXjBoEdTgCNKUz/bnaMETaaiH8F
mbKHcYvlXfvj1tun0mC+qk2Zq1LYGAgGOTwlae4XP1xTDMo5xtQoZ8fme78FLH4gMJAA3+AnbpKI
unG7MArwiDxD4sVOEvCP295V6RD5FREZmZvLNk+9nbKOitCPMbsRfTS5xmuLE1Afzb00uhyw0T8E
3j/ddudm5Oofu8DxAq6zbXj66uIhzmxvEucS2C9Ktf7LEqNwbZ/eKY/NZnNTRPqRySUFVNfwXKc3
jrH+vWEIbTGnVmLqms/rIL4R0w+5puzZ4/4GdG2256jLj/GJ65Ojyqg+cJ6mrcVXXgRpQ3pBtjQg
jogIgdGG8XQDIOqcHA7zz1WXQsKqXJKrZ1K6lCZgWNqasJbIEkZ4qXoyvrC7Hv13ahVBID+HqRvY
Zz6235c5/NKCq8GdqqxmCfNqx1WTyKN6UDtyaz8JnQSkXGZL9R6vdxL3MC8cjUeVF0A4xH43S71b
KgB/f1QWcAR8H72Pa5ZJUKxLTPGlIkwR/eQrw/PZIShOmmBNYHFr1bsB1UZTJnWCHlH4eq95CFD5
PzMkouyYzGtcqiEeJ8K3nSmtvpjcND6GvSMhe9sEGGmLY8xFltdKUX+awrYUjwk0qlnFsqsrGZPe
2okV4xOKATCVA8hSrZCPU6kPzIgVNyC11t71QNuzDxeiTHi49SVnNnNLC5NAQfpixFknGHmWj6Lo
deX7y2M0HlFMAVujXzd2WQILUPJlDVWrgyhYEe5PParYm13EUIaHiKqYVeBVW33WHCbiZboVBiG6
c8jlPsNGB3plLAiSdkRihZBNDGONoudlCh3DyAwWPrGYgNlW6V/4Q3ooQQL/hvRRgZZJrIGvw3mx
llA7cGVIhW7M2auv/eM6lpQFdCoiqpy5Trz+mQD6m/7UhwWp/FJIPQnepTrcT7bXOTYtKiu9LDPG
TPE/m1NMOxWw3cwSHbXV+2p/Lur50vgSVlnrW9hcLnqB2WAq8Vt7PHHdo/AqZJYGJjYuFYzzi58y
zKv3IWz0mkfwykxxHQK4H7NIalEGzcYW1orUtA2FQ4lW+S/m95Kv/cXozhAcFRxlkPpxCXreOQlJ
41ouPBYatQhYkEWQmrdox3N79StM2kRAOJ+mzxQbVUl7FSKeI9pAjGibGg2q4VY8ySSiYCC1L12a
xS8vsZD69ITOvNODCBc2qnxrgY25rfLgY/FvJfXxO2V2NMLPIA2YYf9NGoETczq1nzNT4t+hngxJ
FlV+0RY1K9lqgoTUqveJMkCzr5bjBaf79TCQLphhH7xoUF4DhbXJc/zbewKFz0vNORX/8hun6g1F
sJGFkqAOYL9BBYLV54i33PrdU6pBUAdyD6xTT/q+cwLbp0Yx7X2ObwenNQWJnAe9aYoP4jU4Aarr
PW+o24zqUlVIf8AMJcu/W40SL+389MWM6oYFoajscQYYbLmgrLDOFlFYTvM2QnZ7zCBhv3vuyVmp
SoUtwVN4CSeiwgi6VwCLiYApV3rRfNCQPUOQYBopwar9QRBfn3SBUNcYt7tAguEwE/3fb9ex31hR
UBV9RMw0vVBVld8fSqBPeb41s3Hsvjq8/6PXSkqyMNEhw/cMGECO8le4dCQ04NElDjDSyABIorMx
ZHc2K1O9JrV7MmFuhseVhjEscvPPqvs6aNRcbUQ52RAPpEunkk/2t3qjtWT84lboF+bJXsP3+DOU
ZB2CvGGXKm+yaR+Kt2wOg7ZnRHnWgYA/D1WZzY3lefRoqztqyaxBJNhdC7MBU84yuILoO4/QGl1/
qp+ktIJLHPBbuILlIIfFZgAoMoHgu/O7sgVRu3/0C1pUCQDwP3nLyKHJlI5FuKGd7dnCpVgpWpdb
6U515tdlJQaIONDp8F7nK7C35W+sX/XFRw4LPPLrL4NQQQwrrdByxaD3qdQeBeibN0B0tTqY7kDn
hCgYxb82ngYuTv3ikrC/Yflo44V3mRCBnHMC6qXhj01jh1NcQGcfgTH7EqKEaSPCUlIVl4Huycrq
5LdXgh07ICZxgSQkDOAHMToSkzu4oiLOKljsM52NvIv3CFdNMoXyWBDlgw+I/VSHCJlvxWq/Sxvw
rbsEoTqxbeh6o7sGedVRTl2gHmXEMLf5iCADw6lxPYByL6k3kgqsS8wreZZEd1a3776UnbXsSvlY
kQ1Zdsrqu0kKCdfE5I8XkJ3GN6SmYd/x8jOb8pm2muvpS7q8BypPUAixQX9OVc3Lgr7B8r/PSgmz
l1W0OGtWJkAsUyMhNlPXyps7TSxcrxPxHiDTHguEsI1LHhWiqlvqF3WQp3GZ6LWv+2qarU+h2vug
rFhATRKnVbmwnA9yTAHF6lQ0SuKTVA591ri8RBD/m+hMgG/OUaDeE+Fw1bhUsmwL3I1F5kU6/5Az
A0FQSM51aNgR7qEMUuNYqKj/byWrngfxPszhpmP+aR/Ae7NjSDNHYOlwjLtDE57/nAvimc3XPgi2
6Qs0I9kSSnUmZfIr41sQsRGjsXrh4hnujDnNmpTeoJk408OAlCXYxFUqgGHXbMUgW13KTqlb3bYk
KMyUFM+KwvDvWhEqFGfRFcAJwgPbGsGkpgZLaFHngjZ7xRMcb7DLGJCuA5kutIPsse5rsCU/dvyh
259udSdm808pWwjwDPY6a7CaelHGDNnsmDyfiAiWnjdKr9qztJKJUNE62S3YdP/Iu9gqRxZjTiqd
Orzzz3bZl1BnKCfoaogvfAAfU58DNQYTArR6/qJF2msTHTsUoapmTq/Qfsrt5wgHXhBlLW/SP54D
Oh6xz5R9UKJpMZPE0NMlC9xnx5gQRflqrV2gwerRyBb03jLl4REQ+CT0jJ3hDCWz/hxGx8xf1lV3
WPiH7vtF2JDPcxLjF70bWE/NWeoiZRrO5NRBFHkEmUS1DLlMDvWcaZBDdD711f8EoTaCaQcy5tdx
cjTuAEm++Wq5tcCOXOtwK1TamrqPe1lCgu5GMd3pz+HxOuTbTCGhuRlkwF8L7QcjfPab6nC5Q2FQ
vJG0j2oFYdJyW9lV2xKd5ih+Biby6QBihbE69dpS39nh1QUEDxFonFX3cMVtoIPQnY4I4JTBIcAx
kbY8bBeWbmuymQVSigopFVHUsCp2X5Etk/RjdYA2gcOd4mwxDQ58LP/fKUfC3GzDz/6S+9PDLcjs
S69+bQTyMrtqGwiKOSoEBZtcy40mxxIy/JFCIXtO2SPRCUr3P/zQYcspROf/e1x2SYi2MHfgmzOL
Z3dSUwNk8bdunf88cTDwMe+Gl6jSGLZnAKjnXYN0QckSuN1d62bAjmjxyrfCdpsNBkoCzYoE5TSW
GyLtVq8j/me0mIVVwmcOpb2f5kFljCvPjHEJN7essuHr1HdibNWLBpnLkvl9+6aLhC26430vPjv2
azVkfrLDTCmuYmX3LRe8BaJS/S4DpSfSaILMu6dqwi70MyMgW8U9XbZcbxD/wYWdG37jFOb4mHmJ
VJNRmiBUi+HjL7TmeVKvBhOyYZcUnoP6NtCZ7myJLthP4oiuZRjGncI0vKg2Kd/US4upZRBSCdYH
hVKgM35aGs0IMnpqJoZM6jaYQxuThT9306ODelD3oB7mRUY+A4/QXz9SGAagZ9SUKa8OMH4N5+K3
NCiW+ZJBlkF72O7SYROYEBHGIXUc2XL/8yTLN5ysVfTG3Z0eSzqCXWLFerrU3abXm2nROvlKnkFW
FZlDKYZVyQb0APoBUQwI9vWTdj7H16OjGybFkJSpQDFHEQZEvLWkxcYkluxZ3VhfjwwXCoDSn9ZB
frufYky33iXx8+9ZG4wKe5cLBk7Lxxq5znRuuS/iqx800QVPyAzqfvJ2FxVswX06l4sHC1apgomy
bBb8sr38FtcV0P8IxPqOgsWUqcM8pCjduWfqQKJZbna+SUzxoJqEk7WZJrAh6SuMqwTD/CYe6N9A
2QlCG7E15SAEWr1lATPsdwvrzRo47tgCMIlAeLki6pCM2Frt0nIGd3RMLH49Y6+wWUbIqepRVvVc
yLAaDGaaOX1uTQCd5qdGgqNWbifKGhjwKB0BHFZGFx9VT/uqJfmUbrE0eSC1J88fsDDd35ZvKuh0
J9HIk8IJ0CaI8QQBW/jTB6iG4KRB2dSMveYDLZRvih35CbK/HXv1VNQxN0KBVrIiwWmn8kDVdQZ+
0RIaQkOL9815U1CSqORForfVudvGcbzKCsNR4sJNJSJ/Pnc7TZfHzqS9N1h+HdGz1X0d/+xFAGVe
64KckG8UY39IyeKWJ0d1ZKt59BYFKxSQW9ZGQoYG+eEk/UM0j2vT3+NNjqr3t2gXSuEgTMAj5hNx
BJoeBdSHbm4jJwejUpbJxI4hRHLgXkB5JAcrMtMin977cxu6abvMf2ROfUIO3p0K5K35c2XkeSkO
bGuguBhbPiX8+pY8Dj6Rseh6Cfo1KyjFefNYSdt9qTmqMslSsnN/eeYUngGu+ZrD4bGnvd+aGJgI
Jr78oERKNJjpnDGon5dK5qUdL6rFkHhqUOKDJtg4KuIgv6tsUr5Dp2sCwJAAggKJPqfLYE4vWhZQ
Li0LM+lg5f48OK/VekBvSezlAcuLRzPeyEYplMFPQtpJHaihqKgvNs7SP84+HsiCmP31NE9gKlyH
gVCg5T7ZGxZNrIex4Lzrs3I52027jhxJmR4/uQpeddLb01Ri43jA64cvtLcbrzYodSpV/kFDVYeV
H1a/TY74Y2ka9brSaYwvLKUSp0JC7dPtJXpEMqoaESZvHBHe6wa6r4yxqLsIYuokvn2lSLnFt+IJ
zcWl2yLXqNLM0d3IEqj8kkvr/VU/iQdyB8i/zUNAqM0hYv4snxQDIw7Qr86IA33IM24HJj8bOnby
L+1lJdck3KOMRn8FE17mzEUigUmGOLqlhIems2q8rs55nrpT74azeAhEybiEK06EfFR1gyI7w2Ow
+qF5jiGyDoZqsSJaNq3+0siXUKVWab4KIfVKbHzygLcWItmnrhxCny5H+6ko/wAtWDmWaxm5vDkn
tZLpfpMxi2IFU+nAtUq7fivdU4tC9l5WlHU+ksI72imbZRUGOsI9lGGbBOmXCXkc9qSlSz8/ucqY
wJRrtcRcKkaqLqWgQ6h62ro3VojE+mdNp7jQVbkRhBWyIZJ5afBAqTB0ZZMpmb0PWOg/Rd1AXj/u
Bm08PX1aNcj8SoZl6pIpn636qazX0MNOffYQ23/h/AunFyS+ffml+2MtWKVJgn6EW5h0PO+aXGxZ
vJEANgi4rkv+8GWnDkfRQ2oqJfLOH4eFIMCUfVSHwNmbYmWOnR1mxD06Zp9gO2eW0fBzKCpcQ9Vo
tZXEbeR1E81wljZ/6MB9p3QHog7jfuzKJ9jlW1euJBnRtTlrsznnl4eMTlBKjtWZ3y/Im8X5ANjn
P3wv/WiXf9ISbypnqQzHToIT0AtqOWlOnfvXjAlvqwPLPmTK4JrHYr4HrERxdIukEFg89JUhVBKn
Re+QGLwkrvzFvmllYmIQ9L1Fz+1DJPS+794D9MHYjdPtwljR6cbjmYKxgFIhuVT0NL1UPHkyaFkx
Nxg7nCQz+bJLmeUNNYCxJbiuVnAMzAQTgRx52+fyQWU7nwA8xqHkizUtNGYeN/ZnKTC+4ef16kn0
C0GNwAupMkwa6kVk0imdkwgl6kEEK5OTO7J187DKPeHcEo4zagx5hE6qSSpOfQr2z2sQ6Orq9rzO
ybWcSMPug14Vr+mDydHS7e0MXVqyfMQIfvLOMJQG+/YFAQ8XMxKkNjgdLNavQMgORZnlUdDL7WKY
jc+U//jIwuL6pReTpXR/EzQw2gW9jj+T8po9xGVmoveJGmpVUbEJbZf5E62xags44nViYtKM27f0
nWrfGr/8Sslrfc90R+Pqm+bMSshHaY4ydDIvAVlcQ9DYPZe5ob4Ao/uV2faqpZ+LSdaRECDyX1xg
uuecg0T7H423U5IzmEblI6b6juAEWAJ+HCWaFnfKof8Jb5rz6M3WhQTeFuhSPxhXLAyyJdV0lVfo
khdRPhUfWfz1zCYtrznARL4MRRok67G6ezuekEI3B4ecbzOEmeGrOaCsrc8Exfye/InY0EAo688j
KTkDQTv+i4CJWTvovgk6F61QPF4mWTbRvNEAgy46Y9xXZWUmjI52zQA/MNaC31UF2fk1oZHkPOIl
E9YPc0Grv6aNx5UlsMjkPAJSriVBdXwmX6pokBTND97PnhrWlpNsC+rOAbEg1cFqPwHiqeBiu/Iu
6xC8ZqKbkaukvVQq4Z2EriNQM1tWNAhYsr6OnWycaCdS/7X22CQnN+i3BQ7a/9SiIStAoeiwaKiV
Kb+u7WAxJGJDp7ZyHtuGeZBP0zY021vmRdJni2R3rpbVFcowfM9ETwOts6sdB+HA8ih3D+MqyOvS
bFpWoj8lsRqc77oovqGhfUNH7h+KPIwgV8NPh43sbBBrr2o3pTTyWxgJtfhRCoEdPH7/ARFVs1M2
VxhkC74xXkDPEFAyTsuTJfpZEYiO1k1tGQ4AUn/qOKBXlErhWD908Wbwcd1wWgaCnU9ZuhCYYiUH
RosHT6ZY/0JJWE3zQikR6YL5EdPWfARBRITrWf3RHsKUQliAuhFOUKaSrz/SInbwY2cTkh+IfgB1
BgDxz0zR+ExC+mcJuccYUMCX7rbBZD5Xlo0DN9HVtHLr+pFqNzYJ9powslWgYjLESRNmPzB0RCvY
njsRvTMR+8/+0o5kw7yWWNT8bC8tldVG5elQPy+1PQBwwLtOy/LGbZJI2rsG3pq04L77hY3c/UnP
gCRF0ih8dOQ3ECYMIrPNnb13QGaXhfXgO4TNs0g4qLpn66Ea6pxyvftNsUXyIIWZtjbBcX9bQZM2
bYEgYMvXVqNqvUQymE69SpzDOJTJ9Qi0TZ3W7YwXLrmd0WXGVf35QOHvDiplGmUP+3ILIi3nB1R5
VS2ABhsH4E3QMZZoEOD6MaWRCNKwCYH0CzTcaDvYi99Zu0Ya3GYUDUVTz2XzX4sdF4eXEiPi3J7g
vq1wIvtbRKB+XhvE7eZuY0Ln82OvHqEWoMhOQZ/SegG3jncTEc/7AbAULjxXomDe/t1w0nqIoeUb
R02u0ZFIijfrTQXiBcX9m23rKHVFKOemREcwjRJaIuUifLbAGnZX0AeSYHflV/Nqd5dXnjWL87XP
RyDU1sA9oHtqYFCXs3uiqE7natOSMRjc0AH8KYBvpKUGikIEerrBIZksZHgnNJihhaDHz1k9Aj9s
EdHxeXPyiEfkCD6dFtHsHC+iqTbcpw/22lXvd90tb9qIQXth9ofXp9DoT5SoljbWA1pKp27zeo5i
ODQ2L/x6e8fl22lv5igPXPOUc93CmyTbEI/qz0Kmu9v4dgp9pVTBh7x0lJrVOlZjyJXhCril6Cq6
SoA4yAunBIgwjt4lXOC0+IUJsOLwPYO86QZ3Uvx9bTAs5A0OwQ2KXbQM0xuPH0xYo0a/rztNZS6W
36x+t8pjgom8+c/7zkB8xFEMHQAhrozOozA28JZRzzuVlYadLJfMPmKwfG8FfRmgl+Zgt/Jiy6Kj
9LW/C7ZWN5UqyKUv6zn1eflJWk/cIBz/Mf3eZLk/v6Lo4KW/CRIsm5XevUILCB8NIhTxw9FO6ogc
TkSgeDE43B3sWIWwbDfAXL0PctSXHiY008QK8Ke8E1+NWo8cS0Nnj/7bM8kLk91hCGyA7p4alGtW
mDTvRadiNCFaTumHCJsXs1iDVnA63faLaxUOZFYiEYS3QknamhsxbHAz+KXbQ2QfWljOkHUohwmr
mdWIAt19EA3B/PH8XMNa4jKl4LdqfC/932PYQxkWhbJn7/eLrCiOQin2V6AKSuXkKDRQ0hd4bs+9
OYJV/7LhXw1m9TC5yYKtFUQvc1uxxTRVcfk/Rl8KS89RADCppEe4Al1RW1SD34rTF0EYXb5tGpK4
Rz7/zhmDM0tzerezB/HxQ8mcQr8Kp8ZMDMC2HSnigucAU8RDvMSqEcQ6FUT85OdPRrwrIDr6HCG4
iR1GzPhvG1mvhErzGlw8GLnmNPzZpS0S9SOAEFZ9YEWKqDhie0rxze02UNG4vI4TBQTX6QmwUSa/
mzHy0EmR2YM+xdBNwAUVst0IUMVwoTDi08tT7jqtJ4tfpSUdsv4gEca9iSwVxc84jyFxmePaPZJL
sHzYwv+VWTjYLNpJ8ZOAebNxwPlsrtqQlKyxIEPY+Yjz3v6cQm8VwFh8Ac8mOt65YL3lX63m75HN
maf9nHJuIlumtqytoZ/w0+unQmRsTXldR0rZiEwUn8LfBT8yDZpo9gg9uLgxStnYGNasom0SdBRl
geIaV6OsBZe2xwN18z0IwEC3+/gXx7plmZmgPbVBj7kqGt4ceI95/mb6B71qHobauqe1df340DPc
3t+0BavziCQLULGRieR0wBf96GDG1Fa+bAhyiv1Mz3VWiHbDFNJiDtHuWBD2rFJ8RzqJeJPu1xa2
Vig/LRvlJczR3/7hOa1n9TPvhv9uLaOSD7yIVlnaPxnkb2Eyzk7P86nj+NW3bVFz49SU+ifUoXBn
eZeaElwdaeuYU35Um1QEKuGK+hWuvyiNk2mRhrP/5r2EV5A4LYfMZVmxevd0/vtou64Y0IsY9WJP
fjzKFpVADybAWg1DXGenkaOb2J9f9hfenRrmEEW3GVXmDsqHz/Vz7DrgJ0vQbicdZauFVczUR/o5
MbxxPyMy4Ln05jcecMCScAL5NJVvalEtjT7M7LcOFksAS7liMq9xxXnfN0TmG1dJ7oz/ORFCKaFX
SQtvQn8OWlADGGSTjmOTNdsyQgtc97CPQYI4TlHct1iteq+7ChOxJ27NDEK5iACGMxJ3CW0ulH+S
CkLtricN6J+6u2vp2K1NPbelPRI7sAcT6CTihHB5HGJLTbRCTTfUzB2bs/5X058IFGQA4XQyyhMZ
S93f2ZGmyBMCD+WCH0E/94VQzw8RV++PRZ3juZH+bWXPUWNtlXxjfOfH1bBowPz0Y7fSoHOkkSGJ
l0MmQk5JwA5mWPhpTCwA7/izjGfl/T8vz8ii51tKSakwLuqSKqelWAISL8LB/gnvn+ioqWRwg8Qr
VvxiHdrtgZ1JLN6y3S3gs1iMMVnzl02Oq6+OMMHzklK8K766L5WvsE33FLusDFsyRjAT75FdoJNb
AonGQ65YTBCki6EOw5g4jkhT7qzObSBG7l3r4ph+BjtrLP7JeQ6qYovMu771SNIbaKN79sohq2tC
VQIA+U5SMe7DVeptTiXne2AK8XfpLxjSZUVSLn0Bc6+dBv0tKVZIyvexBCSlKcAnWxDGUHwuKieB
BNIKRaSa7ch1UVfY7tEZan1MVU5umobySbZMxw2TdkGdJl84JT7tsEm5s/Gh8qzMN8Ss8joS7e78
/0Z1E4yKuXRbFz0LPLMFHCorXzamKiZ/Qp3Yo4VOnWE5QJBkKqn/CV5kJL79zB4Me+6ytoTJgULX
hf3Ny67gD8rg8i1Tj9bLdkw6DYfaJz60/W/L21BkWVQp3rm9LDsdzUnDQuLQ5RpBVUtfjFQz+1GB
gssNMdF/n7kPQ0plsRGAiva43QKABwib6CHDkYTSGdB5RN7FqwwoPKYfidgCLd+9L+ut2Ih4/hFc
PPwtxlGpb4n0fi+XnaRlktUJOSIAEAmUvWbnHZwq/2R/R6MDCct4L7zmcl+mP6z3dxgyRS03Mcn8
on6tH/3JlkwjsltWc36dwFDlA8KqQe2S3RlIVDwabpBnBugGN/qbT64kWZqy5kqvNBeOV/KlslQf
wf6ssXcLy4PuYIta1Fh9Ag85iz/9KKy62yF6nzYWNDs+eR2U1oG/N2kBbkCdxuzJFJ7N4TXram1r
Qqlw+82D4Gi3FhIbSfN1liVU8lyVQJknUWuXjg2es8tEdHXp5qp6PLTUOmlJucjI/kx/scmfTwgy
OrxlMvxWFjYmhSwODjccU5QGlw2RO5vGti0e0xEIBLLDbvf2hCv8c2Ow/6ThwsNCwWjYtrXImvNi
VZBKrqtviTSXxGXKK0YX0Y6DIrrniohZ5XHRugwP6o3vbTx37v5BCI1VdbeY4CsqI7qgIXdIb80F
WDv5M/ZlpRQRX8UnIw9Tt7z8e72wWT1s1h0MX4tqPUXcFIlZbVzOPqFSyqDXHdZ7uTRx+7sK2O7A
I+rAm8HviPPeLFgtFmEHL5smAIjbENscniqY9+HlBpB80nFML2OhdjTpJz0e4ha64Kiq5BOFybfL
zc4QT9LtO1Ec9bFgkwDfV3xKpj2AwmAa0UrptCsMAZ/hQB+3OjPv8wDZVi7WlByeSKyc01Xp4+8x
xKO1RQG9I3vnzpO3jdH98UWObZTUwIKjSEl52gvkUvY2nLWJJoN/pll8fDrKz6kzawAYZ6C/Lt1s
cWO6kk3XfOnlWfgQnrEOjyo25Iw2tKuaXbn0EsCQPNQbZDiw8YEin1jFpme4JyMG5wWUuhcBQpih
oRNuxy6CPO4eM7hdnX8/+CgCEmnw7BSLmI1uTWnOgzhAJW3zimBlM2Czn6tqLg5671o41pWfmGIu
iLtC5YMqOrfuo808prWa9fFbXM5y0i7iiKGe3hQq9l7w8SKodXgZdFqBgfIDCUjL3h7fKfx3kM9c
Xx85YQHyJcANk+EwYQu06FQyTADr9AMUkBuNN/4e3ppBOX3NCHRrenuDa7g1vPtP5ewrkimdQKDf
00NtQq5woPT57MkM3XKBEko8GnkhfbIv6TLxs/WNuodGinUctjWZqjD6yUV93uWjmSnPzv41Q9mW
IVqTrGfizs2gTXD36pOWLnHE+l3Vfx1osGSk/fXdv7ibXBc8nHw54gRO1IOj/l5HqgPvAXR6k5Zm
o3325QYP3ELJCFzXknlAc2d1Ooyrk4CQMR69H1oQLHq9G12OBmvUsdHeAje/UQ8zeX2H535mIoM3
Eb5BaifevlL5c7PtckPPK8DrhGVAabfKqE+KaAD5fwA8MJgRp//BR7bjSQo8B4eH8h5wja9fkIo9
OnFE+/RonTdNPU/UOw7fxIFow/s9MpklCKhAeXzYsZ1BEvH6q+JSMwF6O6IboLMsQp9hJnao5xZ0
hhmOzLajgSJ6SKbOpeMeFZ/bRqDb1mwp64eIOGiRT7zbu6oVhFtlzORFgu+gGzBLde4oMPhaRIzI
pL4DoKRMYrjzErZlSUau6q5U85NjsMvToyp/HqyjCfmLmYr28x1gGFQW9vA9sWn5RdnQzl3VFbjg
bd5tCexuxx/ejdE4RHGxuniATPSGU8TftuhsTQnQd51JlQiTH6vl8Igt8mihvXgBR0btnj/TK2zO
+2pUT7GTXbFQwoqbdhXWA944tgpSpNCeSjmkqKfhHhmX2eyH9lslr+W9aXHxG7/5K5qy7asslvm9
0i0whg4jBYyCPG/RJsAS68kTO93efhUVWVoGaVEDYUqpZSXkai0TmZFnRkx7f95KDYhPCddkTShL
+XdBlV2pfSWgTYSFuLSZR7+Y1vOmKDERl1/prhXMIEEj8pQvQcBtQqyGRPybcLihDJFvAdjrlILu
KlTtLnOuqS8HmeJFLFo5I0JWnNkzVyTcsKlylzT6t2jm6TW2KWGstrZ4ZlatERMxJaSW8OFL06Se
NJgBOZf0p1mxCaRXRvJ7Gczv8N78WYZWovUaQrva9EmDDdEZwt56MyjyHlUEWMIAjGxk2Y9bvxAn
/OW5tiHZ66NfjN0sIAlDHDRSCBdhIlBG5ksPsgEMOi0lGnIlim9xeKCgjq2YJVQxjlFiavNS+dTp
REQoMVRTBRu2+rIXARWCkd4try+iqIGpRzsp0dcmF4CiEx7AaX9ZgL3XBzpQroCXIP8i/2ai++pf
/f4tmMlVSuWTCAgyq6B4kncbENFpa86Q+8EO5+C850NmndyylCbTy7Kit1YjXw6j7oSimniT4Qw/
jBDqF75yU8pM+Kjdv5tpSk58E0lgl4jtr+b5QldnxzUvEEQEZGPLoCzFxIDCJMe9b6NHSqbuPx/0
4qBOu+dfZnSjAqGIjkiDHwQw5YGB8sA2qzMwi+yVx+VOxi6jk/tMkYJ2XJoXi8nJxGH3Ija73/g7
diI0UYEZKNcc4bpEjiJyKgDYh0wB8Ft+tSLzKQcU9FiaNP7OnhXBTVTeOzmn4TSY2PMQaPXkA4QG
1fs2yW/ASZ3w7bqJBJBJliAkl27Zda4v5pS4ERFnHiyl0BRAezS8SDAV8cQYB3umm0PSj0uHs6N3
AL8V18FRHxleIe8KTKYwxWwSsL+gRGpgALGuDyRxDJX5s84/rmqGeoCgelD8N/7fb6RKd3sTmnQ3
6erJ0P0XhZJGHGRsiZgDpnB5zAp1hoRnAeLzjDI+IFHzotttj+Bgwv7vOLGJ1lnCc5OA5nKmKsGx
LhUyBZwRupFKOgLttZbezY3uUgXUmfVHTfn9EaROjB2Bv+PRCwcqJGXZEFqGKroC6eWadEavf8Va
C2Ppy/wSZiLZREioo3TCOm375AU2cYvKrvBDW7PmemU6++6uG55rLf6n2CQneuOykx87j6YGKZl/
XzZMZpoI9t1/YSvJHt90i3/Kg64AjsMIshSnt7YLTXbzdgi0uA+qO7BE/i5s2T9FpVrIxR43/hk+
UBunFCtvgFuqZ6rkmbOy1x9etHlTWmOKmaMJfq/LFQ4lgo9XWv37IMyyjpSYRP4sOJNPtAT/8rRp
fr4K3XfVNwb8Ued978YjWiQcYRVeTTulJBAP8rXNaMi/PSe7XBgu9y3VcSUozyFKutDAIWvXnrQR
F1IIwow3Jg9AoMerw7X4xPyUOTHJJPgMKrdZb3BfNTJQWHeF/Fwuy4qbXlqp1mG1kLBKGg095l+C
E6zcaXKoh4b8dGQuNPmq5XnVmJwMdPAlSFM9BrD86TMLEpC7EIh2TP08O4q/xf/AqoErrBzC5F1X
CHLmJaoRkJjXOeZlWf8hdTVvRvp9wiKvm/teXlxtUJaFB87+YLP8RUsZ9MrXdNnw336ExlwExWFI
zLo2geFtCpVJ22VgqazeGvwqpRVH8weZqZUX/U1WwHXVSI8LVkNk64OeCbNZJygKUJtoW1xqB62c
cUauvWobuABMFGfSeOxarE0w8H5zbYSbymxR00/e9wU6MyhuSv3Nu41w8WWh6ClmTtA9/Okja1fE
4kWgIBgP+6XhRXiR2e9qAkvxefsQouR83bed3d6eRlWWcfJOIm+3Zz9p9IqsDX1oZfVY8seUqQab
7b6N3ntq2dR3Q29nKssnRLiJyOHOUq8j6HnMWS3+39uCkEUIi6LiX6xEH+9JOBzYehKrVZhAqjXn
tPET5c+2IgGVUluEM1xFp+4EmxX4WwY7exOWhkqb5nBa63TTyoIWAs+DP2jJxLvDp0mmmylJ0qZA
mGNgN94uG9Cvee5fTfMc5cxL2qdW11p4G7jzKtPWSWxCYDgyL8e4mMwgMwxWobJxQbDE7gCQShNa
7IVWKlK7nEAuivj9FhCbD/w6v+4AnXZJutgU6pkEBgKel+jX4AsTavmV6XR1IBXmJlP76GrqvWgj
gCunZ03HsgA1zA97Hdsy/gPbsaj+lbWuDgfTPCZV+JkxCEI64oGNMT+KRw29JqJC14eXDMwcx7/T
KZc7/KSTyzilGIIlU5yhaId2ItDhRS+WJb7DC5KM42hjVU5IXwXdKWiejazjv1c4kJBQF+oYaGa1
tLJXAUhG8R3lNCBRopAac61XaGD/rJTw9taNFteauZ/7qa5E81FDxd9hf0w3TfZxMwTVKH73XiyH
krZHEGEPoWBVPLsCPCliJOQObdzSme0zDMO1qGS0LIe0Pd8vdGThL0cSPwXlc7cHiE9jehmaATFh
49UT7q3k2cJp6x6hxkZ8aN28VDxLu+W2QYaBxC+QmjoWRAa9/q4Y/OoXObUGbImVYqOl8P5hUSn1
jWGNq/Sc56dqK85lTdcEy5BNLFnxkuoly5VQFVvfp0jPmoqhp9r4WNa91rCmz5mmQgJskCt7zmK/
rSIcAWYGeMT8MGbAT/J2nvrXRwTjwlR6MhfFNafsnS5uWjo92fC/rSIfzfzUtaCpt05RyM9IOvIk
ut36hAZZvenUaHGGR0LE8TKow6M2uudRdWTPRN2xXAV5p4iGbfaFsG5US7pYqg83ubTCMhR5YBsi
RQl+WezLe/8etCo5Y0O5ctoeUpTHDpHO+qaFcijWGc2QFGmsIYMyGUX0r/plAQzKMBuYEbsXTREg
m20S7PtDSt+WL9kpAiejaYsYSQ4oeMWtKKjFRKLMGIBkZPpDxJfqZ+MxAa2nYl/WyHqG3NGgE+5G
LSYjO35r/KcMJK5PrdvAS1u8woCjOK/nFZKlDK69AqCgr28BI4xe+9nXy771FZsqDuCN1/l4qcUu
r6+5gQIrDveifcTtYTXszkKJr2MA7oU11uNfK4/rjU1MBqSfuto4ppCbZK9tFR+XK2KzifCe4nKM
+coYwzS8FIfqQPQCJvFth/A1P/8KIijD41EmEAtMuevy/1Yg5KDm27NELEYo8FIO+a+AoUcYjKP6
IdeuEb40tniO7RdlkFdfJZzzsudGv/6nfsI0wdWQXiVQaWRnd9PkXX3mRkbd4vcaD+BEdrzOC9+/
WlYuA4Dw3nqPZ4LcrJdNDSRuC5N23dCkJ0IXoPFDMXZ5Jk/H8y7ruuPMVKI7DXuSbLDoVok94P88
u2R03iQ1WqjoUk65II683ToUZEB6oruaXmYfTOMHUqP9+2nEH7u0s2kTAUmHZzzPkBVXkI1s3KIT
ol619DoWYNpSwZ4kvG+Ez1iFF8rrRODsYzbVTZzsvSHmG785y86KEsKA3FH9Jr0UcLq+zc1D8n5O
vri9xpaADXjuWkJ1EEnfWWam74oA+6j0JIXwYYSryQKd2sP7CV3060uNrwv3C+KQlyJvHtZHQ5H8
Ilif+scpcm2cVj51P7nOgwIYAO7PFAtbjo4ZI2w9qLKVWfgiLmQ8HRxxGJ6j+m/HD387NUjbY3+1
6BLcmK0vMDlWZMUJrXruAmzW5rDOhnkZzlmbGVbKPUaAswW5ub3lu+XrCUjMjibEOxBE0M0pmsHB
NcCNI8IrHrZtaMDLAxjkCVJqJxPuzj13PT+GDLFsSIDPfJWDDUk1uFKOEIm4AQdbzLKcpZY6svvm
ZJZ0l0poH+UbffXK/SvfKFnU+sOrcnTM2/FV1oA9GThaXrtnitQPGYUCvgopPzweOtTuYP5dnKEN
r10l5cZH2gcP0FeW7zToU++a4s0bF07/szW83QM26Nv0RvYsuexTwT2SLA1CFKISbGhifzBizL2x
5Tk/1yBcf53ZiWjcEf4ln3yzmJ7deRCKvgeXRQAeTdBWPrapLm9dKIHGiJjQ5VrwJys3Z0Vk5lKA
YHKTYhvolygWK31+q+O8UASjWIKqIuo9uH67U21Rukc3Z2ge33szcpANDJLY/mxqZWGuo5ru+Sio
fErwkAPaqlcLqCtRAu4v+dXjDGoXn2YI6QrankxWQb32C2cDU6R9UVbPLhbOCpodT0fAcqRUnZGM
PkHzGC43GNBa/RaEFxLb5l93ZAhAQjQxHTMqCM8oJ91AQHBbSmXY6BMzrkic9QirIX1QgiqvqveR
9mNAGZ2xsCeZj151SI6NoFlJAjE4uyoIMoev9mdd/5t4lMR7SaUQxfvGBYx2ZXRn+qWBI6V3UB5Y
a8i0rbJsGHr0drcMze+LQODPxm8N54vVng8r1rAVb6/+WcHFb3TnxT2Eq0WB510JWscAA8UUtfOA
45BorE5fd8+OWRACeBMVgXAIE3nghrGzuhrnWgqAznK8wjdnby6vUbspxjQuRzzoQh8kP7G/YaeX
57iWVHicYfaYf9DSJESKlw73E5z79zdrEQb7IPOBNe2hpvBdY0vH6lDSGkVWf6IvF9EkSeuDqZwA
Xuxrw/YfmwCAc4dKDOC4EojjUbh/r4w02paIm4RkjX0J/Qo91dK/xZPXzMU8mFOcBTplle4+Q+Ad
0/WSjY8AUkWIPgOQ1QGC6qgOk+LK+9zuwTjPZWPt1b5OmBn2tGAOqqIH0nL7nQwFiVNLYrxBTx2p
hB/L2dY3WROhHsNQfFVt6ohmPvsI2sMFkgsrCrhYKT0M6+v9RNDjzGSsvWVmjiU+ZJpjU6wZbWQ/
kivYjafP+fbjWFQJyIqkkAqYaMU/FejkBvzjEnYR9RWlT82ny7gDLsZt/F19lXvm+ME8JtHd2Dev
+YPDgIWqrLZFC90Ha6MYgOFpDhRNeiEA4U7wcVpGs4YSCG1VkSChOxI6ZTgKIZpT6lsMzVe+0T1N
1SYQxcpX35/u9RgHmTi0CUUixOOS4QEDe2RcBGRv9gjlUuiGxYYgfrUz0lJVvTg+xLGZmzvybFf9
pEfsW8BvR040OpIDl0ENuObCg3RaXUY56BPwn0oSwXmBm+7OnwKTtP4kQNvEPXJFvo1RlMm3OK/G
LHX+FpREjqd0Dd+0sPYkFO2ua6T0URzJM/FN7ZzfGStPikTcf+04J05kCBKVYM3koDW5PApGtOUS
XDpeDdyGTI6c6oCx+fd6Zu6Z0m5nN2K338aCOcHVWxG6kSwcHuLBybOyvrj5BuGoQBdEbEz18DAH
9bD0Hfg4OR23Re4jQCiYEp0ATTPav6AMU/zsk1Ay40TOWEVVd5qkSPvfXvgdAbmsTpoh76gcQyoG
AN/bBr+EqIpN20RdfPGxtR3ql0zvV/aYPRKcJi8jAixsnydRTJlcZygwXeBkIBkBE7ntUKe94jFS
kxZNosntu2f+1BzZZVYTeMSOcWgkyitERiZt2chO3PYcaut5Q8XfhFbrs09TsgmqOqEz1hrtviu5
adxU/3UCpwbXdfy/xFGsaoPx8qd7olX36G89viYMX8QiRHVTjctngnZCEbVFr7MLh5Ok55YEOF48
J97bS/nLeHvnx0nomtlLsV7NhSt+RCOW6OdmnMSgyR/Xqjqmy4XVk6as2xM1uyfu1ZpVu0W0nIZz
LzysbOTCxVPlQfzNHZht6ClUhebCUR1fPv0CHmD85/86yd2v9S0j2EhggXJmNTVT86a1FUlgQmdi
piO31NnH4zlgMaGHR+ZFHsZn/hoRZZGsUhbrCozxcEkBrxCF+1IiOWhA5j5tJPgBzjCuZsI3/qwA
nbomnY2Ds96WqXzHOW7/qk+XiAaKa51FcsscPUmnLoDqBnGkNi7pOGm2eBNIpsTjoFzTW6aRl2z3
rF44obS+ac/n1VMNNwQ1pOuu9g6eEF5gNskU70qO3gldv9txl+2jA76mGkCgucJ/4WRq4NW0OrZt
iTSJvP/GMXabO/or9BCCVSPut7THuBgvZ4SOoXrOWfRQqi6P4zfYFP4dWEGSVqzVIxJrPH0Bq56u
TlD+fnGWI4EXJAh089W1Kus8KysrvXFOU55uoRR7Rul3jHkU7zjkSUwuIPqubQWUoOu6bI5Do5lC
QCH+Edp5Z61gcO3JSig0aZABFIi5E6fPL3CJDpGTboROnD23b6ltrKmvbybiHXrft5dAZ7CdzheL
YJgSws/bg3Cwoe7Z3W3cAimrY+6Biq+DtD6jcG4AN/a3gycTkpLOEeLPv5BjWkApWGsUb7KxnGdd
SfNPxCPKl5eJI8z/SWS+JAApwUpaYVUawqGn9vGIw3tmX0ui57hZ/OhOdWILnb2zj2TsxOLhn0AO
YnW2GAFrVSyXBOArNWtMvy4jOmigBj4J0PVWGWHMaycfC+PdMzw6/wXDnN7QIKISlc0hLY74O7/M
5qNBs5oFIHyReGuKoJyr3TaxuGRYxg76wcjydVWEH+Pzn3QJE7Lc6k6BupPRB1HrBOPOSYy7dmhj
hkwaWI6+kILbmPPtfs/PeHV5vhetwfmsijWyiGEC7HcBrbdzwiVv/V9mrfY0mw+qLE9HOdwk3Z3d
lAtgd5ifs4X4qCprTlZTG/ui4kZ+Ikq8iTrB8IZJpa6il9SSHV8OcZNSR6vj61KGwAR9Ah9P8TZj
qJrwGpFmDkKbHOOrPPaL4Pg3N0tk8M1VSUFrWyLS+UvS4yxwi0yY14GEK+ESAkMZfk8j8ZmhdXir
mGZADwWrqV6EG3aRj8ex9weXLn45bjCPWg6p6spfxLrh4JpOK66kvVYz8/GZ32z0IwiSrom8I75T
a+9J8QQVM1e5/lD0mAk4V0LSK5bv0j9mCQS534ZIWdrWgLDcShG9GmOZu3lTEoNolAUHWnsXeruH
YKjwUuRfXVRCBzcJprvBDvss6ZQwBhkRIjHbft3iuGmCuuIMH6myYlNQ7pkIvMxZuX6GCmDctkSg
6QZu2h6BqPLoBEIopiaI+MonEmZhgE3ygTqVU9iFNYVQDuQVRIGme89dw/LynMcdUdJmIe7n0+nw
XP8bfKmAZRxGttq8GkJrLqSBwgQfoCoDnCRVqMYJAeCN+O4PC7a5DyZeWjXwO5GyxX+uEDVVMoWx
4+fu7FuSnyNsa+2iERju35L1ERPPpJzFxxfNvFEzzisxtiVYhXs2Nfu4IjTWmv7xbEYRsBQPBVAF
hOA2eHO7f6UbIhxErwk8Udp6IFTPRqtCKMNpRCed9u/6WIFu76mILMJL4LKHV3SbhnuK567aHE76
bxG//QqqzKW01UvAB+sEuCi3Doen6NUZPZDpnRKTSYsWwInMmzvt+9v9k3be/XIAnK0fPDo0OYPp
v/KqtXOpHu0psoIXdSIeuD/JKxew+YagQ+V13veOvLXPiD9BcmS5R6C7DGBg7y07afRo89LgbopL
VnUnhuq0hsfGcjN7fG6nZW+KJ7lIvuaAVOLSF5ii1ni5DjUyJ4e0HDe5R4iibslXzoDvqwrzO5/N
ZRsD2qWDfHAitslvHBYSNIYdzQfrJvIG4W7W60g8tY9EQaywEkq2fupHs5QueNC+o7ngkP8/nBHw
hGmIghDanPOO13eX/lznwHrj5T8xF5wmWmgt7DCWO4TBAWqHQFbfnp/anx5izGUSixz2d9PrJMMY
gxFGGEyf+0fSjmkN92ZLRw6xw7fh1Ke1jh5rRVuXQI9cHPtJaQP1Kz51ss4W6DgGEg4xMnnFgv2i
XTUp75FLRQE97xB3eQ1YYLNdScQqeZ5fyK3A8hOrmJ73CrybN3ppzQrlKRyGlnJkpUhnq7hb+LPD
f/FKE/+1frds3zx3OCk/EdO82XNPmZvlE73PgmGZ5c6u+bBm+32ebxBQ1V/swy7krUHD7vYu6O3e
fdDANJ5CpMbDdSzMOhv7OxtAxENWvtTSxdDdzzRgNDNP+UIKvMjxjMvx9/5HtuoquHEeg+nu0FGY
ONM3JR+KarH8arPF73Hj1ZrNd3etOuqOPepyd4mQ3yYfPSwcQ2JH4n2woIIFlCir/1mYwXZOdNaJ
Z5Bg+hG7eYdp1lH0CY06AA+27U9hetRPKyPrDN6JU75ZeSeBMBt3VJ0bKeV4NaQMl/2mXB//yKNh
fK9nZivN1CmiNOvCcZA2Vjag/k8xzDSH+WnI4l55eeCmSAggEHvcnwv4qbsxI0vEzHSWM9PlVYAc
68ATAB8WSkNoAtzYUIGyeNEUvGI0X69kOw8UOlF0Yahz9Uf9iXAHNEKvpfJLcx2OXcMFTf6XBqnE
EVKS5I2V3BzpuPX/vQSdqjZVaE4t0ob0Z41HsMOx15Puqm8BHte3UTIZ8lyOqYXc9D8ljksfACyx
39QOUvstFl5XIFN+DZirus+Ntowvjuq2RP37RJaKFoWmbkXdUwLbJhR2kg2sOSFaDtHkA1wpAPWt
FFUGEEPb8UxSJShScDRw52kvvHaRdnYz8nEraqmQlHaA0fRkfk+0GIBTZ5JPRgQkCWYuqvyhqooG
clgosZLLt9piOTJEvDOC3KVtDGj1pKyrmletsFeZdjDyqzQ0S3Viuf0ay0FwEcw9Enf5ppY8N0lF
nPbL+oN4kzV1l9YJneOhNXSettCygOx/If0GzVlXZcyw23nlzNK2VbGQBZYk+CSuy0EkMJg6TMcU
n5vMytks+tasYOnGUq2uW3rEBgp/cVa3dmuimdcfdpuY7/ROYnFNr0nmQrkea+DaQ+oMHoh/XzA2
K4p7V5iMPF+qsH+X2/Wm0dXl1IEpu48m8cI2HrrMybdwohz8QiMTyXgp0zWgzms2+cwjlvUzROEt
ETZ3Hy8kfzhR6xL5/+LYagdfTYxzr09ggUfA5cUhPm1aegCZ7Bdk6CxLctHJwMsbYN9mdiJ3nH/z
ZZORH2auWANEEsuBFKiMPWv4g3W2tWvA+kvgJ/DuWj6C3dOvfRUq3AVEMnzf6oBGbL1PzNXXx1Gf
wnfZ8siD/H6tL3Cx2n15XzrCRDQOAhzohKO0r2Ff4bXheCphTxVFYUADX1E+LkQtYAq01qmPBNW5
sdElIYs7AhrBQrGNCvh5HcBQ7hmBu858SnMAPN0i0sjeq45dE1nZ21cfE0BgebxvrHXMOv8x9zlI
+IUbHeo8e0OWPj0udlyTv4AxiZlFK4Zyi9NP5dj/7Mf94PFlyA5Hixyw8TRqDuTz8Gso4QeZi1Ed
qRqnZHCUj34EIyhl1cYlZqdZg8T2Qa45zJRZ+chow98KELRbJERwHaQaWBZpaCUzamBSdLIUPkkP
eVAMeeynqoKJtRXf+CGMyvSUMmh32YsjyglN8CHTFUvqq/SljPCh+Hcii00j4Oc2kPNF2AMboGPG
UimFpNA5dZWPeCQA8G+Yy4Yh9vKG2mA+Xcr+hCzAXNFw3LNto0fPkxdMNlViyYC24c+QgVh30IM5
oFWJ96dqFPanHbXy6ySpIi9XV2gezq79wiGozIjhSsRuUiJ9TgoNiPxecPyKsMpSmE04W/3vjsub
cFMkXhRyt7kDPy2ShKzJtUX/dJAWHfd3KHlapZBfxG4gcPZxw7PueJiZYCco8/ILaUip6RD1K/se
ox3ZOSSDB4SCNgWGgfVDZJAd4EcF2vi9QVgO1CfQuhUo1aLTtxVvuyK8xKnf2tLgIV+0c9P8Zvey
tB5Bceamf9ErVP6CwDVZDSRz+odSlemr2sx5tCcvVM4rX7yktV8Ccl58rxvki489SXuPVNLwLBtm
1NF6m6Pe/jrEEjUn+jB9ZPQVMK/AQR5lmK7rkTtPEnAb9scx+hSmtY4MVmvDjZ+77DR4BsdkHvOH
50BtkpyO85JaHel8OvVpHSpvCHBMACpU1ypVaRSkpiobjdBN0lG4abxUyjLRvBIte+XirvKQZh1A
RwaQmoZIP0rRruYApYd8Hq58FSkY7uGttdehtziEtICwQpmejeeRk6EV308qcTeWiQ7EKN0+i+xN
rq7rw7mSX2DwXFA7xFgwoYxZ3ES2NQC+QKCrUvILQoV1UzcyMKMdZaJARHz/zDys969NWhtgNWLz
ffoCuBr86f5PrsejQbdky+PzTNUl9hZcYM+mCQKJRePsUEqg164piK0pK8BXrFgiLGLYkgZd+EkZ
HX9COohaIrNV2RJdUVKenz7/pC3K8pz8WC7nGoDdAdg1pqyu55KOupuG7oebeL1mFOp0eJ2wT1fi
QAlKI2CGpeXe+BPyWT23MFwgRUgiflkOa2Nbybd6qoCPJp66KEWHQp7yqJY5KjUjk3R9rI9csyo/
W8jd/a4rivn/YnjWb4a1EODwNmlpPgcAMUeK6eUaE0E1aMQAibsj0jr+x5b4MPlx9NAHfbx/pVwU
b7ARvOX/H8csVr9z5Zkmr3OaRzymg+CSVQdP5GNZGMF3Tr2a9/YOL5KD+ENn/qG/uHHlbpYZ0l1i
VXqTcVPFx1Ihy8mlQbMT3e5B+kpPBZY5mRttmt8fgae+jzqVeX1zRCU8O3FJrr4aVtr2IbCUwafc
IeXAMqoZ9wHX/iWOToUthiKAkvQYS8FDfZU3uJXwgHMNo6OafVWPEPGnIX1/ceElx9dvW/ZwsCgC
6zstQfRO4uEWG0S3nt23my/az65WbKWBj6DrEiMnAd2ZqflG4yikAXpHM8kghWIZgzLYm8EkdREK
+E3uuoQQIjdv0S/5IQzdVsWiRClWsUvAEXCxS/7aGgoa+G1o2bTUXAl6+wn4Z6/ewcfc0j/TkmQ6
UJ22bLd0YqobRgPvVfMgJxQDvh56zRhD/UKqhfBy8fqnEeaqvVGiHSuE+KYweXgeiJ/NVHJodiOx
BUBgBGSOdFb1VFG51kQeHQG4rFFVqlEwahVEYH239CPxwIkU2ZFeMFt5LGzVrQ9qPJkpLUmJm34C
bBiBn78ljV24YTOTfRNdQi+H0y2nxDjN2nHr2uGbsrjVFwPMNIVpnIhzYYjTAbsNCE2CfXF1BHed
Nx66MZDhjM6mTSDM2imUa1EvAHh/rKUZWB4IQgEjAgCs5L/tosfP5sIievZTeEIDtl+DHIZDaflw
3KVcljvCRvbnHxQWb59T0og9BVHYJG8xp1dwAtuWHRPUKxMgOOi4NcplQYG8NiksZF/mixicgb/b
UIbWHLRdqOJ4vzEDVe5o0eQ0cqMvfqldePp9dIFf0xMwUD00mPxojfA4ycVXRczHb+9PZsXXRePh
M2OFcz1S6laF0GmHwB0gDvj4jePOn3tbbomJyHgQ8Uc0Ou3seBs4SpNPPRvxXW1nztkoikIzksey
W6K/IcFc31ke5NDKxjtsniySUMsySf0L3vOU3c12y0oSpPPrmcl8lZ1sRrtHzc98oek/P/Mc2gIZ
18o+jB77gH87yW4qghlGido2urawqgfHW1gYBqna/E9OXPe1RLbi1PQ7/8XUfYX57qrdkialB9zP
2IQfDDyrmyXmwHeX5POoQIGpOKe1FFNp5mJc6UCiAcuVWMJP0s1ce9ApPkGMmLrtq/649LOpGI9X
SgMpldeNSDKEjJe8EssJtHSnr7F9DoYmPtDBUneGtUqFrrp9zwkP44gV3tA7v+wq91UfSly3RJio
yK7wrXq7PdHrAwHXlFh4hPr6yk7xSP/T6hH1HcN0nxgv+9rDPqog+4WIaThYDHjmcFdYLI3wz2oT
3EcmcAsn6ij2lavrgremE/zik92D4joq6Il1rLTRX9YQdK1hlxx+58rqg2s5WBX0JVyi4qA+PcJ+
nsixVx4RnhtAK0jyNs16Q0LEis8yF8dbBTKsczriJuS01L8AJ7fekXWMrN5HL4r2g1LHiDslX5cB
pxp7I1X9zl6R99e/p0K2Joi+BTo64Wn09LpHs6k6HuT1KjkEj11Q8D2XDV6sE2Vo2RwlN9wzfC/8
PVAub8RswHkvHAc32W3H0kSMMcpU/WxKuVYWL3P7OsdX7bUfaArXaA4Y9V9D3HJJdxk1vjF2QZBZ
pvB6x6CDoZIN29Yln7nazr7tolTsjaN4rx50GQrZOkfxKzYycO44ewHo9pU1r+iQPc7UZNxwsaen
IW4sKANSMdqMz3XpTatmXn4ijKxYS8jKDNLQ4+4cNlVHn3qY29b7IyIvjIyKMLxgHwnstMCP7/t5
ZO342cC+YQH2wjPNxXAiVDoBJr4Dcy0YOnffdn2w6y3xsu6xsoJb/LDmQ4bFV4rome4odY+Y5q0n
rQroVoSLw5bvyaCeV+8oe370Og8Dy5djdnaJrjRKO3Mhl/3jWi8uD+9jV26/PBuEM8NlG5S1su7T
nzPbwiY4tlxYNj/cEqpd0TQ8q3LE1bU3hvw57cB3bsJs7rClXL4MLUkeb7Hs1fF+0LDwF/ToJPRK
X042s2ZyarkLs17Kbnz7lsX4N0JlnMw40oDmPOgqFMmc6fm88isQ2QopckijlEM6bZQ6iCJwGc70
hXdgfL39Jv7HilCO8NxZGI57kQMpcDt05EAbmwDtPmvYfs1hf8g8I1z18Yps9brITI5ZVVx/F+aT
nASXUBB5tGbuAFgJs3XC3AOnUAE8XJp4+F92WNXLOjG/FlIl0zYh6cYkcHonozfZfP9xrjLuStb4
wsaAScBPVt9v36hdUOLJlZfrKBr8PlxstQ7DBG2E8B2yCFvdJc9sotPdrGY84Loqz6h2Xz0N+OcY
UBjIU4f/qMHluhARYdVMYdGnSRBDZhF0uugTwtgnNBilJt2rOCGYOtAkpekwjgQpjffNUCfztkFW
xeZBXokm8/G4hX6d7S/qYE29/5jNFgFASHp+8STzuO0TWl5uDjqztxe71ArfRYDo+PrOZXC4lWXs
Wh33scbwwTIxDQWIwn21ZXmp2bjM5MQircDoVoh4eiufLPPcyUsIAg7j6vOMdidSYbOCIxaJzPTr
OHJ7wePqhbXAdGhWr/L2TDc0JJVbtfQTquq/t5HzbyskdZWjIbxPvVhdZx75QSrN5Cic4LBuHyYe
l0+UwmKdzqyvKWdaOLxaDmNxXv1sxHbOM8gvr0mThYTaXXs3ym5YzM+85xX6RjwHfGCJpW0srWEG
jXRnxVMuWNR7DekR+Kglj5VeZ9NMAKIvmQyYe/HlUz2hxU35siBO3R/LnD+uFmgod//wzwLgrU/V
EVy9AG6cEcV5ZE5uGMrOEwGKp9ZZxOlcr4c+NqZk/CeAyP5B65bCSQubrUa0naZVtbyJ9F7R9Kar
1OgFDy/erjYBZyVClYabCrlsUy7AuHKM4prWBQ8gr+3oIURBJTg35Rf3g31CEPwiQMOtxKa3gsfG
MbZoOgqR5XTpHHXlMwxX+ixfF1LzAAuMWGC3PrTKnoeyHY7k6unEQjZvK61w+dtJIFuGQ8DplGNf
zKWv62e3vCZ8mfy9vRFvj9CI6bbCki9nX8XtU0w+vVuZ2ppCoBtIInRXdvfKzZiuaSyff6cpqfli
jjJVt2KPgmsfF28OZWMD4kwDZSDxj6ZNwhrA1QWn/LWF+/eVOfLeolHithzQA2MDf4j/XCHG8qQg
3It0hm4tbB4ZXLhKrMEdYeoA24k+cvTaENQAkFQMIdGyUNolQ9FB4z6kYNPhPEARCXA3qwgJiuxh
cQPVt3uDrG5Wq9nEEJSm1t90StltXRMfe4cR9E+qpqHVnthIRiQ8X3t0l+cTDBwNzX63byUgVVR7
GCc7vP+IRHwVnQdJgEnTYf19lMJjsekWGNJDfKVf/5BFXxMCKnvN95o7IXE/ysE2d6oWH8b0FUHK
JUKWVrHlnHKOAupuhXikBIaqWwcW6kq99qF2FhPQ1smpIUC7AIEVETwhOXje/yZTXXf2KD7hEzam
l0x6PB8RSqaviwZdnDZ4HSZ4nsf2AnSGu90wLkM5mWf4ZQhOgWJMgTTGAxEnXQtNxyGQd8/7/RfI
DUSXIpQfVyVIQvRcxRApvGPIZA0ao8D9ccxBClpTrDjLUpdo1FNkcjmq65Yrrqxb40YNpnFoFUCA
bDpsndbK3Vy47dPZK8G28i8SgbDt7cACL+DXs8He6Ij4GIMTQ/C0wtBG3jDapq2zKFlKYb+mQQOu
XEk3In6RrhlB9Ksyq7Xa361uvf50lxHnU+bVxBsSgZmTvKnzp6BKRq+/u3H36lt81zS2Y+lJmz0/
B0S4vHFy+7ngQuLT17IspRUYCUIqvhPrNYPjMXykiAhS8Kdmyaw8nomDwhGAEL+mty9zaLwm01Yr
qEHOt6dvJImpOnNivR0QmZsTmClzpW6YOF3QzHbogl0DqZ7XFCNsUBWnV2uZETRUw+M/0HPpmJUS
QMXanRH8Z52Vs/LEViu/O/ergwDVHeh3HxFyQDzm2M2EHuoXE5SbzoUXbReN1Ns9LrqjnFHp1Ugo
q0E+eA9bAHVMuC4Q2YLPVk3nYzndQ3TXJhWOLH0fum1nUG8BIDvmnBDGzVr48kcbKsko+ywiQrce
jqdv0FgjxD9/qUajBMq6LKAESouPx4V/sxKjSY/US74LiEyc0B5eI0webAJlT38YBTJ9766nKnAJ
bPpjP/apda29eZ95ZtQOSO2EA9dbIC9y0djHoq0CUhDzAffRIyR2xzzqURUrG089pIRbYY3L+BvT
XPeTj1BytXtAK5AnVv9VGBtw+SFkFgNQPPNJW/vF1mi5hNbOn1sv/SmIOoLRHJIs1YueDi98xVua
LH+VQldJL2XCgeJyb0K6qoj5sji2MbsxmjPUpubwe69iB24vmllQE8doX0WLG6x5M/lxtP9NYUVu
7bO97aaV9rltN1fID0l99Lftg896TDDs4JMuWNsE53L/Ud5TI/y5s/HbIRkxqASVaTpwjV3GT6Wn
9I4aG4H8pRPAlOGWMXo5nwT0C//ug76haHKe5k9O0F7BRrxDyAxiVpjacWe2UIe/jSWnWpa0jFFR
kSRmPMI4e5Yp5tWMFrDpKyalkMAKK4hXvB8TXzvJKqtPN1UbSqR7HsAc70kBDMlJlpTM7+6Zw57e
lnQhbJcgvlZWhjXFkU/CSDlXEvvElshI+CxgkaEN5EiqbSYUladbAZYUofSbp6EFDTkqoEjg6AB4
3Rgw4ZtF5RpR9+ydC4BE2t2o06zmUwr7iUcGqf67u3G1zXSHygux/qR6xi26gBwSVKstzkqsx97s
ajSPLrThoDqNVm5hkaQVFKoRsxAJU+zJe3CNSbFnQDKqqGY/DvHU2NBWJ2/JnOXMVTgOlSrnfQiI
ktsUJQ2Ka50H2076UVlJvL+ni/2YzMarY+usn/lzUru33GH9CZYXiW2Z2O8NdcLzild9DU3vjhOh
C0Fq1If7+LTsgOkWAMXpc5aIPyTgmyjGDDqHra9cnITuJB+BtIM9OTE/YZ0J2nXGtsHgbHXxynEM
WPJSe/JUUvqjuuf40T/wa717WpOgsU6CvUkxlFJrsZVf6ZVZcR8ioQoN60/gMym1vUet9mahdbJ1
n8LWYcfzNDyedNB6xPei6i8FUelnVXygrZNLlfTpSvcUgZ+G3t6boIWY3doFA+/eGdT0tcTrWEK8
q/PXPEWPw7biuxS1459jtFDs21sQEr+i1hbGc+WBl6Y21cOqCs+gTADLap4rh39wxCzAtIsomBdy
5Q6RYy33krdRcwaMe9qDA9vXZQPLecONtRBjSeLvwBOV89P7CkkLp3qwTGnRUBBbOrl8rwx6r6n8
BXTYqH17tLLOE5YbkDz1Zbq6lkfeyKMU+ziwr4Kw4L5Bk9yBkIH3N84IolPb/GrHuZuWprVJQUBx
4T/bNk8lPfc9ENalw/4Z9HJ9ZDXuLUtQjW/yepwipLSm35j3+4lKL74LrQT1LexnPnsC+sSspVRk
Zk+DmX9a0ppSzJUubDXiMeGjMouJsv75SPbAw2eYyVIX7LERCaVzFqvHAtNQhlcnZDgScHXEpjXy
Ak0UOFk7BiGjhjUAtZxgxaICpdOjMoQF6BfVzoJeqFMRvCLgJf934MfHP4BhyOhdtyp0tDqJ8Vo2
koBhHgbXmQG9Pup4OIuaB3rbbs0wSi6t42h5VKjqpf1ruXcjCiiCWvV+KYc4ymeKhqvX+cTVMMuo
L+hw3TDgRbq7y6+SzI+mN4V6CTYgdToYfgQH8f9TgIJ/EDkpCi1ISB5eL444btGxY/INYkozqD0w
hos/p5N5coFpqZ7yTWYo/cUqe5rv4J3ejOhRN15WtbXDOPEWnfq28pvE9etfuhDahkT8wzPyBEMv
dUSqnksshp+UNlpFcX0fDxtCgLKGc/OlmL4oAh8d91TzYD9e7ggBWLImHDJ+V9f+80IKdlAsOGvJ
lSiB1pndexARrmXlP6B2nSWFLbWqhGXMsWs8h+YYHokyV4zqGeaFZWTUQ1IaoH8aHTV2eBHb9obc
ZADjfChI3dAoaBUwGJbhXvf8ZMpO0BJvBZdXRrIVal75k1UKle5PiQqpA37VnWm35X5id7utI4tN
yOGEyoUQqIoH96ZWEP15355W9O1My/A6Kv/h9UDBb35vbZlxkxSfnBHbTOddiECp3pG+eNZDjJwn
jPoZlLpNWNBwv9XiHUkMZBiQ25+thHVROcebTTrv8b9uhVLuZDQy7XOXFBROo/Y2KcrzorsGVvdu
UUpfE5Z/wTQph3oqBScVKORnGDnj9XDlcOMmUuToUj0nsoqeYDGTBHYXd9vrL39OR0Ora9uVx73o
kEhMwaojkN/2SWMzwQp7a0SxZ0fgT+HiqG09CtthKHgjLbRvRyXvtAxkYrQzD6LUoqL2lZidBaNz
Yb2OrdQzbkHw1W7FlxXUVRPjxl82IvAfPNAO5bAtVRAzuat+sDqH1FYrj1sMRu6U2fvlcH3DEnDt
Hmne+7lUJSZ8O9Y/nf+ZRMPmZH+accguQDMTarsrLN0nYpOsbZN6O9XRBEWUx6pJwzA6YKLjwYH2
MSeDWxdJ2J4w+kyBpH4rsB+FaX8bH6I4bbEiWDU+sRMnh4jCorkrXX8RpedCupc/l0HXgs4gE4TG
6Ub9OXHs7SWwkyiFjPcNPQJ78GQhgCAnMdVs3ahtlrLAfjEw3IpPZyoN7CJlL6Z9yM7Hq6T0CRNB
7h3KEVw9+TtJlt79vaE+WyA7ClnEJb+z0LIZgj74SjVKLJq1tZjYpqVLms1JY5QkGsfyjHYOWOo6
dSylMCDYqHeenB/K5ijWZJdKo23dCOuFbFIPvZwvlfmOZQWHTnWILo8XonWXJGi6GJ2S10VMzxaq
HDB0HPFbMWAy9Ai3lsMpPMGuoK4BnhEk+NKsgYBll2VEu1guV40VyNUnL6X7GI8drht0Y2emA6Fo
tUaHdrEy8A2Nw2dnsWmU2k9rF2QNy/jEhGp+4L4FDsWTCP72qhhC1w0h0jM7MNWleMeAcaMaBoZp
oor/ioPQF4dhhIuUZ27lynhDetYLbnZRixfTQ1lIPigChVqLxfKb0y1zGi/p0wzfl4hUWC942W3c
vtBTb9p7Ub/YQQRE9Uxm/PFMsxY9BUdwyETZ/uVimrWCAKuB+Q17w7hxc8dtx+6ClNxu6TrobMWc
M+W+9yCprMw1Rz5sgN9+RIueK9OL4CJzKO/jWMnVk1pE9qkmMpXJtGLkXj1aY11251nEJg91f2le
5R6l+ORwmhiT+WDBQPLLnas3AVYdqcGnk17o8XdyXxDexd8RWAtSKu/jnr+nH+ZIZKAFo8cSKM4J
ZEoUi91pcrMYwN+MZN9YdWN+RNF5Tyb6HgZ4Xm1Jixp+57AsACdWs42a/SNt+CYrGpWOT3gmEhCG
tb5ci7eZdqL2Ylq7B/dLcN8B+LSD9yO44I/iqsmZ28GjNYr96SCTsd+TkhfzL3ofOKhEM2aAsNtK
3kL7/GJ1l1oZqSDS7Fp1HnoOgsIHxhBUX0Hxby8MEgFco2hRVKe8yN5PxOAu3C3VtrfSo3d13s4C
fRKEq+sTFITKFjho1jPW9TPCCYiX1A6h/SD0ekB0M5hCqayGQPGXkvl7s+dyf6kQYAL/ckKCYknk
5cTVWuhVq4l9ID87L/Ph5FLnvCeRM352/LupF+0ebGTKtXGjk+G9fahoVZaCnCLZT94adjj17GuO
n449+0r005D2bvX+j6dNSfUHyTh0GdXlUBsCP+c+AelZdkKGXy8pQrYlB/e4vdCIdKE1dKAhkKJ6
6QRnY1b1EVgVsdoSwnSu8IArV2h+ccsktAbBclqwZxKr7TRLGCfjOBgr7bbkLKgPB2NTY6u3R7EC
invR1rDvcZsXOPfskzIkJyStHTrZyp6c6PImZVMxx1AbOAtLeL+l0cPornJ6osNrf7egaLKNZ8iG
MU5Gy6oF0BinGUvrFHhl/36Fr06S0l6wjlwionmA67WtLlYOVu74nx748pm0/PnT4u6rL9hfv9a6
DX0b85C6Al7Hwg1ZM8Gg6afhwHexZUULr3yIVx8qe6X9Pc78Ncw4v+yzV/7h0g75lKe/yJeJgWpU
P+9Cwapjk2l4Au8jBaK6HegXppJ4fy20kypn875LPwTq+lcWodGKgOfcFnN+wfdLJ3m3gHnIrYlo
wdfEOSH1DRCOb71PvKc8pMGo+MtOChK6T57iqV75kT7kItmuAJ5NaNtertrw8ELlbiG/rXeYnx0f
Hm8WMpLEX9zqO5/3ibgObgSulCI3fTerrRHILyuHPcW9ZTt3ehw8HlcZjgBK8fJbCackWSt7d0K0
bgCjpr3/VdtwKNVsGCcKsap3NMx7HpkV0EfWM2slQp+F94ISsaBiOGg+Q++2mamFJ8Yt/qeIergf
fj2u+YVA11RWkGciped3HBUEkRCmjNDvOJJ85oDF5FmB8RxMdRVnpwt3J0JeDlb4OjiaQYkymUu7
GB0BBz2ekxaRHilAP52ZM90Fx0TlF7DXUmY/Eb63xM+kNOEmVpQH39h7hr5fuKob3JLIa/YDqGq3
udYFwdRiEq5b7+wImi546aABfEdffz4kXuWrY9A6psYwpXUVGha49Gd04dGxERkHUw+tE6eb3CFX
JzCDucNXO/TGGdKM5oIwYIgjmn3hZmi6UrdgUyyt4gNw7+iDAV/nMyeagjldx49pv4h18NEcELqT
RXgkqcrDEjoi9/n3eWEmG/mmW+6RStJ4RxTcg9yF3fdror6dKdILm6+0rl1/I4oQQd08w11eug19
IbR5Izhz1wxc5vIpEoGO8H+shp2YGC9yJcy0ya/Ey+SdwbjkMrTUWEX4vLIyrZc4qedTYAM10L0y
rGkXjetrbq1VhSs+31RlHTmIxRIeaA3Jnsoe78MmubToJ/Sadp3fHNs5OHP67RTunS2KG5nC2H+P
Evs4ccj0OtTem9crW1YulHlKv6crcGqVsPlkjtgBk1HFygGabMD+T6vNgoOfs3PmV+Xv4iqugo0R
zKTW8+oB4bc+54FTwdnedNmBgK6smuARL8+1E0J3Atgu/TVGRtqLpOZnO0F41fhuEQ6DpC4WrF76
PzkZ5YaB4q3cWHJHRMeriaMZTqzZ15GjYdkzHk50dB7//S2agbfFP4rmxaoFfHdVlizUvVRSHOm/
WKzqYGVqNmED+4Q2MOnxq684mR6F04RkwvrDVjbJRcKX96FWKgI4yoQ6PjQyPXFK4ZK2pXxHE/qm
m2TDqthj2v8+J1ev60D9jnouS4FE9js9zfRbsYiUiGfafFRMOACCip+oNuBmmu4oAAPPg38BIXEk
U60p0G6nUhOhktOOnLhgJoPHvOLoE5ArmaIRhEAuPhtMLUwVmWWxnLbR+lyY72qrEZU9c42yRxvM
b4PpZAoC27TyobP+vkEwrMYa708RI9RcRALKQtvmN/Y0ujc2G3ElD9AvsgxkxTO8HHLmMulqZ3xw
4XvIv+OM0fWMKlJDpeJix/xDhJz24bL9KE2cWvzst3SvYp0AENqHVDqN8nNcxGxgQlVT9abz9n1u
HlgbcHsPsDMZHhluVNdOnhpcSennIbea4HON91YeKJ3nYPW07tOCPzvcafYNBiCxNYpoxoZBJNh7
o0gbbQGp9e9X+Kltz7zHG0u1ykXmjYmtCH7DHvCzhbaI3cY33yrPnhM+d3aLQZXSKWLKm2FBXC9V
IUhkqmY5frRSrs/bDjqp6rVHtLhmX0wYzMiDTc+rsvCpVHTC/Bj2sSi+yHWzyt3swkFtyU/Sjqq0
0ynExdv4AZAvW6L6YdosSYdgJ+cyxacj86h5dvp9VdMCVut0Hjuaq9VGtMUAobpwmBVm9a925DT1
kZe5KHPnOiZB6Y38EP3YF9TG+gMlFwS/ctpf7B4qd1qhIDlfZBE2hYG6hP3xfUdsyA1nSJvs/7rX
EKJYqunt9tsSauGygkvLx/9nYTFugIn4lcZtsbkR8iwZcb9j1p9pTZqMh0R8W4NureX0ncWq2/q6
hSDSLYsMiCUiTdfYZGHnAeIv2RnF3TODH89H/mWanR2A4oHG437Iq/XpMOBio/6pV2sjpIFHMaP9
7ovdAqr/98olp2uSA7ph8Go8sUMvfX6xT1H02VpTKVLXzX6epqHiOjPBCO8/dhHIAK21BaqA8Tl+
HNaMUzUMNUJqKmGxrrvkuVBvzzzlqJ6YieRH8srumyjBALXB5PTd7gGSZCG68pNP3VeLFvR4y/vZ
S8rgrUtM+lEtw6nfcYVI0L8sJyIOAIEwlyXcFgLFKUlTwtx/pnWLy3YCSjiGeyuaAZxLQr67IDpR
GcTfeEGHe81CH+XmeX+//CDnbBpwE02TR5QISK2XKT+3xSa2e240k9FQBC8LtJl8T2s59qkDMVAz
ZfcpDhXGVYsPA9uLPK24d2cH33Yo+ffo6Tn6PuKQ9Yof37HvvUiITZGG5KAa8nKsn4pI51dFP/b4
bjh2gOa6aYSOgUap6lcmwUU2nT9aWjkGzJOwXYAe98F9ODaA17d3hL9PCqyivz/YFFaK7DsFA72K
7oRfnV4MU/E+L2dwqZjmAVT80YpPcQgoGFm0OMvXcp9th5FzkZFY8sLbWL9Xalyt1ZnZr8gu/iyJ
/aF8UBrQnJu9h2NX3jDjdOb+v430XJ8ztCeZH7ZyCbmj9RNW3wLzyDHgcYewh/jd5bXoM+vvM7+g
6Ki0wJehKOvK+17AQCkeJWb2Lmdya6YoVWShzkWhyNmpJNLtGJlVFJABmELNsLEPJfSpgy1GkD8y
5LjuFUoZpErF8nnrrBusZkAPjkOXzsb5wdclr0ypi7qLbT/47ov0QJPA3ONvrGb/RWVJ32nPdsd/
rolUCDvXTVfN+0b48/0toSPabM7d8UigxddvtvUhYPq+w/aca5HT/uoc8iruMEKLaNXWS3R9HDJf
Elxxban2I5yfImr3kv6fXCMg3YvPNThYvQi7WWwkljWYf/Xv6FOnXO2Z2igEjZ7rxwKsXsOQg2A7
s81PCXyMTkON5z0buEybbliFtS6ptyXlu8amc4lgN6QXPobnR8g29oSCVtjprg1et1qQvXhM4FUv
ilQ9guDScZ0WfMjL6o+wU4+EOUTwhTkmHAWbhvJ7LMs7N5bLF28eOaWaohzN/967NHIDoM7vjs1d
c9T3jk4qZU26f8VAchJEg9l3k4BGFlZOKg30uop0N6bSJTCqczuvuX518pVZOZ5P3ycQKU9uZw/R
DCXSBiIiIudK8Am0mr3vNeGAj0iev4eiQA2JuF0dpgEHE/3jgK5msbkPmzJc1FthYCmXqDCC9y/r
E7ymzdF/E+zD78qiYfYTqa538HgotU/h8VG15LnYNDhJAPHbLJSj6gO4WaxLiVS9GyjF+suCwO5R
WxDDz/X8sZ25XUvVDGcd+4cE7zj1zsPbO2AbFSQEBIutGGa9yOrki/K+mGyo3SPmVR9BZwQmGzl7
bk2QJkRAvcCnjwNCAnm44IhbU/fQwXnFe7nh4EQHfHdSc+/VjDr0eLg1AOA+SNcQSeTdnUXcn7uG
P6nuhC9cVsuZ91xdQeBtN0cmUkb2JwUn1JRvXTb+l4wfHlrqREDPi4bjtJefLT7C7i/wvZRndJ5Q
ljjJ+Qfb8s2Z+1CLkLg62wTnC/O8i7mwVG6EiYzPBdEa6n20PnwWRjgemUiJ4obQhCOA+XdlR/dj
NsIRDkw6//kWCNzP1e6ejZZNt2pMXoGx0ktnNq7nf1UYIPAuWE7twG2gSnD6vnecjrqzHolwb4gz
I8yX3LJl9Vi9csw/Qcn9K6yeQrISELJ4LtkP6DSJ16zpsyVYp87y9DaIm2xMeDR12q4SN0cqSqxp
Pby24HsyxWSMMQCQPqj7mETCjyqol9NE2Ay4Nu/2JjEMHBelRxINCy2dr/tgKHMr86+PVz2wH0wb
YAOnUhmWlTb+z+wK/RL46acm2PFwd08AAFUkhAOQblrJ2a8T/ZKH35G3a528eiarH50q7Eq0vCwq
P8F7rl11MJlYQ6JwjJCfA4Wbr2sO1D/7uvWCksYTLxk+rNVufm0ohYY8HnG3fUwoGUbrZtXMrozo
8e/MeK6rKErTMcRwT1b0EICqlQpiAbh/NBuwAIh4twL8U6IQZGC/P6bd1MHpjkqwmM3vfX1TqkiK
pd+GnM09mca9eJZxRurdYti03+Gb/o0J69GFWbYKEaIsYO/vgN/BxxAjksmZcbzEWqKhlSb0NPQo
3uftiykGFqdsemw/nvHR+6JYFSakPNXNUGH7vYTvEy4s5jagcEHSKdYkiRh8PoxRn4gaYKjhDE38
n04uZXKaxaxJ4hhcfksX0cXSXWMq73YeGDEeYbZVQHrpraa7y2bPVTAev5I3ve+giVNGY4F6aFRy
tGwZdkiVfpuKjyUnG6erEpAymzKYPEMPzpYkfTmYvt2lGUDPqTg4xQ/ZWMWRSWCqxaWmH78T7rKr
Yd41J3wGEHxTyzX4N4NQOu727DEWnmTDtAPcjzj8wpF0b5efpcDcN4VygvwhK4d4XVX+wDn47d9U
UM0eWWeSCOT8oWZmL9KpMMScXpZB4OQnogWlW7NDToX185mSolqaMTM1+l8PqaxyeMaHYo12dM74
uNL/bc84rq2ijJmwIigbTOIAD2IKZ2F2NZMiheGbd6qoS1L5z2N3sx5Zz5Skq1RvKbMQM0v+t+Va
AZz6uQ98ag80Mq7rY37/6NoGYOFtL79hAoPxqlQbo/Piu4QAJohCeCKUDflajaiYJXQwpBlXwcSu
25YykCH+Mybhidat0XF1lymHdZBNa6AXyumINAie+C69H4wlNd8v8JYnjScHOMFwx9xX4nLoIXT0
zSapO+BDlKacxE5MHTEOut1I222GyItF+O0Ka/3H8Jspz+VtaXkjblZy1FueUM3p7cedp8R2w6NS
Q/sWRN5DtxQrG3Rv1patTeP+6LfsFNeC5+xLIFrMXig2SCPZhyu+Obzyz6YGqqxgOWlA5/YDzopd
0O72iEhvx78EUVkcDh7vUW5o/dNId6Q5gRg6LfLGhhrSf1SQmnEYk/z5F5FNT9TG/CuG6DgvoJLs
Oyk7j+2uutWmN0Sq1kF3j+bnEmAURvJCWBw5RIx7dGdWI54dWX0hFFMEfLkzm4YZ/Nxliw/7aL33
9Vfz5RlHJF51OmydebijQxcJ1wdo5/gZg40jefovqPvveyUdgOt/q2DXu20mwtG6XdDuVCwavgL9
hKlKU2hNlUYTk6j+VQUL1rtI8GZ41B88S1RnACi0ofxniSPRMrZytFTGLPSh/bh2DYgRDh5193fI
jxVlCIaxrh6kGfIyat1g7jORKwwjvyVirI1Sp7y1lKtLcwLnhJKEkd2ey/4skUWaDuIQBgVORCmM
D5hhr5or2zAE1563z3S6RZ7/lheTd2L/qlawT0bfMRuMzFCb728Xo14ZuCHAaw9MbsRJZJ8YIsNO
bMut9+GyXz7jeBG8G68D9X3qO2cBdBmWXyV8hbnCAo+EBusImrss38xIdbo/fWaU1LLEQAV1EULj
u9/ajHbVwlXealEPihBauaFIKJ/+37CFt9Q2KK3wkXw/SCsiQaLC9TU3Y04dW/bKXvNkF9kE5juU
9DOCf6rPSIy8Z+4DEnot1VhP2HltZH02bmuQKqvCW2TVjenPtlvhAfI7whQnUi1rwlHYC6hJ1pQw
P/LL5k4YYUQzY312wNNTudvzeX/iizm8pLx/a5PnTwY1/ZLTt7Da9FMyN2u+DRI4RRluQ7paEnWl
H2BMjAVMUqduoaRSb7tT8/DPtrQddFRFSCgLBC4qhib7mNFcaLg94n+M6Ow3W6yjknXZYL2BKSTf
rksxpk2eGh4ERDFZPF/hbuAhROJWTcBgcMwpmS/kkJRT7n+7aj8BGNPE2Q8dZ8K8CQglyI/KvD1z
PbdNO7BFWpDloH+bgXJ95zjFudbf9YigynKGqoPcBFlVOQnLSUBBRbCDMjgXNlWKel1lqElnIdMd
d5Ijq2wCRDfhFYh5XIv+ksuqTqsptM3Lr+UweTuzpPX7Pb2jHHXm31ZgKTAuP2e7nJuKteQudv+O
QdCG4Q1cx3lUdGHDTVlKkw/qkRp94hCNLHwd1ON5sVIgjJm5+wEXeVfjfPGJZZNSxdnvh9Un32ds
oC60QaBivQGAlBYXS7R2Twn5ZH++iS+vi6FQPFKrW//3PJlkI5TY64RduCybtT2c3upo04UlUX+b
lpvIo9Is6TyV9SP6aJERMuebZgBi0WIQ2W6UdF4Ecn+TbHcieZqzqksiNQLTJOggrKoyUtXmOBVI
zYEcoN5OrWyV8lDUg7a7obRWxl0Z/8ySRN1tv8jUqobKA+JD4ZfwHUsY7ALtrDq1QBIq0jBERd/M
Mms6kOOqb/d4vqrHj+hjfxlELxu1cRL+TXJzpNRn8uf7o6ixb5yV3Q8BqPfKaHU0ZnqAli5wG5Sf
yYsnCKkDG2ldgLbmqTJsuIEZELhiwxFfl29AIxBWqSh5v1/Y4XIi5LxP8ZsYB5yGnIXNqWfnIx0e
89dnx4oBPh6pJxt4LVatKYBo0ebeeflIqUydqcxqm6LjtWXbmFdgcWgtwvbJLqNx50k9q1uFSTX5
qjXNmepVnAobwraZ8Wz5CznY7pweUPsW8LVYg5ZUBTuVAgo/IXAaqhgXMYDCe9wUARCDEPJbiq6O
BxHV92tfUIcDSb58PEJFN43eqwKJqt7Ngic/EuESVYc1A0iI/zopDNXXFVWr9wFKMdDgJwLsUywC
+mPElg7mKuzKbWbwFhBIqOSYhzxZymMyfJ9ORq+In2CKkpvjRMOEYNuf8rtfugFn6xUxTkt+1H0J
2VQDQ4aOcwSJEugc/IhJrbk2B+rRPu93nmz/mptAkiWFY7N4gcZFH/IWA1UYLwbutv4cEYGhF+gn
GDAMpph0GeCKv2cK3V1IW4gz1nHZVdOlsLxkQQXo0QftGTL9SDl+KEhGassHdF5jw+GGDHyAs0qQ
ZZi0GYIgF7JJCTViVpzapT6CoRaCyKwaebAXrrJW6m8tPVri9b25424iQmFZm2P4AKyAfj73Cuv+
8edIEpEagA4C0R+8rXUG87XSGLaexNb+K2bHmt0k7OYfqjWgM31Y7Vfsb43TzntKxNOb5g5osjKE
UM9wqMeElGfQl64AjYJjKAON9xbtBVSf5Fd/s/6vhQQpOTddhJKw0DQHz9oIpJaAVZ5Np8C56/Ql
7cT6kuAlpy3yCJc/Kp+f1pLizrmOtEB+FqO0pNzZ2ofa+AGaQ5W0gA/asfpPxvXZNinqMWwhW/wi
EFfxJ0VddnwvzvOa3AAbqmtwSU0Hk2vm7FO6+pZVLQdlkdZ6O7wcfa/FgC7WAKwWvxSjTVdlPate
ZXZgTuEzxZOjGRG22y6igT6CkJFcSnsa79nvUnG8NAn+u17hrHSBs6GpVrPT+pluheN46jzF7rrq
M6Y+veXHUThB178kiVxtMKAfGZ8BTRz45KpKQTs9872F27jLfc6CeYI2QImwKo5lk4Wprn5SJ4lD
4o41+g+RQ6EFtxD4grKTAxXdXnB2etF5e650KKnQ+TxuQMyRNeoQ09PKi1Wi2F0GJ7hwbrlAW3pg
3f8pTSA5iLwRUaotlmlinlHD7GjUgn4QscVT8IDuU8UPg7FLM4/mEunI8Ngv9er8HYZQSayMqzg7
cEf8EQDblbOCf2Oy1ZQFQIUeSOHxTp3AUWcHgnzYMuiarKKPCPmOc0XcW1gUEFISjffTmJPDglsg
im6MbVlTQPoD0b0AWrnPkg5MBVX5RYC8Y6H0rx6D+w9T3IZs3gtvZueEj0msDt/QPsFoTU8T36vH
WeJSNA2iW2rKX1YQLpTzq1btTfAhYfgCqbcNb5LPWZ1XhRjcn3/owZZNyfElQeVUs8+hhdPfUCP8
x8hmzypR5eauXHqGK0QkiLdL3peN3snaY7oUIrT/lPOZax9jTO150lY0c4UrveixbtiwjXM6cvqE
Ig31F9q8MH/pknT7wd10ZMDxkOvMTV+rC7swGh4ubDW80jWQrwEWoJl2trHQJuuOiMcbVLcgBky3
kXJl0+FhzJEw8M/2eThHl2gMrqwnGSVFpi6gPhCRk7HFK59u55nOCo4sFbL81cMR6EZkVzFYLt/+
L77pd1Ol5syJxRg+7HEgld2jUpMSQ6GmHz6WL0b2YPLrFx1kwlOclXwQ/NeFxh8GRjOtU8JVU/K0
vyjRh9trWoJpTF2a1+WnrUVXOiViBk9wkEK971Pg+QSX6sqspc5GFrLxNvwhSjV0xmUSUcXIlyMk
hh7xBcamkhhun8K00Y0uBfnGGeWEWqLqS8CNt2E6OvGRnUBCou2d9v1T4u2wqpBF3PRd81Qr++TV
KXuT5Tj0BgRVOTqPCAKzvft2fmW1jtKFVFTpiplRHcvTphGUaxIT9wePcJvoPx9YutjQkZQBRWRq
91hAx/+RkgDrCZDxS0acwOvEn8/Y6M3QFoVNcRL17PdwH3CRWCbRFyp4bSaV01xBU0lt/qV86W2q
Le9nn4QerYJb3h3FsIfXkQd9fXhowCShYhaBFmAvRQ7POpzbh6bTTPzVsnf07bp0UmBxR3ibhlZ2
OKLY38mvNpLoydgEIrCmElRiWZQCEolnAvZm3S6ciwiXEmTgKPZ7C7eIcZ8bvwSWHHiooAd4VQcv
swHA/EY4vLCkqpBCj7hDbHDySxzXWfLlRF8dHV9j7Mkm2AU144aDdMvehE60QCrerkJK0bn+reBD
kK/yYpU+WtWzCGBU7TmJqFc1gM3x6xU6qUSVmQ01UOX+/c59NkEHTRB3v1P/OtefaYXJQwaMHbzL
ejmYenRPplc+ZgFP90wQoHmTJVNHkxG91UgFKlS3pWqvE0EdndIR3vMHuWAY7nC6Y7nJdXe9uZzD
vFTYQkainUVO2AxvcUZx/KGD/9ixwnM9Aq/c/Im6VDJxfWtr4nWfYECjxVkuOG0vfA9wl6IP59Lb
Mi/Kb+urbdFbhjj8D/zzal+aI0e3RTm1Eb3IYanR13/y+RAKgZDYdhfvXMNu49a7lkhCK4u0e8gH
h9tr99mGVQrhys4psS6nXDCM1l9L6lsIVgjUVSZgQsJpu5EqtAO9R7lpR6J3+ldhYmN4lV8J/WjL
wiNaAWoPN22YVWVjt7rupP4/6Bu3DX33P4bm5/UvMYM1hv6ijfuV/sx1mXOwHFS43iqNCYv6E2vU
gzGPmpijhZW3gyy8RguPFh/B2h87q1PiFh5EPCqSE3tNJgHRqIsx6aB2p78yFaKtxqJqWGMZgoqu
ZZg+JXnS2qVUfuV121/aImYXqqw4Y74Y/cOh/vfZN7Me7rFr9TLVAkdCWTyDGJfHDfPlOASIMjVz
R/+yyGFK7+lA2LOrT9D1ch0ccd+TcOhIfg2zEFe7hdMPDc4FVy7yV8PNzqZgt3P5t0zR2/3n8cC3
s38nPETIPLTSzl02at/zSc706Yv0LmsXkcXn4eAkVt643YXGe9eZ7KD0DUjn90UzjiWsF/kYwWmZ
4CAL4WuyQgpeUazE4b+HsUUayUTRV6YGNoLxeShR2EFwsmicCcuQEj3CuyuviFyR8e2vbElDTTkC
Ui1Q5XtRqH9I+yMJvgF7FmyAM8urUhe8ql42zxrr5gh0iUR4eKmlZtyh3EL5pRFKClUxRs2G2Axl
7iR5Rjvav90RXh9y2yvIWW2acG7XTcU2Wtn6o08h/2wZAze4ouFAVNNVsGxQCJ0Pmc2fISKLdbd8
jgSngnU0NbbG49Acpr3VFLe4MqsxpZI7PeDK8NFjPvqkLomtuEtYHqPnaX04wdv/yEPMu56QnCrR
/tli+76a3TnyBtGC8zXemAvzOkUt0CsaB9CBpWCrVA3N3Fm7uCc+nUC+U3aeX8byGroaOIPByPXz
/9Isbv3hwMnSh1qoHSutAK0vrQuJZQfyb1VBM0D/KSr8UQBgXbcgMd2WeUCfWWJdebxftb4e1sGg
JxgAsXJ31EbkFUJ3owqCsmh71BovHeilmnDwbQ22jufsUtjnSVJrSpLr57fOxqAQlgdBExxYBHc4
gJJByB/KlB92NtWizg052/a4n5WYFgqdBEJ4Cuqx7At68FvwPoWKoRmIH5Zqt8P4umsygKYaNXv0
ZCO/yIRE2Ql2BMeqzlr6I8NUO8U1Ioz3vr4xnBlzBzG7oeZVXKiqaW++j9EzxCXXSrsrkRTAEBX+
/KeloAPlw9gpDobn55N7wUOpp/SC8hvm9ImzhZhnl4V9/BadAQOGhmYz7YAkotMi2n0c4xgj60NS
KrPsgEprwmwD5TEDjkzSjKFAhK0WSV0d2ROWahKEXVMhYkpv17YBlDxce7grurxDiTvsrvTQNgIj
qkbMrauq+Ew8kq/lmU+ue+sC0SIPBs1SC8ytKkDgatoMx5mZeIdzwlpbDuvXRLzlPCLi+3t8gweW
xOzn7/K0Ba52BD9REuS6lG9tX1owujyw2AuyAZeLzfvkjx4oIx2nvZ3MISaXD5qw4D4vrJcLzGFb
W/ulWkUrYAzviX0OwMADYdTvNJpVpfkavjDcXWlRy5purKgv2+gWZTnt3PPfVww0wP80F+JOuUK2
/SJwjzoHKN7toClJRcWhIa6D2KutQo8hBJeg4SPZ72OIVjZN4X8Jr5Yx1CSc0G/Fw8q0W/thkV3M
8/mVv8DQ+KPQBgCwwtgBdYQrETp5DZRhJ6meGOnSAnQErbGk4eGJI+WUmuZpOGwphHEqLYnMfnny
wI6fqD0NMLsMq309j7udO/n6UmkvANkh3bRhgVizR1TC9ve8/MuPgEHNg7UiJRBHIVitqtrRgymu
jUIKadrDH1JE22vAxcapiwc1nHggTDx3mEKZS090tY/kujYCrC46adDObAGmDPTjr3n41e46v+xb
Ao+9bOPZiJEddW0dlDiHaSdPsjRAEIlwtuuSaH7cxKNuiFqn1TI7dKex4fBTgJGZtI8FnxrqCuRr
X2L4eEOCMM0tux8VsI9uUPQHMZNF1SGwflImyupio5TPw3qH1t06oRRa/hUQQVzpZnRX0+1E5EYU
AdBIg1pn3rOSqkD9qy/Ku8Yf17CjxWGyvUZOFkrhFP7YOupGuwJM5iqfs/j9ny15X4XeOMqefULN
+IOyKwpUIuGfh5MkfJJLjsWDPU4ceeIgxmWcJYFKih16skVTbwdu9WAkgVsS1c7vDEMd5DfSnoHZ
xmGbm7UICJZCBVX+Ta5NUllCPmE7vMwtUjgjWVCA1rxr2KxNCSNNxldjCxxI7gC1zNVAQy/iW86l
fHkSRf806w3M4e+W/lTONbnHwAXEA/JBYfqvumtL7a9XrFDqO8jx2r/f1C29EeLh9OL8ib+syq85
6anWQdSrBmAYvyXNgom5v2jn7FgVSR+/5UEjtvkTdV1mcBwFmggH2Tbtn+lDTht6HAujkCtQ4Zei
IvCuCSmbc3ngegwd1XMD7uKioV8xqU+OV4U24b1IFWf+7/yqAqDEv4T9gTooRPoEzX9tQje5FdTn
Ct+p+LfewasXn8JUHkFVvXXP5IfGac4JuPRdDLmBClxRt0ho2rPDmT+QmESZ7nIlFc39C92bLOad
HgjcrcxAH5pNRZBsZfBpD8KqyiCk4ewH9OSoEIujqH2PHWlHhNVT/9dLXJ8+pJumC75T2abvmDB3
edP5rECcCX+Y04iA99qJPvg2cA+ZvdIDh1LzAJZSkt3BR+0ZmRiLTdjOIY5xcaxh2oxaSfy3m/O6
/6zQQb15kwP73oRocE1itearSiZiKUj7hAPHyeMpsLDSpTcmEifvTEXQXn9vT1KZWQrMhHQkv25W
lOCzeANRAlYr2P+rVACVKkbGuAheHbnDaGP2+MDTnbnqzdupn6hCGbbQm/en0XRY+xg4imadkhJU
TktvmBmd9xVU5bzIVBMZdkI/ip4emiUYqhF6DCMJbB0qTNfnwOipGSG34lgFuz7lus9OHfF72qT8
WCO8KkR3JdH9ZNTyQgJTa/3Lfb4PY8aI9Bo3aiQIv5XF5rRpnBI9n90sB0wtTgitclFDwBOyZQDx
kg6xB3uRVgMZeZZf92jOZU1JGQmqIZiVZXsWUAYDyCJyJQEsvEIA5Qt267J2DjGfFcYidMKZl2qs
EO45C2yqYU7cWr5Y2RTXM4e9nZRaqlXV9JNnYpfl8dMWGCFAwUIuR0huSZ/bPhGQVdD8VZAPEhH/
AqUP15KmOJYZfZZJgOQm/ocCMIAyq+/JayeAMF/lhMKN83EdHjkkH4hTyi+FBdCAPHnE5ETuPlNY
NiLya7V0D4TzJVCaPx0cl2QPnmOdGw0LXT7ZEZ4FieoqL/vLMQR0pi+CYdLQLBZkllF3LhieQ6Tj
KPA6htHdvwhxuE9GXIIRbD5K8JfNt25x5Y2Pc5UbyFi40I+INPUgWRXRgUjnHLYNqo01Qw/0hgH2
8yI5SnEK8mCl9AdF8rgEbY46L6idJynnylsGAyj6bExniXpWnHmtIDZLNBiZvMXuHw6TaYY7nxtf
x9deoqe7hJSZkuKci89iQHJurPpet7PRFrnewKLzl07AF1u+BnEfI1nlLElBpNrX88yMmzjSteCL
37CRykiIury7wZrXyil1B+Pohsw2rhCzVEVcTF2njjXKGf3kk7omXLpOqGLQL+63eUsCPCY5xxKi
F5KT6HW+VI7l4Xb3n8QIkwMOnsNGGq6bou2uV7YSYFmyDQujwdVDWIrnE/h4poowqruDx+N/Mld+
BCPdZDk6mSpaEzRyhNC8MEOATXRXBmQi6rpJIyjChmd5dXSc9++JwWZZzGqmoSxpMLvaEskYS9tK
k7Diw7Oca6WyNugyiNDw/zu/skYuZXR/QUtXgNDQnWPeVZny0XrutcAoX09jB8VgVILBALJgqXhS
rLuah/3npEodMR4wDsyh1rVXETjEnQw/pzQA2PtnGcNNXjtixAenSTVtB/LNTsIWxpQ/THRaPh/4
kNNhtqT+y+llzIRDjRSSsXXdUlVtThWPqYtbwrrNH3dmnWVWG+H0CRHpKYR1qZkkycqLFqYg8UNc
RxXuiYPL1B8UIv4LKKFrb9vo8fouwpS50bTOKVRvOe2sKc4ADyOpeIKXeQ5plTPe/cVxb5DvV864
C5ZNOHb3/NBFjumn4YBboZrdiiVSXO9iCvMUS217CvRKcuepGpp0t2TsPIs7tVzNOfeH+gR9RTXl
1FBWK2zf2bbuVLb3NRX1nHSU9SNVO5desWtNRVuZHXtRFV6cgMZs10cqM5GJDSO0K1TMMZPy3dvo
b72X8jZ4azvGIBqa3BsGoxOOVC3DBMOCiOnrXZjNCcobZnLP8cp85qGQ2UTPgk22v67bskC6tiXN
+bkwseeguHikQfxx806eKglw1K4Q6bUA4WHFDMRYDW4qoKPY/b/EY1bVoFoPUWhMBRb+EWE6lmw/
14uMYP/42it6v6oalaNG9jnptD/b2RPjoKyOQfLmfpfI+tabC2LtezBVPLVHaawFuoay9NbSa5it
9Unucj7QUcRDvG9vKNMZHSqbP47p5S0Q0wRq8+sj3k0lzxXxJ19qFxuzlHbmtXqAkkrGhVzT2vDD
IuGB91Vyol1q8xlUCWUgWoeL2Jhblwaf5MkMddv1spqh1YAZl6VmXJSf/LlhCF3T+SRXVB/eJyTX
IwnT1oMLL0UM7BshJ1fUEDaw9pS3YwPFd19ydbEoKJLnuLpntM2YQjzcM+H2XadtsHdvT7ZdgdI2
RX8uJXWwKzu7EfyweGVNw+chtOPRgOaEfNiIHHo5rN6B6xt++Ui2p/ZO6pMcqRnP1EC0ASC5yBn5
mElXhn+GZP1TH5tSS7Bg4NyaNK4N5xO2wVsPggme3Ml4YBeWmJqu3lzMfBCq6y/hnRpm8AVx4bmO
PHFnd4dEIPL7IimQGShf8BynIcuu07uZK9WPWm/MkYGpxHZqWGgSq2Xu0DkQ1eaQ75VSXsF8XhxJ
sJavleoX2wLsgOQpwL/Lz1HGX3KsKaaGDZNfjlUnvx+qhBaboyqyA1wjY2tv9LUPzXcSTz4rz6O0
K2dOSfxEs89r/d241lIt9veO95k/j+q6KFncgqQ5DbHYK01a9kuj6GPUutctzy5WgLNKR1lnai1B
fBbhwX5NLomgQKw8gqAU1uofRV18G8EEq0Yl+NhDeEgl8N9/OxaFE6BBQIK1fVKrz8e4OQPzgo/h
I86PJKTBJbpVETUV8BQtrgQrlNBJUtarhG3bBOcaB4iC1WdbE8uBJEOPTVuDbErTENDQ++IjRMvR
Bgu0s0I7/qKIdOoYImCfhF0QGq4f5akITpB8mAH3/VqL1Yf3bbBsGuEgMM0HgOAPaKTVG0cxx/ef
htQoJ5Z9zIVxjy0W1Vj3uAoHVlg1RncW4OanMGNNZrO/5WpTiMbSgmQVkNrZa+UtM9TekVsIJKJT
nvJiQPWHSITTH8gxLU21OL9AV0R1kDmbfjjNpcXndaWqBvChi/qRmUx6p+/e9BlYo5OyyKJKbLeB
6gEP/fNmscHSWsh0X8PyiPPr/N0wEtC1URO6P8GzPolLZXnYSLL1n7YDr6DklH8pBgqVYHtjppfZ
+M+Lnm3kmuffymL38G4FQsZ2g+Ze8Y0njwIeIeQ8Se6ifGpdML/KrLk42jEd58vkxgE2f7f9RVjS
Qz+bVSyxcXJ62K6yqBHUC8nKxqRNWjyozfAQ523/0VC+tYr5t20LoKrraitP2mDHnQdpTAKvmp2I
FPYPoshfINPaojGj7F23OoLe4wO6evULB51CRmW/oO31J8WfxF5CBDP9iazNkYSV7Y3RzQskw0qj
grz5hhho8hB/HG0Quk1PHSbEkH6VJb6kiJfn2hUuiBxDKhoIdjTTw6SoPoW1onXDnAdnw2334jIf
tP07wiHeB29+OBFt1ti8YcATkxZaXX7jaI0iNmIjt6b0DfLXxPMJUctacyYl+8+hR2LeLUYV2Pmh
AVohS702uRru/5moeWez0s+EmvfnJhz+LMzawOyll+WORIjsK36YbbK8LQo4NLZHUW17rJ/AE4LF
KTgC4cZ8TyCoIIEL/lXnbIPpHwhLmoO+mSn8ql2LKRezmQ432bGqB6iJOw2/xYmZ7dwROX8cyr54
nBFbk5mmTJNXMto2UTs5N/mKR/0+K1z6LcKjL9p0ucD8OJH4TSP5hozCP8DNkc0lFBfjS9jYn3Mb
MxRCJUNtiICWxolAhrfr0QjpAMWD9lyFhV2WO8Cu4z5NPhw/7xS8EaVCkAIomvjic4rYDKKXWdAZ
In9sQ0IxgUsiCMONLGn6nwjKsrklFTIy2dY/Hx5tfvgZfoxt9M+1TavguSHEVeMK0wSxwXn0FpJg
4e/MQtt2XrRPuEB57muhyG1n5k+xIUy95Bfyc/LHTUjUaMMwbx4Yy0u9a59wNDR75mbpWKcZRHK8
3IyccJhHJePk2EgNCsUG9tD8bqsFbH/oH7dLoUcO5AHIoIO3V9c1s37qUJElCy68du1UxMHoxmT0
U8tzlKaW2G/k6gOjlUtnqe4JDuo2r7GHKSCksfboarbflhszBmD+OBC+zFmOE1rAuFSgGpzStIUl
qjx4C970Xv8VF8Vz8tlzPZuc/tMRcvUwrMWU8L7z8RFPBa3WlxFJOGuemWJfURfA0qvRQlvqv4bN
fKQEQvJNTUGR/37AgOMS03psDJPNJiD5/kZGKs6+sdT2kQzD3WQ6AmQ9eWuWAaxRVBJM6fWprmph
RNIdjJMho6qbqsMhI/Juq4vMyHHZkDtcr8WSuQMafUzPbYNwIz/Wwa9sdlUk/e8SrGslt+9B1sNr
Ak0zATBg3vhZwiRf8idjs44z3Ys5Fdub3+zvFkbi2HB2gkk/2AbUv/kXyJlCqalthVACqUXT4LdE
hqZfZy6ObJZpd9mMITPg6SXv2ikvs1iMYH0SCa+QmfSo1yaT6kZQ7hdzBvjTn1wZlnQ2CZnKnoqM
a2E9gkgpjVb1nboM9BbxLQ8rwZMwRmCe7YxhOQq7DMP3xy0OF7y7j8rKsZVcAkMW1wr7fdBf5tFB
U5zQeQnY+Q2X5mP0neAQ+ML39KyboEPOxF4dS2kWO2edIhH4NMPllW3bgrCDxAYDDeQvcpOMVVyw
KY2xBGr4GuFtnoDoCFwORawdild0Q1ZxwHfoIGaS4cTdVAbgp/O9xLzV7upLcx1/EldqqqUyp1Fj
z57Xt+p9v5Ve+igz8M3A4szRu0tLsdM4jFFWe/os9Dy/rEoq8ZInYStVXlSiNXrdoWI3tSgYs3if
chZKqk2q1hzM2mXw37woUvMNTkr1Edz1f4HNyW2ZAXpZLZtAkaHCUGjeEKo0eDakkzDIe3c0q6me
AFwuoRvERmaLUuvudpQ9fAWEHLxDUiw4bcDnkCujk+V1GOYTfFCxq9j/E0KVp8sxxdIvE1700wHQ
8VBK73rwXD19N2u4YEFeeyEDpay+TDo6k1JsE/SfzKkmbBoD8wW8ROd0ziqMDOekkAo4d4MAJGlS
7LrgxSNTrSKYrgB4OSw6KqxItu088NrtCosbc3W272h//T0SgKU/rjBKF2HoSrW8Z/pSjCVR0rVf
C9eEqgtkA2hefPCT59KgIKR3lw0POUyAHgU43OBKiAThD5pRHIBaBKyXVzxiF5q8J2jaMgw6I3N1
b5P0wp6JZz1x6Itx0x65rtckcMVPazSAVu67J1GbhQCyALO3/MjRl3pZmDSGHLYAXil/FmmJiyYV
oB+f1A2Njh6CdKxBS9/Ao/7ISeEtS3Ps2zoPGPudECPxotxCZiGqoJsNOAihLB29h20H8+ze3nWN
+kR1kzXukZUt3L3cEzuK3siGk+TEKxZQYG4Si5D/99UJGnC7gTy4Lii2LvnVeMFrbFe1LKHPzutj
Yj3YkkhKJBOq4ylVHCjExHCNQGs7b5PEEfTR3IKNar9uo6/fB9F0FWpJyhuCD616OEgX7+Qx1rzL
3cYerKPsNQL7Pvfg01kczBbeWYrnegp99dec/UeZfGnfF4TDIcgeBPZ6ZpU9uKpYv26ctx10Mm2V
J1A3QyizKCyZl4ZcWJoJCc0yXCQ8zrYe3Yll5jdpZUQYt1MZasoPLutJggnji0kJe4W9xroVy03A
eBQ5UB11D+KOzvHFkM9I8PKpu8UGBKTxG8v6K52Azpn3PqgdZ19nXXr8zQ3bVWm5PJBxRzxMWPnA
kEOz1mjTkUXxbRMQLczTcstA9lSngJZxTRuPLv4QvFr4xETknwmSXVWC8bJ6cKdGULNIlS0JA63N
7wd0fIWq6C1U6n+heszv9/SqrIN8H4oGKnm2A9GFRbLHS3W7Fj8DcbJMv3TO8dew5AOWZYl1rt3+
bsF2irqQHsfJMEi4OBGl5icsZ0MJ8rEE+N86jxUSYtW8wHWg7iB4mpArJdBQvjCD0bumGT0bJw5R
CyHJRcdv9ZpNy+fMgD0v3vw9ZyPzkn2SFeLWe70hyb+VUXMMoVfx2u/RuqeLU0dFJ/ut2//KOU1D
uiyA9KedsabE5QFR8C96e+bPX2HjxWpocJ4OR5o0b1dkDHdn8QyiqrzhsIoyMei4HE+Qzlqyg4St
pcjY84CcCGQTX/FrnxY+Rdv9lgmlVyIK74aqmC6Jh7nRM7oYa/s/52lPaNxR9x/eOHcMlOu0Ggpl
AHvZroOTCFk+iBACE7yRu1OjTIyWJF7gRKzQOB+LAlYoqfZONzABExkfGHGtg1XFFDQmsZsxbq8c
Jxvp+r9nrLLtO+JvXBNCFFiFSJspIRdUbbhpfgEzgM+9NcCbE9iIbfGksKblhXcOvbYs7Ozvo6TR
zja6ceVA1PjaTGWSIsB6vHF5QKJ/HtxbcYbBJ4cZ/5vqPBMaJHSH0CNvIKKpu8ZnQ/GsmR6oljYb
mbP4tjXx5FiVadKqM/qhH3SXOyFj3GpOmTJ9bwBSbgAMntgqGT25Y8GtGqotqkpfC+Pff/AFtDTg
iTkq/otvyzGDGPV+qMd4xWvbt8ViYs9oIiHJhBx+fhti4OCTS5JO3dur3PilsTDnOad3qBHAnppU
qZhaysHXmqEfRJhPqjm+YZ39a4wOXStlTeepUI+3ftMas21RxspxG0jxYU/iqiErx31hnIcEP7GN
Cg1fWjpENdsLx7y3W9Vw317ftwVvbjnwSAbN19NO5MnZuHHuju27fWKKXlw9+jpGLKmVYx8dRRmX
pPPyhB4uYJ2huVTyBdRBgkIe5axG+4b4VUjUJVhX2ZuT9J37cEM8LWIdmgXdacYeTc/+OH61sHww
j+J80XGgdobUAWlWDa1ZlMKv2nX/80sGFQgjuagrycPP11bhQfj8h0xRH+3MoAXThMnW17/9hSnu
Ud3GfH1QlWefkWU/NrWCAPaxJN2PANL9mx/ZGg3dVxYSuui3F/VQyuqoJ96sC1JqXaAMwOymt6C2
2OS7bSL0ureFeuFUoMV4GMormJFnYyGFjmj2mBW7a3shlU+IzbSSWpfeBhRA31unG80EBDWJJBMU
eG7G2rkgjYhaOHdmYBPI7TerPKvXWUTcC+5momVr4G/OsUgMxWnVlUlhbn+R5sSnmiHEjctQOTbo
6ZffcYKYxazPqSfMHcOL2ZFhD8+9ST3SEcz6OA+kG11DupQDymf6/L0aEm6Bx4zzkSBV7g82GPY+
xYfAryi+Ah4wIVrvN18OSNZN3/BDkCBV0y/MeCLD3CKCTo4HeJYrNUaQwuCZITe8uGWT2x6ZvWmg
YbuphsJqIxqx3bPDEQHxJaSW9kMVdWpaTfJd43p1KT2Ks6/fnqZkZ7UQvpvZpuB7gW6FPLeOdu6w
JgDW/Akir6D/VQg/inDthBT5PnCYDxUh8btkP1xpokFSVUuf1BUk5NtUExr/yQ1cMYaeZbiDSz3B
D5hpWF1I2NVClIag/c+Po8MYSdx0jRIZjgwECzekoHfQV1iIEev9vBFGP4xBXD73cmLsJ08jR0tM
3V6zNfMe79BTi187NenrfKEdly398s1FVkSMtN22/J2KJMzY5EtvR4ibwAxhBGaPI51keMUucuVr
ZP+eQhupn7k10x4Hzktc/ByKBU/lSFTZGMoxunEPCOYvfo/giOxBDBm3aPfYZPGHpe6cQSRUYZ7F
779Msw+U6GXFpi0/1/B8st6/62H8C5H0DSAbaHhnB0gRjcihoUY6BLn92cU5S/wSMmKqu0Bv+itG
ClLNeFsshzs8vuA3tIdEqYohcSFOQKRs0DeNCYPTjX0NfXXBnST6BThDQwicgWFc1Ny8uSdePKi+
/uvuhFKi4VTYbaIAmoAEqkpZYe5Exffb4DLGIePJd2gtAJeuEshAz20h5iFPkD+edkzbmIQR60BC
AZBLhGdUMo/pyf2f09Za8OYTbfzArakFnmUBwzQ8U/8ldsaoZXaSFyNoJlNbcvh7jStgU1H7UPw4
RrWwjmC0buB1jYywZPSKtLx26XZcvxd+Otmj0C+Ax3nsh0dEvcDe1H2GEP4DbetwjJNcDms4NrFp
aVPIfYYpdrXe3ELVL/5tigYPlCachj4wIgSPqGau4QHIvtR7eS4H3wUWniLpFMHx4/ZPWm/eZ757
dxj55QXexAsdD3ar7f9YzLbDXR//A2S3PSSbwsW9W0kll3+MqIgUmeEn8LNvCJmJNDAPXPG0YQbs
x6dJUVtUWW9K+9jI8kcuY6EGiYTomFYMdAKvEyLSe/6oPJ8lx+60nDl2O753LaEqKzcWhHiL1AYZ
GxfqXjNB7Iu7r2DV9KBAEnMpUENBLOIYb8UDQQ2j083UEP0lwp5qh3dFGUr/NCB4za1r5IQL1kZA
1koKcA+AX+iey483u/SCURsPoS4BlAOaRfZsC+SjF2ijCQTmZ5J3UoPR4+JFgwAcfNs6AT1nfoDR
yXJ9u6JzWcrrKp4PNXVw/ikjDYl9ROs9Zu3KPsNukfc+66rNF2ql1Q/0cvlSYUbzvblAUClgMH5B
Glpj/xC1ZOpT6VIV3hakquw/BQQicH4HsfIvN+u2soR/NY9EJ7hr/mDe+wiDsn6x5VPHcjW/u9+p
FAkM/9Tq2hvY7wQRfCPMOwptLK80MTIp5QVU/a50E2mHzG6DqAo4EbXM4/RdySXVDzWbVv59leBO
aVrOl9l1xIxIi8hJbxHMQ093ARwcUeSq0eZwW6B9eXnu5XBWBx9LMVySsIcuOi77Ta0HKXqRi7hj
GRpgzqoYoAyO5MBNiq0h8kW6WENFkpWib72ZeQYjXCIbq0Gk/fbg4LDN/5RnaXJed+Bluga5jYvC
hs6qVuugS5QqrFAB/o+b8Wipvgm8mmLR9xTSj6rUNf1GIH5DuXNZ5raToibGZ8bYS9AQd15wRXpk
r2mUcXci647w6GV34ZG0joO2kwMzZwQBcCDWSjl8nRWa36xzjuj8b4mKqLdCUdgylpogVzIMutQv
sPOqcLNXonTpo9KDqZzOG6akqnnGtYQoDP1xLlqeV9MMm7HZUto2SzhFbWGEqHoUza66sGFiVDjx
vZP9m1TAGSQHVupj577cv7r1SdGpQ35+zzAE52Gqi5i9OQvF5hL69RE9leMAJASlIvWfqm5YS2A1
WRNZWHB5UOYpQVtyOXohVqtHj2V+7Cnr4iFR/z8cpbz/xyX8k5Vd56UAv1h/piQrg6FAY6XTNn9R
ZFMQUiuupDaIdT2vI+N9C2kSd3B5emGSr64KHjPIYRRCcZjMN/MrLSxnbNuCs335EcxSbM/wf5ps
q6l+CbO9A3QurmeiKSFJSqoc6xADNgVXXwSKHoWbRWrI0Ulxi4+6o9Kv0nGr5mroqDegGMsvvszP
FaEo+ta2gPpaA7qs1IQ5aWZNF0rC4jqlO6wJ/Uehpzx0keGrnQrnqZypZncK70tB47DvKawiGwGv
AOlBCcdLwbBFX9lpivwQvm88Az+9JQjO8beh62AbgMImXxdJgWxpQEFMz2zjOiPC2UwnO6J8EfNE
ozixhb5AIV+1cXVoOcTAOGfOH33ac838vrrlIQPH+28mly6rYCRqd3Kgx/zOrcqyXl+rSAUtov9l
UYQvrpGzxDB6tUD1XwGl3wmq3sup+VTwEUCyeQr/m5BxXZWKRj2exeGC1H/8BCTgldNHI6TnKP4K
dOco+llXwhWGU6V4nEhekoe6+zNhKY4mSEZU9gv9+dowLyllReJf1LPrJGy4AgDuAHma9syem0gB
kZRKODr8o7itgrfRH/EOS1fuum7vX9GF4JWEXRTcuOEIRSk2S8PdmBteZrwXpiDv3IPYQ+vTVxUz
BX4BDuKLLRWAnlA9lomEjMVdK+dagInKMgH3ghWd+8fz0YOaOR4Fh14z2TlhUqzT/3OcHn8e7IZS
yp/2rl3M6pLLXVDfBxQ+d4uDb67/C787EFXFvxAAFmrJ3i0nUeDsJLIg54CY0vVhXv92F0FPSYV6
tXj16JQbcNXO+QaGYSUg69b3TImtv5H51rtGcfOs2/+eJ460X9D24ooIW0OR97Byc52z/fC5MlAP
ilQbJWnlO+STCmSCDxxZ1XgFBBtdXm37pnMMl3aLp15vORvpIiwxIYObPf6FSIY/7IeJil+0zkH4
6glQB1qeB9iL9wUoKos71xqY+0/VvkKjMDwwQeNp/NsgOrx6YziVd2E3DmMOjz3s6XJWzzhxsSDQ
KkDUfchLV9p4P/L4pacKM8gR5wgPfs1Y8LuoPw25YhV5rnK3E2X1Nuxo1/VGi71v02fGcwqbK4mq
27m7sByLUl1K7+zhmKaAg1tPVjXkPKq1G/DbPNTg1M25bNaGu02zaSjN6+AgAT672qRaPgeezIX4
HQN0momYbmMAzfAG9vurn/xmClI9QPFl6ReRiQT0x8k/w/jpySi+Jxxu9uRLYvpgzOITbt9om8zH
qMAmQ/HG2M2Lb2OLqLDLozqMmFR9o+t3ey5vu2teosGxhL6K8/bod09HEW4btGWRDZOwY410rJS4
P4Saf5/xK07GbjujD9od4RE8ssR1aVgYVOSWrIWLFcx4x9ElX+tOx9VSnaWGeX9C3iqTA1ICblxl
9OM3u9tctH7jyGU+9WAJR877Wjge57dDK2tDqGuZgN1+eEytPqIE1qS1H0J94exAUmncuW3SlMAl
iZCFQViThso7Vh1jtmpXV0vWtaOtny6AvEiP3Kdmd383W36J0YRsLHU/Ubtn0w2mEf8ib5bvUyzw
l8O9MzIlX5GbfW3JT/qUCM0+9X4RRWoBi4GiJV1jPudS+tOtsE0ZLHHMk7l8piK4ne/qOwrsGJth
U2nvbeIs5z8ETNE4H3ZZFEfFbP/mfR4lMoxfSSQJo3mUcZfQD0XhP5A4T9KAkKwPr5CHrM08vN4/
xJZ8K1YUhiYrVOB9YNDfdmhfVsBxNMs2MbG6IdgnmjCEGYkVslN0KVsjt+ljZQtzy329TKhZoxvz
ueg7vgjBQMWeIcDD5YzDw1UwCL/HEBuxtnfpq5KZ0xDH+WOUQ05Gj+at+YkyS4b33Zrbps4ULLCl
ZjmGc75/j3NH/waWRwZvu8SPiSkwaoSRKH+T2SL7ojxZ08e1RJE3I5g6J3dp2KcgkJ32RPs5Vum2
HRAnNuOk1y0IF336u3dneCLdYGe0vX9Z2YOotqhHcvLGOfFs94gPH+3XSgpbdExHkuGXUsxrRiKu
g07PaQaE5vMRpyIUFYhhvLNthIxDeS3TQiJU8FeQnuaSiUAZpo/kS/wTlsATkySl96QrrhpN5waR
CRxaRnFu8do7pWydF2nuROlwExHKbcpaINtUi6u6EXk7E+UOpF2xx0hNQhlmczsmy5wGjFAMepFN
acuddju/f7rCT4zm/84UklhanC3HccZy+SsKNxw/UdlpDicFPV/MLNYO1lGdjWRIidEX7FSzq4iX
jzEvZKxv683QoyvC4i8JF/VjlCk09G9b3i/Ca3m1VFbTVumVvohUcdxMaO7X11PkgnT7mQDZkThR
v9E2Q4nd6qSddiRMLErMKrB1Ab5No1YBrEY7itVoEDKFDXdgmACAIu3vV5Lgn+IP3ERis/j8mUtq
zEfhxH0oXcwX2vic8xI3H34OoGLe256rlj9I2u3mMtOeJhcal5WqX/e1pj6VHaHCU1DBR86SiuXH
p1aRKqGyQV8ALnnhWR5KWmPzAnOFlaxtjiabIYydd/7Q1wwhLgGRgbSYs1vmq7fCQEiGc0L92X6a
XaCdwqYSRZ5G8yefzeN8Xf131kperdcCBwFURVyZjNEVfcFVCzy5i9jf83GNfAtVMNPgBEH/wcM5
CIQfPalitvXXJncnW8YKBbvyDpXJuCD2FsXTxOFOVKvgiU+y5GSm1JR5Z8Q/atWg1vNxx73rDoct
hesyr2mRNV3+DOMWozmBjg3zuPRJs3Ekx4/MQz+miv87GoRMlBjtHO2XhuKPjKRPjuaetXBq/t/C
CIuvkbP/U1bwpDIDAYWbY8Zhxo1GA52/P2CVwBrUr4HyU2ZpaU0NxAYSPFE1RR6goNVq5OOJeJbf
jB295bPGrrOlu96gHiBi7BA0OP3fhOWcAqmzNNx57VOWhIyQzpG3Dc9oEfU7q6EoPgWroWJ0ackV
7AA3zhrhv2N2IdoET6dbfzt6sHDgqjAHbio3p6eV8tC0371RB8c/G8Izc2v9pFcWzdGiotK2kLhJ
n/+zARWmouQXYRolJhiIws0JmmgK++NKG5CCPIXQpTRwICbwqpHhEiB4m5+phErZ0gDTrJa5TKNF
Muatml8trBp3aSzl4kh5xZcoQC5wo80VxTI0nTEKgLHDkLSJek2Z0yEhu38/WJayE0cFvWCivLra
niGi4wIHkeftA4kuBQ30Jqsm1GA6bxETvEzEoc/X/z8tQh55ZKaLsBn6jP7TlwNr6t2eBVRfCMg5
6en8bMahahbZdHJJWqKX0jLFStBcUpT8yO+OSunyGP4zyRaA4eFSfrcOYGO2SoVr9zLqMc3VHFJi
tYGn4Rsxxz/6ewQGMAiw4oxls171ajjZ4IAA5Ly8QTLVWzC9ixFhOEY+AA4SSYZeaTMpIjozsfAq
EdjL2+/z0Pram7pmi2BEQ6ArAG0PhvaK1fWm7Hfwm07NiEx5ze5QPY+gxdQTrTO1N2rIT4P5INh0
YqfuU98iQwyHmQmsPd4ggUs0Env3PPUKi1YGvTlJQNFPe69nwSgBBV60Zua/DD13HFPx5NaasYbI
LkaQ3gm8FYxKd5YRiSU9qOZYSjNJJt1156gTNSi0DA047RVONzXX/xyfDpYw1kNmqqVK6zTeWSRA
bdW/5Vv0HOeV6pyznPWJj5juG05cNdOvaId0sAIYPW+iymuqoIpo7ctEVUuaJZxsBTqLjdhNZoAW
YaTdiwAosk8ab4w0kBQmLDIqQf2iWbOLBh1W27eP36sDfulLVY4KSwmsoRmsT46mzXaLIm+JQkUa
zMbaM2lFZUyl4Gty1unRaMCKEKbms3whTSubfq2vNLWP/NFz/4YJnUaMJzqm2h/MrkO5ITZfd+Oi
TCFw7IW3h29WRJDTV7CZui6GOWWsf/s3IFENst5MTSYDA/m0NC6IX6Yl9lSlFNzksIU92jIqyFjD
i2xA3zie8Cxrhi77wzAYnvlpf9S57QXCXF2PmaM/cbE43Zjs5+wLyzlm2mF/zMJvhWQd+iOMTrs4
d2Cj+H7SExaHtntVL6PPZtEYttr2Ko2t6Z/sEl2N740G23sKcZgWb5CEtYbZK27bBag6hiNDZwsi
j6R34h0Z9zC6R2eFybASEOoYjH5pTzPET0FIiMT4L9wIP9yLt9dh8aDQmHWWgmv2JUrft64wdtzX
yisvBASLdMUtH4vXbiRmKT27LpZ1L1W16EX3+uZP2H6U7Vl50MGYQw11jT3cIQ97Y5ShL6AJEQCT
Dvtr9IC4jcPXjnrPM2QnwulmuK4sAQrHlFkIWlWO1Sy1+CFr8FuB1EH00k2kAM9xCYZw8M+J6E7A
cURrF5nc78udepaDRRuRZa7Zk147tFNuY3AEzx9IZ39yyS+gA5TBYV5LqkG/LOU/kv4TU13kcLR8
ancN659T1LzVEGUDmo+tzqnyJc+gDoc/l8zk3KOykYb7qn9Iv2kBWGZ6RV2555uWOv1ndjkPEfil
QyZY6fj2gK+hTR4XWmAdyBDKKImfKhHh2YCYiu/mj1lHepam800/YkBSwc/o9uUvg10IGYoHMmJZ
deJvKvu1VQKb9snPB6BPZzS4+a9lBOG6xhts8tGHDIZDfekcArPnvSqax9bK8q3AiItEHJmT+sNy
jIyTKxs67UjV4aZsA3316t1KcxRtY5NPajaTafQKor+v+0CaQFvIUuAS3bJopn37dsXmDyB4mOUj
RJFU6YVb7ZTuhC5Urm8++5iuZIG/OCz+JFERuEIgWm5Qy8OkY4+5cAMXOScZfciBegd2JrvdJQU3
lhV3l2Yzx3I8Hu5JYsbCcCVjwIon+BXm6PyKee2Kun34wa/sjcFc4biVJk8FGrwe4AeHXV8npQ44
/9LartbS5ZXiiD5QkowP2iXZTcCBHqPBR9fQ8aRW2j419HIpF3xiofEcQIuGDNkrfk9JU3hcTPaC
H6ltBNzJzkG2hs0WAYEd/Bni5RwFxUlJDfDhiRtqHd64cTVn6r+Mk1ZquVdSn2EdtiEITfOyC82v
pHnRaDcOPCbp3yCb00fjFh2NqmiR4Vtqyk+s2/871+CZC8FNqBjbqI3fNJ+SbYgR98QEP2FoNpxY
hAt32lhI8KHKYnVXxVRNpF91mQaYGYysz2pPnozCQ/HURiZknndNDYLp7w+IUHdMMei3hqEhgsmz
LH19nObR3Hkj9AZR2YXk3F5l9R6RkTspfD3bdlAS/UqI/DWH0eWoyCtelC7NhRmiR1RcOdkuDTVJ
tYDKOgNY1a9UNYa+7tlHyaAUgTIPcOAqiCT+6FrcHin4Xp4lYOYxow9CL+geQ0hufUEKdgx+AVxU
0TLrkEQdxaHcnBxdQ3adlIVtK0PaK48ODWUsHkamJF4+oXhz/yVqggFUUOtpnTv85o91a902FNLI
jb9Q/SEPzJsH5SR+9++h5lRZHpKjPvM272+hMQDY99/67vlalG60PFu+gxPUa3OC7yUxmGkM0Dcw
WsM3plfmqZNt+N33VjM2O/7LKm7QXGZgCFH80PLifojxzvzsjZPgM7c3LWtzKOBC4uFAMuNKYZfv
T41wihoZTKkrWo99Ip1BtXvNQ1bp4/bwmw43K7n782XZCB/bXps6HNvxYYYxGWm5S+4A43X3IMhe
INeuODVJSt8RR8d6YYwiQAMrgk844fVK3fTuBWQwVYbPDFnlX9VunbNmMM6twq/qOWOEDkj+Gxb8
kdcFmex47MhJNd7kJgjmLlGmq9D5AeexLQMcYAB5OSZgqHr4Sr3tGa+uuXkTFr9KgdkjfgCxTiVk
FC2zFL0nHliNokPz8OKRmls1pCxTlYLfx3NZC33lopAL9FjJSFKyiZVksytoZmK/6PDi+y0z4Lbh
KhviG4Ms+wjiypiZwB1jLCdW5ahzwgMhrg6ah/U9qxMuVBG6NFx0G6EWxz8FyueP7OccbtEDKvGt
+j5a5Z69oWZsrhi4CUQC+uIBcc8SDb4o56Q01jhPSuEa6wmHyXyKJ1hsCrjzfDO5GeJBE1iZ7obR
4UGi+exwmNH1+bAzH8vV6r5KX7jFaiWoBjTiScWbXxFaA03ArTSR3OVKGls/0w6E4hNh3Nie+Jsh
F/yjmkdot5NSVNJ/1kwWnsbLU/8PfbjOFCehss3boHXb+iWcSYFeq1qhQck84OC6D807EeXrHbLU
SsNKODVRT5gjVPrRYls/iGpFzJWe+VGimRkm8awSXgOvldyyfHmHtKMqTGItb9fKMmGs8CUUkXqc
Sp9J5G6PcRb5+6ct/IZAnf7aPjrYvhN9JoelWwihe4puzSkJEgwAWDhdzn/A+bjc52cMstsx5g2x
z4tafRezEvHYT18O0Lt4gLfYrQlKVtIGQDH+LKKRsLCIyrWdCyMCa1lHK1PnORb0meuyQceNlqfv
KbxNldsQnfrPlqY5K4JLt6sPJwBQee4MidFwreC8Zp5sL4Gze/boHvY3/hkIv/OV2tfdGylOpfTQ
HqGBhXke3BccbP3F7KJAWpTiwlnR5O0ZjP8FOK4AkUsQpQeGYFkWme44nHEvq2WAxnLfk3gH7Mdy
4V0cu/MCY6cZNBQaPmHAS/nqYktJCzrxaMB7WE9h2R/Bv4g7f9pCV4GdF0n5DkBcftEV0YkrWy+d
y/CFvaBucI9LpMoWAY3eMR/17vM/Lro8NATFIbRDiILqNZfDT+/Rc8jLObQHMWtwTwlyYh92R9K5
3CCzDA25qIVjmFJgw9nHn1M1vrgfOnO/8zDGLM8EYmV3cx5mqGfg0W83FQbVU+o7gCm/uP40nVfN
EeRIUrAYhd5j6yO35r6SnnA2GcO5qHFxoBVr+wcCB16VwfxJmLhuVt1coDfGf6qrEtfDc+21fNbQ
BeT6PpUld19qnPFDSdASF5PXGi3AgJzjyib2uxj2BuXiP2z1WlNxkVWC2CQfuXNLw2YSF9CWu/vF
PkEGsU1RP0Pbu0FAaRc6hAadwAC058JM2CQ90c0/XYWnl2l5hezjaRVLyhplMXI1MoiokQFOTmoF
xddolTs5DIcOXOIdng5OkSCrZulAHzuxQT+IQWrUgCEwY/qp3VF4E6nHEwHQPD4q7zbK6vrCPQeb
HOkKxe4BUb2556pLQPEwvcd5eM9sKlkAkWPRerrCFwSVcDFFlfcwS7ClnHSGaF6wOdwynKpI7QLn
uxWX2pRDjQxxq6wdS+ftWw4/CBA7yBM1j2iAy5xMF0O7Bjx8sKXXZN+zytjEBkPX9n4MqYhnlFmq
vqJl0Hha3Ak0CAUh5g+45pnyjsdzatCxxskgvQLFoDb8Rfw3CEdKdzy1vHku2xSJE55LvGBjZ+ch
ioIE0dujsuLQIo2c235am7XZAwFLNr4eVfy88imGIJ7Ln5JfQ48RHyC6i8KGsiA6i2CM6r+eUAXW
AteSJhEhVE1Grsg38mrTMzInGA6D1z40RX7YfCZPnI7zfVjaqljQ1Dlr+iec9fXmkf2hMudA+H5E
hVeHNr1/JzJcgxwXRRGCUNFa3cdPVDc+zcHA9nQi77yYk5b0BU62GR73/nZQgwlERi44yNxHruz0
m6+n1XXCqpL5mESBWTS/DwUSRtlDLAm60kbKyPPnKp+LbH87Wet960FqQFH/PMZvsXSNBl/gCmlC
QNqB64Zb3qw6okAkTgznDLSNNkc98RdMgJAXEpXHUASaLh7uhoJhMNGFjrUv6l9+1UDpy41iDKTU
qwfJcw2cYULDkYQPsUsODmxAcq+HaqH5XTtLxWjCTBK8hVlI/U6ipk1v+X13tH45mT7neYeDmalQ
I2YByBRU62ymrwlR27Y47Wy6wIY4twXPpy+YR2WqgiscWYqixNMwl6s0MDVFD7r9U9r6khttou55
WC0HWAAQWKxUkDx4+5dkXu0qrh03Vtda8u18XwDZB7ceqdjOaTd5t94kU4S/Jk6QL9jWOWvmlgeg
9SwKt9dGkyAkhP9KIsCx+BGPTNNzMacpiR7OgXDxADo7b0Gctaw5857vH7hmzWVYQM5daIy39Ccv
C/mCZvMKN2UwqvW3vDJa8IBxRd0XC0Ly7LEb8jptAJeXBYaXWe/ujyzhqUFYFnWuuekSmvKaQLMN
485A1cI2qdB/NrePoJouQrKyX1RJdEkk51p4jw2zYeA3YDcSGCiCFAQLc7nyWg2340qu49dN3tWd
cZzv4vvouLcrPlPjHZeIB1RQipanXMivXeXbZCkdaunOjp9gJAEHdPPTXWGtniaTK5CocUz6uOMV
5ErO0THud5wgWs4Ml4GCrzkIP+VrXgxo1wFgWP9lylWEtjLZ6TFAIrJ7LHy9ZqOuXG8fPvdXmPp3
TGvZ+kAq4AUebimofQU7G8pEpN+wV06i03eEAdIaxPSaWa8P+FSnbDwumkczdTXefVnquXaTWOT9
/zLn1AsXxC8q3ATOa5SODVEAqIUjsgq2X6+cTq6lTBbrnIiPHkNRPg+xknglMdEWzUSMeIYQVIbH
yR+ldWszMdISGT3i4WUOHDS2IJYnQZAzFTSnkrlWoXHRn488oG5buuBEbEG4pAm8RAOzWvV+r7O9
1bAW771V4uQDRkE5pMGqWajJm6mJcYwSsu5N9AfhDSeshmxGJiKTRyE3ILcm4pWZKOdhFTrHjG8K
aqfYSL6phkiuLf7LCXrmVgmNa0H3Aq1DoWUlqebO5fi6KyVpeNLJocAImgbQCtMxtsIGYsYubgWW
6lxuLcT25GiM1jnKS1exK96X0Iee0Iy+zAe4ZRIcadMheA0YuLeXs4QsSlSOeQ1Ec7JFet6HuFms
r4sv5z341O8t7JMeC2AY/5ZfugiNCS0eVS07rMldmkwBwW1JnScKtjhq5dXsR5lrMXPjE+w98e7p
khQtAnsKlCuCQxRThNnkJu7lry6IvdqhbzrmuE//bHtKolbn/uNRKocC2tG1MZ2Fm0YiQyoYzdaq
ffUag0YgdonUvRvYreSgtD0Yj3nO03WYErMBHHfVdnDFeNR7hMjXfncM15EatHIOzUldQKcaB+tr
5Mmpmm1gFyzSbhSYT8N+F+5wA5hacYYLap1cInO1LMqUSCX+wMJzKxROyoK1GDHaRzitY3F/Km++
/R8UQ+BmoGJTphSeUFX6IuHFUO7ShwyVCbXsLLO7UXFYmkfijwKPiFBkjOYdAxY8HBIW5NQe+Who
R8LMPm3BPgIrYcse3BJRj9w59jDV2AwwKGQD7KUZvi9tQz/56rUfzx4ZvxbsigaGKcFREZiyZspk
Si9xBK9By129s8qoFXc+GfpSrEc0wAhNfMuM2pwwX0SZ3g1ocMXQ8EZTan9fE5zMMcE/FfUUFW4Z
M/4xuL/5oXjA4TD6vUqwQnnwSuX1xJeUhCgzjt8224pK1fY7IElvUefi1bl9hUTGlqgnfkGWjVnM
hTQ1rmPSOfMy82pmBJnZpp3EfYBLwTdZ+dRfllrsdQ9edRo9nfcSEeMu8mI+q4ZXNdkG8RoodUqZ
3DVW5mfmNoO3s3c+oOPYkvuWriFWcsb4p5nLbrEkwjB/VC4JYIcIP5r/34gJPrkOyOe4xtybD6ut
iumciCQ2HDDf5V85RKGKlU7Nm1Muvb7KCG/S1nWP3BUyaoXUpVFLfwoVDydNddGlizTkc090UvLW
au5w02DvyUU632trKYGkjrzwJRJy5/UAtEpvU0ULWz9p4acqS8bl788Gz7DONiZmnjRNYXCa1ZFg
MpnvbgD57GqfHvKxtcwLWJyPbO57OASITavBATUqoO+JX/9jjYKHMEgwVs0qRhbUYpLUq4dwu1m1
JiSaunn4jiM9SZYkJrohncptpAfDdu30MbXucNQvVQb284qQFuQk4wxGlvsDtkVJSbxGBmA8z0j2
RJWTBmodaazcn/tnpKdQUZqs19UqnpZ/twLVHJ6fecIpe1xQazkJZ9m8eU37B2HaYxazDnXY1HJ7
iJOGd9TqQnSZnUpVagThe49y3MBAZttTBbST4CCTL7ZQ/FebBKJGRTpSXFQN86Rym81uzQkQFMBM
ZzapsMNP1WhsIf0jxdh/aDMC5lFEhzpQzXwEQF4/bQ+1EqgxphgHO6x/LQTA0VwS4Ozn/AZyrsd2
vWZksSCCwBaqVZIaDFd6DxTR7sY27rbBiVFqBoKLtySfGxySVXqwis+zPcMVFCdZBpD91Xc1Ova5
Gn+ABhq051G9YyovkVn3HFD5Gk1RV/VIRImybiCDMvCzZ5gQyxVZ0Uctb3vapwcRK6sOxGVI2fSK
+So6WopvEwbv3ULCmfHkDQedBFtGp15lOjuXZrmPVdozNlJs/sKdVLMFT7h+nvuAXBx+F8bhMeN2
0YYSOisycY5TS+m1YN/q/Fdw0l+DndsR+pilT2RdvFOQ10dIdu9LEHuhRxw0b/9A6TeuJjBgeNkQ
CJpt1eSzHCJYm9rWF18m8iffZrdrzfpwfDKjnvX1dn5mepG8d4ouwNud1z9TkJ3Uc/CI9cDEn70K
cj3ULxmnMUZ6uOVz2sI2w4HJZxW/Zz7sbz1XLMgc4x+janOUAUQiCoWHRf2kvPHAdkOPMDxBWa+m
t3qtkLKLQZPBtprjeYezBb65nEEh0JGODTIG3z0UrW1WTuxxbXSiWGnIy+qf9zf/9oSV3s+yHBxd
HzOsW3E/r4izOKQiyvbDcu7U/WPPjJOYS7wty2eFALsghndQL5WYqXUwXUiO7p8ZwsTkCVNETyK9
cj+bF5oeDqyVP+P/HLTk7HUDlVmYUvSXBwWRlA4fkC/JkAfqjWhft3+TPyp7OGQ69vwxK7bqulhG
qf7J0/TjsalaIKz83EsseKROQeiieSXvkrh7ptCSYB/QKoi02YZ12vnAGgbwQIvk2gyOx0DD8wvH
1fL2+g6ICF5mDpcUeoSjwd54q07FwBaSMtBbntk9Sz08QlnT6X37WWOQksLhmlpZFXinmj8dqHia
UIIjv03fMDl1xRuOIa+Roc3jy3T3vvE72DMjretdF6dnLnWhra4U6GHjnb790jYSb6CLxzRfuaRd
RMVIBbVvrRf2WEUXt3Mc1oFcB2tpRJdxO2pTHcn6RqlgUl9CxFSpvpnsCbdifD3/BKvO0RzVOFCK
wJQxUpTTV5XulZJz1TPUhTTIxneNvYE7pD3RF6Y4Q69zjkamRLJjsIJxDoAVndEU5njyxRyZnkXc
FmKneVSYmq/G346ZiNRScVIBwmjIWuMR4w3yiqYWE2dbDfvXUfoOtfUMQmBEfY3V54EWR4HdrFOA
Kod2hjcd4yv7vTHUR5WZMZMrUoOvaLiKL+Bzi1Vl0GKZoRu+KLOn+fHW1J1z5ZghubKPcmtrOaDK
VvRAuJqXZZsnPtIw+PUokMFRznkMtDJZ8Uin/DncrO5/GXKrswWqBbwrDKSc293j/JSzmu7N/c7D
d5cnZj3YqaK2y7qKMQ9CA9OVj+ZioEnjesRSIXGfik8Z56stJjO9gI3sQ5hxyopZTOaAmpMHArbA
UAZuNobuounU5CjjXPgOQX2WZY/UudoCVGTDaKkaBqJS+uavkDDCGrI8xQTy+OkqR1/erSWHVqaI
VNYdvfvqnL+y0Q3lBnqb2tFM3Y6JJ3HCZmNoBy/Enn2FnHxOKhDwL8VGCrr5aO0t/UVoY9fbv3Mu
r2dnPYjS+gCHSxyHN+oUBePnEXaE8A5SDvSUCY5NUPs4KahNEBDD+aDWDihNmepk4uVKOlymyJSs
NUHQiZndY3hMPlBwFtpl9oMTEQO0sRDl+TfiTHpothUJqBu8Ukr7f/9H+ORLPowup3RbUWYkLZrf
Gdjia/Ml8rYV1by5w4kgWlkecr+R8FkL4uaINqXkTwI89C2Mn5NmxGL9DW5Xap0oSRlgoOUnHA4X
lUE5EtWGrWD9tdCzEzyRVG4YuDE0WA2yH1x+ZGgkT3MGymVKl+e3YKifNGxOvdkBF1HFGXOO4yUh
FsBY7qkF/oLlHkelXwA3Ev95QjQ3BggEQBC3iUjIIX+HKIFYiEymui58KM+1oBKqfHYJ1vl/hjgX
toLETv2d83ZHbu4KkfURcexhsjgXraLTKVRpD6qyQSus46pUBdlE2o7F17Ya+wRtRd+fsMHFJO1A
kfdyjH/mlkGtg7tzYBDYWd7J+p00BOVUfYlPEUBKGy1gQwBZjrN3dBZW+73lXZMcMh9OkjXvyx8s
kFjPKhnr8+fclHDrrP8pFaovvfTBF88Md6yRYxGiKFag5vRDE+qx1DD7E299BaVp4b8dRh/yOHC9
4swbP6f8FwmryTwiK9u+Tixd4UlWp9UZyMey2A/0LIX452UgfcZJXaijbPPFtlfkGgH2T8d1kRqU
WOPjzxlVoz9eU8luqCHa1KyisKo2uoQLX3tVOM/wL6ORKcuhNcVqksMyHfc4ipUdBQKHtweUguXg
/ZcZd5yGH5g7Wz+EddXs+4PUhOmdV0uyzcYLhY8sNlibWk583FFWS/X9+5XMvs9uLpyMxPgXru6/
EoM1omBuEXe7/jnS8kL4VgeusEFb8AGNYHtHFYMI0BPN6iOJ6mMS4ckTQRqJrqj9QHJ9YR4BZace
sUaRQzu5HiqW4LId7kmGjF2ikMsU6Tbet2XqFb6j4lOJMjUMmEogXEqBtQzxP0OwtsXpm/+UYyyJ
Qwpvaaztq1KYE/mzrySyCl7i/nMNGOe2JYFkyD+bcNB7X65PmUE5qa95EoDiHnVAxAWcr31sEo/S
Z1ae6cD7x+aBXDVZYsohDmX5sVt42w6nxng8knX64tTvT4FBMlxIKNYEiQJP9ksr/sjb6lvvdL64
cvJInLSjJaOxPwz7wIlnNh+37RJONrxTcHBs7jCwVx1E840xw1P8JSe7IS3ihmTshppKC6gL6sYT
1ED3gv6wR/SqZJpbjFiWNxfbDfu5YOblSUmRvIrh1H2I3SWv7+O/Ehjl1X4Z9krLgo9n2Hwvw9bj
5XODbUhRIgfdK31kOIBgFHBEmtX1Ux9oBiMj2cs2oKgzFABcXRXSg4YmOijcON9N8S0oz7JPs3EE
h7/f4Sm4T2i8GPMVf0n52/G9Mfm683pjwHEDZ6Z+xp0R8wD9Ns/9xvpDcCMiGT+dAc6d0KhcDF8G
RNZEC/0dhVpLzYCwnZ2oylgayZcqRnI8mS39vuWnEqutLkdRsz1r8/vQb3pLtf2RUxxy5PjY15Iz
TW3JJ0M0hF2U3UtN3FrGZDOz/jWQkH8hs6ZPF5gGVRKdiFIVAr93cKcr9PvoQ8+MbGQ9RTISnMNq
BUQgh4SzYMe/2vbGIeKniVv85q2WYediN+E/MB0KlMwsZjSgy46SOApGt62JB+cXDE38Yh3cFIiS
I7YHjcV52S1NLkd7C0Ek9JA/bkXj8FJO1CnyOI00o2pJmUG4SZINpjMqlv7zkij01bvPM3vqgAsg
FvFLgrAKF4/D9DrkCeaCnkz+KReEUX0lDNu6uAU84e2ZfjtrMCf+d3VNymtH5K+YhBzbwcH+/Fx+
uIPBjb1QY+uq2CBkXJH5+XTKRKoB983NdfL4vn+/0PlL0NOCngcr8j2f/RM/gZMYEBp1sKX7Qs3s
Ls3mxBEAgd3TKMjUBg91NzomtR4f5oe/yiwNDqD7AxTQV0MoZYhAUzIKNqeZicbvWKWcdl/n3NvT
u+zCisocUPRLPHqMqUZY4c/wdF2UxMoJEf2mbUIz+DTWbCn0Eh2rG9GS7qnFr1DouneutZH53EcG
PStZ5n2wZwEsfYXF55AptXtRj+YZDHoHQhOlaqq96nYx6VmtxqmQRdqTJPKT0XHZkE1h/ZEAt01o
OTtBb/cuZJJW+QbaNWE3FSzWiOyhQLU0Sx8WpcZd+7WkC/0kd3SWjW0njwkDyjxUDPg1mo7iykoR
26NLcUqq5DRwvCPkvRI3hfJaBMS6QHx2OTtT04ATJd6SBm6keRxraxe7lDg4VwZOM7QVFFNho1U/
wpW3ItCFl6EQ4rsAROmngKXgR5kHQGZbl5s3G+8FC0OoqsvqljRPYNSkMlkjsi1C4UAjuMrFZr9K
FWmxzMlD8eJOjpekxjeLv1mFKWgauKaMID8AIL7xd7FCEcUhOx5R/t8Er+jDbgeIQdlnSyWeU8hH
Rj6EPFt3XDH04DGD0tm9lIovx3wLJcFGX3WGUbRVIJgqxC7cmg9TWBppgsdqghO3XcBlmpE07Lhn
7j2aBmFGuulm3EAusFG4pZapymkOl4R6qEfYh/GykZqlG9sXqGaHqWLgc9KEvTxABi+3Y9Myz3Nt
tecFCFbb8aQ5xBUx1uosKjATnPlie68pQCOWyY+d+ohk+Q+dFiObjn8xm8VPovfkWHIsgeZ8Eu2a
F6e+xcTMZmGeBK805Zt5wxpPrHk+UzBxrRLHPCBsVoCp5LKCfmySUOyo4gMcpl4ngBx1ksMABYJt
fcFq9hDUvylbPqxpyQCtH4TCcFsT182drENn7HNC5d14vX4eO+KujKWAdlNroSX8JpTgZ0oZqFyI
5ObhX/4a29bsvnpoxyo1YOVmtBHqhtFmgs2wJzpYblsEYKM0D9/i/9HNZmyX6RCiYtqSdO4iiSiR
FS3oM2ZNB32uQHOVwavADU3hFzZvtRr1xaRszh7LQPfpLaylQOoMK1hUbP9r8ePYOMQvra+jf2VP
dTXvovrNb9JpvAQKBhINzGVC4lY6/7ppvsa3OqAFWYJb1Z+fBtRVFJVL/h/YnywR1FtK6w18qR6g
xh0iajzCuf7pBZkGZbrhRSqyukNiP8amOPs/HQXqJfHnPh9NZL26oRYfHpDWlN1LOuLZDeq47QFd
8GjKwBgXBO9fgH/UuHxyii+nFm9oQnwzZ+h2CoSECCe4ZXptoJkdRi3xuH0JZ24jLznDgQ4eFDvf
GhNkEbJmNftf+CRvD/BetirabXOOfOcEn0lVIUA0q4QPFiamjxGiQbslt2TDt/Z2YUXZqaa+E4Dk
uT4+OYTMmHaa2VcPAajyWsM0WPdsvps14BG+OrJV2Vt8WNfjHePDa2ED7X/HnRXpcH3t6wopdsOv
HJtyw3fzeKo5GekaIBGO+mMHuCmJGaU8lJ38IoUmDIs2XLeA3ZUrf2rSkPLcNNhtmBQnSiyWPl3F
s5UckOqKnfRq9G5RceEGHKhs4iQLJyUIgpwnKtcNEkYQ7YXDFdK7IugMBzsI9mkynZVIRZuexerp
QYtI/KFWZ84/xcsfcjHLxRKYK0Kuls0VSLcAy2w+KoQAVX7HbTAMtMCvDH1UG1+C632NqN3pD2Lo
zKhimxVYUGk6m+2LON+r706YhgX/qNJySCk5S54ZePgon6YDFZA3QPF/5ZBrQX221voEUSldfEQT
Lr8ayxe8SjdFbOGH23an8f2+f490aotjUIrKkw+i0pmRVglKjnNHPiP/280HJFFQJgE3b9NDvbn7
JUwqYXY5YXXXx1xC4CGDjhifcs+yllDaBKs/BaFFkH2AFJHxOUzI3kb5OlFPjgA3Cqd/RYF+In7k
oAQ1DV7rrXkpJVFloLhRLTGACVdnAZOiE6CGJTq5w67vJnV3drFHosjSbkJvwyGQeUYwBYtE0EQv
XRB8vB2nzeZrlqS7WGvnUIs4+bETRA7+5uUmlEd9UkSB2casXWqt59A0EqhdtIj08MFPaniCtQsI
z3iNdyJyssiWq2IE7jiEA2LO9Z8kgdQLmRuxf1CFP180NdUBtRRDEoSkha/+FSrXlzO1Kzwxqdyv
bJtI+4T3Y3780ml4RWOdXK4ASIJfk+vmqaDykcdtVNZbce4WSMFmv3fKEU/stJem+1b3RBwSE+jE
cM07tP37opnod+CS5AKTm0i5YX1McaKkk4JIKDg5qCYTrYsg2WRW04TSz8bihm/jJxWVRWbtsD7v
XhjZ/XG9riFI2DJF42pxCzXTMERgRDOmWsRB8mnfyv6sLV8JXGOqN1uQK1524rMDN1mWV7h3j9gO
wbi/DuF6bN+tPEWfkcB9FLXLEB6mzLfonXFggsNy2/bpRXpIkwX4I5s/eaNb5rVI1D1o5Z9sWh8z
6MytuX5AMLtcayNSeEzyKQLnSGntYnEjtqyjkdX2rhutetcr8j3/LAQsBZN/8ibEay+2AXQI+5p2
jxiYy1LajQ24YW6Wkb0dlFgZJ4O75dMY84s3CUK12JRmVnPnsqt7JOCuQT6axsS0Y6mEygMa8ybR
NrleE3hjztxlvXFN/jqE0YnX3813glqeb3o2YQUNFCiXWsbDzkIJN5bTt9bJgQJKfJxIbX494PXU
NzyvSWfQ/iQbQpoT0riGu5fitym5EZZcqN9wIhVJsq8MZt0zT+tjGCIouiL8auE6up+l5Qlu/1E/
/loxjlnB4nZdQJjnn+30660+NJLdhhOpOI/TosVKbSCwHyPD6w1AhMY5hKiM5MP1nWIvMakXaeET
6x4jnodmP+ULzitmA11MInLEtJjUK7l3KMjqXktXHCkudJNrSHi59PXIOKNXuIZymU/qPOv5IzPt
CBJVyr/z2vI9oqdR33XB1BEssvftmL4+5YDM4C0eD+ZlY/pOC2X79DPK6HW7DWKd2IkLJFoGgq7Z
/LhgKlorm740pVqDVsXdHs95opfYT3FelQ30fcx0RneDA1W65+VVFWM8xvCH850SHiNJX/5v4gMu
TQOS+ZHfUuF3AZsm3BB75Fzl6X+PTW0jeZ1vaDLUaVrpWkEctEoWkylKiIGtlK2Y2dY2s6g8h+Po
WtjViawt6Sd+lebXdWrVpLKvwXoRLv2GvdtKLhGQwfFTULiWBchhMRiuBQdJrqHI0/VCH7BJ5JRd
YvYe4r+kGa5Xx7/NBAklTWmGSJQLIDtLjUZNuFKLpKujkEt4wYiyoGLonsxXq0wu9HFvxc5kuH9k
gZZAGyWKJ+qox/kxcQ27UVeRyYtAcfLM0aPvsKeUIRJrUIBquYci7c0DPRUMwfXBr4Qp6wHwF4pZ
oHaXjn4k3XfDuXmXkJLgZqj2+IF89Jf1KkUYjsg4jFtZLjA74jDL/2wP2okAkiC+0TVrSKJiVVCF
mYRDzdBeim3fJ2xDx/MC5/5G7uICHk1zEWnHj0DPA2boe0lmFaTVLwGr34/m5xJa0KBhZ6MV+MqI
dDwmi8oFENj8LUdbWuq9dgXvClzBYxB5RI0ThlYH/x2AqvfrkMfCuixVekhCEO8wOmzvBxb6zphW
kreNYLqBZ06zhj2oFy6jojIhV4iTG1hYxUrufcfhytW5hYGSOIhqD8/VmEL1QPVt4l7wifvcVlGi
giun94iOVdvfMRUlRgVeqVd+jObcYe0Pm3B4kb0dnfegPgGX4S62oU3QUl65dVjI5y+UtsV5z4EA
d7rHo+ceqjzgXUrF5hQpbH4nGR3fZFeiaCgFBHAKIDUN9c7VFK8WyMjiC4Aog09BHy5Fyj10javR
kf/8g+rERuoFDDvpyHHAxqBVsK0OCD7c6/pizYbxkDirjcqFknrYnZdkpQORG7HZ8vsQT079Sb6b
Nt2371H94bCdlO2yEy2BgUCuFfllB9PtNi1kwa0J6qpsuVW4de2fZ5kQCMpNqURD1UChO8mpnIrD
uZU91QBHzKTToW9j1l/e/I09OzYy7Iq9LvxUGa1lf2H1tlCX6bo1QzxFU8bRUTmwBdWe3WmETPck
shu116ndhSrk4PdoDP3ZJkChk04jaqDfJ10ac3bKvYjxaYx+zmUCzA4ZP8C7BGe52AA64jea4wtW
H4G51hs8s/4560rILWQJ0Qh4xRvyEjBYh3R0lqlH/irVcQuj6yy4HMLSTPcWWsjm3TqPsAao6FeF
QB3odMU8Jg725X83TlE79NU+Phu8/w4k73wkLKoVKWqplCHJ+6/znL9LpY/Le71fguW4j5ot8qNd
z7tOf7dFa6n0xIIF472DPkPvf1feDdtlaiYXi2lNgFWwJNTqw9X2BFrTuecoak9BwRRUXcNnQbqF
4P5f/8hr5evL4GVoYMGnrUTufJl19kelRQS4sa1vKRS5Oqxpv5FJIHiJ8XSgQalPSwZPyz77JpJu
EgPl5BkNJ6pdG80cI3DYkyzH2iEg0H7GV//TCh3ZGwe+qbkEuaAoIFyF52YwAlGef7ssA/pc+XiI
QbIA3XBrI1tWa9bUPksd86UDUi/mC7wCsQwx2c2V6JIHs9r+2yJzDJx4HcNU9gj+2zeu/T8cov22
KwAZc9JxExhC80kauSA9utkvKAOBldz5BZv16RthagPDxzgygG7KNBUdU3trp7zD6xidmxOd51tE
3+2mF9/88I+G9doAOHKmjAdhueZPPtzKT1Wqb430w0uP8FcTF6lgesBZzbfb8gT36Jmmvx3Ze+TK
pJ3+QxrgGwIlG4HmzO/qIaNkgDUWxWMf4+pLRe7PZS162BXV6jyKW4zDQ04PePwBtwyqQLrVDxy7
u7MrSwfX4cXitL3D1ZJkxOuK1mpzzxy7ygLggAC9BLvgZF9UWjaPC7qKHs/ki9nO9hTaN0ZeAbT3
zXoATh+6ouj3AyxK0Hdofohtt+rxaZsk//t+pnsQUA5uVoHJguVlsOShE9rCVR9+g9hJ00b7BSic
rKTkbQ5YTyil9SmHWRPMZfPR9MjX1qsg2kxTb+7pjaoW1Pj5I4zYwOmycefI4J3eCQwvhcVELCEh
js+JbHzqTXWMqFH6SCNg9FCW8tHWxc96XfFabrWrYfzZ/jWLguGbN61Ppi4HaquM/whgpHujid6g
TEL//ERcqyQtgdWgMaxTGKhLBLelXLgM6hhT8qFQXgQbUrcL/eH/lGqV4m7Jnc0oSX5t4IAS96WH
NgcoD8PugKmFZPQOblnl3ZyVSfRRa1rKpnI7oL9dE/+Z5Jw16oSWJDyruEraytaCuFXv97/TLtr9
tjJlxaMvaVnKX8vLOJdXfxYm+hdVI+B2ibTqKwi8Dmibgk9hTCTzp7owROg4eEbC7e4DkCS8GqIO
cnNE6UEvw26kOPj76F4mIZQHz1F07YRMZHLx8y53OOAMwwvFRwKlTisShI+2ZvSD1nRUYOZulOie
faH+fDjDprjcrW/lqeH36ImXoczFC8QquH7TeBq36DaH/Ok6V0tZWpcMfpPgl07ok+iJJzsu/pDp
UJVJBQut6PmN4VSvHOMWvHNtjAZ4kRJ+SwLXoO90No7nGxXMxoCDn3V7+hHhdnM9wZ6ueM6u0VDw
B1ZXDji2ZWQyrJfipTdLdCZyQchmJCSoMEey6fj2OUOA6nPb8GeT0JWzt3g5qETN6YabuIt0hB+o
nnptkMGNQZ6yg+yYAFmKV/CcGfIK62pHKvtHU8J+NhhZlrWOjX/NKJnpbk+dDoYemt7MeMVGA2OD
xuBPtsLYz3rkU/WnWMEXi6djqEBj85aBL68sUNYtDM2rUPkHaMtMyEQl/0ErV4D93SAQa+CwGrtl
CYD8qe3MK29wUj/ruZsZiZiJ3WPBthW4O7oiU6VDVyXb8DZQ+zDTb2at3qHDGvqcCV1FREjQ+wxJ
J3vPIQxEz9/yxSPyz5eA56YsramY6CHvUZ3tV0jhKd5n0Nh1VCWs1BkEosndL2oLkqeYXeCUpBZQ
psHb2Eag2Rq9d5I9weg68dfiki5cC0W7jdu0hAP2dHeUozf8n5Pstg0N1zglDveeK5CUfDfbZ8Eh
5ALSKUgqrUBjY/5M1fswdZ4ORNK5YPIlp98lI+iMsU3sfHkxEYythfPjmeSLQHsyoQiiSGc8qr8J
DuILyXlAjbeg7lwea60ukqc8YCJj0mEaEKsVI9dK8lvrkw4D+AoepLxUJqhnOL6xzSv/9YCjTsSB
/PH1KZV5TYu7cvcK5na9d+M2v3MYZlP/BLIPMh4VmkX8M9joQ1QlWjfPezdzmQl+GoyOLIy4VWPe
1/MaSDPVy7Vz/RFpbefuMqPFbvR6yQ8fgwddx6bC8tUv0m+BP9yKs3hqNEkfeGUOmqbWYNoMNXbM
n0nE5guvGAVwbLGTjQOCEyNkU5P2y6DcXm7XRU3s/KLqYsC+D0RUiFTjQYhLuyRkgc8gyCPkB4iR
gxY9AbpPTVJ9vbFnVMBlrfaxXXqrwM5N6GppapDbCG12vl+SdNzhMd1Ki2eI5WljgVAQSZs9lrlB
58Wa0H6bRs7e1WF8EooxoJzBd+jTwMmVxJw1v/x+fCaaECiGnVwkNYs1w4Uj6gKn1HHLPuai818r
PVTG4xaUYyCaL1o4N0HlglvkubJ60EAfaqm05Y3aVZn8F6EepBv6ASxYALZVtFnXDlblvCFf/q8r
9qDJsEEQNQ05JQ/qV/pqn6LXf/h0cIY8Cr/0a6/TDf1tfUoc9uzNEFz2C4RpnyjYtuDc1c/5p4Gw
/qxhAy21cDihHSOcPtMuLgMv0UFhsxT2qVxQkXlhPYvkXf2vB3M4oOa0DJ2IEZDmO6eJYL/YvjKG
pB8hUs0dTD6DXEmO3ZVtRDXTSclwiKZWnf9isMoEHL5g9p6heFNM+2eLCiAogTGhV5Aba5jbKZCx
+TIv7bxOFqj5+/Cju4zj40Dk3vH5OU4Dx4QnJPccj3cdZtkx5ziM0DbbeqeUwvM2hcZW1la1feBN
wkd6YFghTfdYNmxlYG6DzkGikBdJQjGb+Gf+Ha3vsWJwvWP91IV4Kd2iCFHCFo86MeyHgex1wLJT
X9JSTKjuf/rBQRWrd1ckGuZxEFwKbqTQ58P+3p7WZAf4ozhN4J6PwJl9RHNNwJMar3ImzjDCvFL3
teNWCWP7uQlF9bMCyLEIzq6o0co6lbjrpvFOYFcTm350r5rzA/4YxtYPSJv3XTzCmyDAMKhur6rE
eBIKSnBV4c5LOtvvkxAWHG4T2pqz4ssvAKm5lRhBBXWpzaUlR4Lq+U49LEDJ4vkO7odpf+47lYoP
Pk5YS47ubFKchedZ7ONZeQDEa7FxTsrNa6pGsEn166oYljm8rE1FkfSuXOIiRw66TutDDGVwlEmF
nflTOp28VuGG+bYjdt5rh3ic+WkGEf8X5rEr+YmHScXKRR1PcAo3QJ2ifaJPSwbjge9JOCV011Pl
zv9USRhTtKrXK/sOnjEN516E36AUILDzb25WH/qcs1r3/KhdwyyDtPfwc9RZ3IQXNV56QtainIlL
FrXZoKwgyjHpZXiKgZWomzJLlwE8ErXc8keI48sGVdcQmv0iEYaLvOSdO8kZfAYqjKBpRSjfptru
aMFcoL654dQxzQDVWZXcgLls6HSryKaTD7CRTYC4uX+6gzYn1qcasOaiA//aPCUvyyYrF2InypPy
Skfuz3lUsx+3nCU8ZaIcYmIbqRME/xDAb2gUQq6I/22BeDtcj/8eOolnun5LGAAnBGlfYixOvHc5
v+s/ot76mIwot6zyGRQtq4UGYemxX8XEUIN8G8pF7Ufvj7XtTajnM7sTaM1JV4/WYEKcglYr34am
rcipjZ3L+UcJVeeMqbmNcvsKQVNOf/NDc05dAYiqKBR21UOkHKQypvrjetoOVMi44IAWy4lpZNNq
lMsAbbb1jwYL7oeHcnPDao5G+kY3/KFyAY6Gd8PkD2p8wavteTarBqvLFVNl/V7juJR5kqfxqm/W
ckEp7VWXYUYeCx/C4UNjXfDrn/v+hCU8cSJw8yXa+x3WXNXdH/5KXj3ja2tEgZZe2Vw0jLgfHzFQ
mkrEkhjVbeihXNX7lFUp4DnhgCXUEUKTq/Jk+whhqQEQ6N4Jk6UMShDKVhiMWBhfzvv7X3W/y/pE
P7k0hJC4ApY5QHb8cWxZVOxnQObU2aPngHl4g0PbOF0oGYHp2ngSH2MzLlGvPrRPASC0V15d9E2e
33z0Glc4JjMkuOCPQie7dSTkDv7U8Nlyl+qKJ311Hgk9+mztEBsCteErA33kW8Z9zgbKO9LHsd3x
Pvp682G77PTeYEr9D3v1uFuTyEv3LsQ2iO8FHLfHxQcg3CuWGL3H3p7hlrd+P21kVmgJE1ehElPC
RUpF89rjx4j4Qw2MJTOHbKYTTXxO9EAMBLD+hXx46+QHdj19tUeb5oA87ThuXWwaISvZbzxvT72w
qKpNM55VVPDCtjNhpzluuT6FR+/7Qa6DP9/2y6CcHYLh4VosdWlKG1Y3kFqYEvHqOSxfmCIW7VRN
9VwgmrRzdlrzXBWA6c9tfLLNjJcD31KQtlUovktb/SPBBkWJlkZnnSFM+Ywm2nqSvpk4WjTMGaxg
cSHp+pRUhTxxvBpsONwQ9C7aPhAqD6t1jVDK15jqpnAeXQW7ewAmIlkWG8HGw+NJllrUHuYZAU8p
5lWe/JJactELdfOX2NROrrwxUsLbDFfmL6cwkevIsiNiUtTE1BwuTFoM/7ogGww0DdwwbmCRvqUq
+kz9+rYKoKLl/9Hz+vtxwpEVtryBjcs24vv92MBbE+A3YpjQ8U0JepVbZb1vHSgRONr8yeh61ti+
+9S4Xwb+jVrDDxPTrRjaubZVZ8KAmy3Er7+V/fFDrvGqmywzpUaUAQrDcjqPHwDVxPQUlHHcDOUH
naoL8FxyHh9m+b5oOrINwy08MmG+lr889SKhoetA8EDO9GSosM3pOh4wAx1UuO4iiJiLzheumcKB
c9MU51irWd9yoFvMnMW+f1U7DRJakdVERQyeChxyWO4xhb+psAj6ciZwbzEiNE6zoVwiilsFKM7I
LZYy0uVIAmfu5ylgioXt7Y555WIM8Cz9JK67EtkLNCZLitKnQQvFUCCxUOAt3NjfcJplzSxaakGi
xBqWqGMuVr0mMxootkHhZp7ldKxT8o38Jcrw8IYV8gbL0D9nVkJg7e1YoYbK57ZN7HYmtUmIhISf
q4fcXNVUxX7iTkfSGNsZd1scs1pw08MnG34eNYdi7K9ViiOu7k+hJ4uATrmdViQROP7fqo91LmJs
SXtubLj6hhbItT1lJyK1Xzv5+WoDpNax/Lwdiqg8PDRoMImYEXR/2r/8ibT26utlGylURWDcEa1H
3nT1ZCLgKUi3geBRMn7jXH7IjcZQHYffmgsutVOinrXoSSdT8HXs4rI6L+ovOdyrx64afHWw+zC2
zpYcY7TKwPdvwgF9co62tLwKT51APAGYeSywxzwmlt7FaZosGUFLXuUm5+uxhXuN2u38JntzQgMA
zxlQoJUDbGObPRhwTJkLp2iH4T3bW8R9Npd2Adzvx5hVhL0DfT3PNvi3krXQ36JxSUhCGsu7atnk
cd4rZD7crgVV9Q3nKF3bT6iK+H8usOyH7zEyq8oHQGDvSrP6tSOdAn3/LdMXRr4W0HlAzYSpyI5W
tJ0l8Rp2CXaO8R5FKCq2TEsqPwt3CZY7j6QdHCSHjWjf4SMebtG3Q8SjSB+/fLIOZoQY4TFHIWyr
ODSmgKizpwiNJY6WRwyxYWGrmziz9xpMG2Xdy3nebVssmhhCykyzLpIMw1ePxnQRKHpZk7fDM/9M
mIXP7/U3SgWpELQsEQQu/ssRXxQRCFuXCcGDpR/wlHYYYcCkkM3qdbzrlQMROHY368wtpwJjf5TU
ywgZ1pMZcg8KlA9abpeNgquK/qxqeznH6Rkc8r9V07bPWlcXCX7CIuMhWNNeNJ2DESPajfTNYTUC
jDFsazWJ7AMN+TPKN8cPO3lqeyR4KrsbjIMGVJmXdA46uiSFC+uxYJFptsS42QIbibUHDm8nkLzZ
CKg7i7AMwygtz1AY6/ATPtu/gdFt0NeGSCozGU/Yc5/XhqMrSsueZb7GHK9EQJQgBmAeXCdFI2hT
Tsy87L8yNkXpo3thnkfK9nhZyMUUv9ShjmzdFmwA3ozWnwKE25AHAIgNky5kFwPZPNKi00hoWJ0e
iRvEsDflINZ3MpJhRUQtClhpx/uqBd9OZhEEQRVxAQqDSxiIpItjaIZh//euQsLsGOg/6/4VWy4V
tVSIy1BfgRWKs2054xH/H1OkkrNGj1iobls4q//W9Cc4VuviQJECOaiuQuUi9SL8J7e4OGSHEofZ
/L3t/mNE7dWQtyGQ8t6CIaClo8YcOynapBpbJLseQ/ZjC3YjXlWa1SB0sEAl9Z61l2dAZEihg2nL
LogtJOpRhsUS1bYtD7UtKJECQFV6279y87I+Gmfq0Xvs4szyIB4Z8uiWgUfYEhI5zRZHSmX2ySnY
nYMGrer8hR3L0WljVQXLGaP7zB8HYN4nMN/b0lsM8/U9gHdSdtTa9bC79qg/cAiwjlvW2ldY5UdM
aMRUBnVuQmBpwc9RSWNV8aPrmkA0mQZVcco/C8K8M+MwouOUvWg6LCSLrKMmb5j6JOK4KldBipll
TlDdQ5t5KfbZ97F5Sqp8gke81O/8h9FdQOHg+VGyZItp4R2jf6AN4e/BndbV+U/s7GflbpUSujfr
ykVJSPw6R6raDfZJuJ+Bk5AXTVVlNmCPXxOCLuvkAQm4cC+ODfnvi0nqY2Glac7NZRvScjMq1vmD
AbUgSu6Hss8BOZNNdMl3uWo0B+C0SQH+UCnAb5t9qXUoHur2oFkDxIrFktzLdJPlxqzZRryyPmK1
X/QUki3wBDxyH7c7mrY9jssTkf0v8abv2C9NLtGOb2IITVeYs7WDRcDdxMSgx9XwJzVR7KuPnHOO
1e7jtPhs5eELWtbmE40vuvXgjLwxEJnvmS1qJnqvmYbqIGH8jLhRuJSE2YY97HG6v7G1a2Wz/yDD
eLAxcN/arghQAnrrnR40JLKiO0qDqlSM4Tw/8XpMWe7cjDSnNkogv2lOmHuM72LKNhWyT/CTX8+e
0yrLfOCouA+RUIANnKoqA5jFXj5mdxaA+AliXp4JnIzdyiS5vUG4SJUrt/hwMhy9HEAKiRpK0goB
05Lvxy+ZOkbgjTwIdkahGa5UJjgLb65gDIB0NW44+m3mILRrkwQx1gzQFM7VbmgepMe6g5rgMwz3
JKuAa/fPHXXUB3sX2v7Kvpbk9fi8DEI/e2Ci59yxFR0bTCohbGBVRsF+D4JhgmKFFVpLkd64M1MG
qqu3APWtOmHW22jJxVcVJvTOcqKM6kpZf1pWZHNqOrdk8ZFoCBa3oYyUhmeVwB2kHT3kPvAkZuZF
svy7zNpuGUg/oh1gFF+g/bL85u9fanOD5m2B0boMEKUFNyz9Eqv/eCxKcZCt3fWiVLfHsTQPsb0f
Zlk47ZtNbxoKVh1g1GVjNiIgDg1XJYTSBepayPY0UwUVvM8sRgOz79gyoNo73yBCfxx2286hVObE
n7gIxX5vENdgrEuLnq9DzHGgco+zNq9onVegtrvnDWNeYTIgMMox3KcwA7QL20QfCthHn5TIFHak
PH9HYOAzQRcH64DUGqLde4SoFG7iiWMgiNzWQKEOoD8+64ZKTa4aKNE2IA0yjty1za0IfnPUvmvO
3LpRcucV6bMos7+mPWSVFp7SGLSL7ugpLY2pb2uW9GvBjYpGEYRtbORfYdAt7WRX2xZhthlhQa0E
Hod4lTGXNNHHxe34GVOQipbKkzH1os9EQ5qQqeR7OtAF0QDTbgjyf1jEYxqnWruZKFL0Ns6AHAzH
eEGM+HhQdEygD4bWsH/v4RkmhS/EN7OQwAI5y+BMu0CtPh5AHlGjUKHW8XNk80+cPWpVVFNQWKB3
6ftdThVbTXbVo+86yzf1bK6rTT0HyMfwm/Xxeb93zsAbtPbzCrtJJTB/lorzMWguyiaVFJc/ZyZJ
O3rEWMXjGbYfPAF7Cqnxd5eoS3Dpmyl1r6sgc7B7BsbPTxKuY0d0lcGuUf22LEsUetc9wxeT4Quo
eUz9ip6OZrvQ++ofis20VfmZPpnrh6ELmC3qyvoA7d13z+/9FmJWUgx1TyE52mR68Okx0a4LFwOr
97SGzSMD3M8nzp+l3IT0X/OuSb94M2S7haQJ4Zc+6MyvOeJ7/eaHsk42SFnIHXxw0+S/FsYEN7L0
1mQTLO8QClZ86Mm0/tMkjDLCfrFu29P/0mR6GNlblzwKsg+u+3Sy7q+Ck8ku8G3CSAHGEc9oLTon
CftbMn8LVRU69uswS9cgy8hvZ1q1n34d0PtpGtfi+ag+T4CAECY2q0I8bQAyNB1jL5ICFzWSo378
38u+Eu2A6r6axBl6ByN4oIq+YXuLrOfXIAa6Zb1Tc9fj0115yLkLKaAYOFQSBaGvcQ0OiWlUPpph
Xkt3sylMfl9ZhT8/F98vc/ySgvqumzQbEcMPA/g9x2dscWvY5QSKhAaEFrxdv3M8HtN2HhMW/lu1
cIXqhAfwVokJCIYq89AW3h2wwD4+4/ow6frhJe0y4Mw7pprAW2O43C+F9ZQkVzKDh0aeINdtNo/p
rbK8rz2mVqi8HZt2s6JfKrBE0/UWq9Qv7C6XA7WmZzo4wXZlYE5lFvf6rlwvIKFdQRRUbHWNudwQ
pAvjxrYYaxWkPBovoDvOnuBeAqW+W8wLXDaVtnJt5KUwgdIRllUGK3N8znrSsQ4S0M1PqMeYL85j
drsAlmPBqnGLKMRb3vnSGii5qq+pAZ8abB5M1jgbtf+nhodrlmHhtiWonTuQel3u1CNeMlGGL7al
MUfGf83LSYlWmB+jvBaSUhr8bcy9GvPImbWLXp6ihknnnZW2C+wgIm8c8WxrpYSxi8R5j952xggE
2QFRAjyR3GTPIXDGnVekF796TuHWoS2PLFy3GRYgXISTCWhX5aPhtykHMabCYOyRxyQUpJadiHmW
v3t430Ok/himKxm71Qt2AgTrKdLyFCbAbX+2JZDZvdfVDtRgwxxnIJ4yL3zmmlbk9aih/lOe0/VI
Bck9idCDgmD94MMFJEOKhuqj1MHKoiNMoO1MA7b4C4We+52LZBbeEQ+3oJ0k5NbKbZCMafSbZkmq
pDq9o2Yi0ZPeNwIZkr9ZkUZmHxQ1K3Na6wYrToxnCVLMZ6fLnt8K2YDWNbXWF27XI2+q8cfqprbT
mhXQcp/fXoWrv8ULSvyYAM/bFxo6eZqclC7RmI1pIExbjbhKEjo4ilZ6iewtBQ6aA7MZegRUZKCo
AFSRUSxF/9rItgoqdfpDbfLoQs9fjaWiYUTrUEiAKwvhIFl/q60I8++j3pjoMVWP1y9GhvKu0SM3
wFvwKpxkU0qL6C1z1WYxy6Ln+8G4lokfWLhQ4Ao8El35rCYDqWIM/Jyp6UimO1wYmFT9H+5a22vi
mouk2uqp7DM7ozUjtpDwEPXSoUcHWKZj7par57uqaldw15tFvEJ+6mkJzUHWW6XsPfyCuHAEmaWw
ehlgpgXh/0cMwOS5o2/BAkx8BgTmXeVmG4GCjTeLxqBfOm/TWoHaO/BwifXCzMMJaqLdsWeDyaVE
0v2H+zTrOtzcJU5ULWSaMq+M22BmDptSGkq1qfzX9LaFav9ApVIjwvANQv3w0gtTpe2tSg31UDAU
5H0F9zG6DurL+1Gco3ThlT2NTiljJ6QprRuNImV3OtTY+anViTIkeuIXnr2UbBHGrfSKFq4fimVA
aeEjkftu5sidumdZ1RqdK6YRNLdW7CfBHNMkWWQk9XhUS4sdtnm662QTt7+qcLJKm4Csw7kddJ/p
tkz+EcJ3lek1w2DFsY04jL+PHoF05+UEgN+840VyLQ93lrL5R0uG2reYVSV7V/3dLwq/JZSAYbtS
XL8WYXkJv80vavbl2PouVuP9DBzpZU2GEoZ+zjEbsXZyfToQ2Ep6+eqA/D0pnwJvHt4l+E5/VG6H
w4DrvibREpikjM+HDXYe/raFdCSiy4ovcyCH0ZbeNKATmuftH4ySIoXlCdk355czzoitbfezT9Gk
hMBAWdbn4TGC42q1iCyqtbd3X9bKRy2v4mA2v0K/Q8xV0zKfOBrfP6Wfpb9r3sOFZMGt5kK74+Bq
5GzKKqsZSnHCkWVoIpeV4y54m800iCQbUHD3bCnkLOk0WPljTHBsBTHTN2epIZ5PHEw/I17dMDMF
jcsxnpZ84XemoW1zIT0cVgJ6Exbom8zZ/gfIrlcBRv+gafnMQhPRF9ZRLEnFuzfej2YsUZO/dlSD
mNM1lBw86jnyvjc0pDN6CxSGn1cCMf1OogQwjdAqAcdUI6oT78wdsiG78daSSueEtPVml0O2gwnV
d5RhyW7UrU5ulw8THTwlbIQWZiQ8iasBbzKL9B2u+as6jcIe560i1n+FMOTDGDpXsq4YyHIdl3xs
0sHUaFg3iEmok4vjD2hkIl+Fv1DeqxR3RoWkRCy15BnAVPFjnPYdq+xI0ib8Ycb7ymdPK0FtTSD+
gReWdPgN3DqkAqtMrISSCnqCG67l2YIOvH5Ojiim6fzv+6Du08UwUNsGviGCQ6RiSQJb8Q/5HXL3
xyJ0EbF51lSXj5b70ReRi0xSrD7AtOA5e9oGYdAT5frKukBEhlrN0evQvAoFq1IIcDXuZw37T4Kx
i1D+X2G1QZbsb/hK3vWOkBsSTpsYk9op/w2EpYLQZrNgST5B2r7OPXgVG89PT4reD88itpYSYpt+
ke5fMyoQaTAJuYBXye9o0jPwqj9ickL9lAl8+jpruwIj9WnJ3fm7vvAbTI2HoS++u6qfsqWG6EL6
w77R4OhplMfz9ZQQ0iPra5gdcaJyZNxLcWf0NSziYxs5ozLT9fw0WZErckZuvVX1Uq7H8BipAG7w
L57AyHzKVzKP34p7r3VnIAhun3pAaFdt1HBC1GXXIe8fYsOuZbWKhdfnrp1KunGHBaof1a08AnX0
OFyS0sYx3dxbBeYCY430edUr7Lee7i8M/fRi4EQGkAi1lI+UOEUXQh/kYSUidD83uBwBU4cuFc6h
QO7Lq8obYvgiPFJj5W0Ei2Rx61RRLwQNxY97Oe9vi61kj0wltWy8eYtO5STz0SlDaP4T2q7EfM2e
KuDyT0Uqs3mmTZFkr9X9wLVDHNTKYGtpz//c0sbTPCblABs9HApik5JQQMxM9yygD78oPO8q1aBU
yxPfu2snr+cJmqvOsGAd7MHNwznpoNRh87K7v3agP4YfND0mY0zBy/Jjm8LGm9UGTOtYersVZ68Q
wh9eiWHcp87zG/FPujOCl9mK3O0o62hjFq2QfFacE7kZ+axQULkwGcsxyasovkZXrW+2eGOvo2TU
RZTAjAbei0cCOlfaXN+JpoQyQnxBSk/mp1fAJE0ueb+9XffapTFeguP8KiAWXcZ8pWCQNXdyRZ99
hTEWA3g5Z358cBPzinDIkFVtMnZR95yV9bxJyfiO0+ClukcgD3cTO/osSRu4y1EbcqIrhiCV9hWd
70JNub+EJOst6zdvOdOZha2adQ3lVoynJgYV2LksVjxVw//MYmwiWV38P0eB/xdlBUqYmAFV5pqB
6jHpgdE5Ac2S/vgjkHs8jZcGw3/OQJGgUZBczI3MkKS5U1VzbtnLjlPUaScjQw3RzoskLX8Gg64r
D9JOvjK1seEIyF1iv85p/XHR/rePjGdJoEcHjR57VrLur0XFsbSF+EFGDTdc57uwxkRhOEnfoBJn
noFeHbXucjWXKENiKHFdsYDqd4TVKmiyREmOf6EMI/eU6vihge6CwulmSdYzmBGpdERImwUrCuri
E9p28RFz8cq6CGHu3B1qg/pqOSsTQTO2giXdMmgaf34suF8lsdTwH88YoGIf67NopyxRa4YzAW7n
0dk+gB+dLPAXflUiMycuwdj1Qw3FFf7gTHh2KLu3ABnpg/KeYvGRCyzNoFcQTRlKci/dnYNKv9PI
NsvylbsU7syiPz9x956goW6hrKqdQ0gf2hPUtMik9ont0NcCJYkSJ7EhaPM0AhuS86WC9bRyycXA
VudwVHnHDdrRFp7dWM/vt2i0yQmMzMnIDE9kjDheXVknvAnrdHu5w0nlaB1Rp447VMspCsPB/uv3
xWqO9CexuPfcWlUeckod5v8OjMNU+z3jYObXbClAmoOtFNgxgK4GjMtITs4rQhZr+4YhNxGXX8u2
yBp8qwGwYMCCVRTRRHlnkquuKbBqx6yfT8KLYbljyXpDoNv64u4KaMsF8N11uj1jzj/utAvCsljL
LJgSRNwO80qE0UExfeNj2GYuV/6YIBUhC4Zx33dkDF0zmfmNE3RdM4m5fnuJWu6rxPz7G41WRYjp
S9S396S4k38lO5LbDYq2NQE49S0fHgWhYZm13pjnpPf62lS1Nn5GooJ4TqMn9W5mB/obtM77cqM0
LJjp57zXbqAIaPSQ2XtUFHBK9kWU+OnUieZC0twjERpHWPhXMmBH1UHqQvSVgPN4RGxio1yB0kpv
OYGkGVOs88VQAjiJFLOqOHxmyoRr3Imkqna2ErP76mMvbuvSMBvEj3/7u12uLOV+4FOCnNObOCef
ngw187DndniZUt3iL70NA0Ae/bA/GjoDKMPcnc6y+78cHUbysmUgleGW1BgLOA5Cm28zyWw7l5Aq
N6P7Qd0AfzyOQfdAL+WtUU2fUHSDGHVqBgrxUyWjWkiWtYPUSDc747f8taPhZbB54O6lqxH0Z4ii
DjdW2FPJMcI0wgTNL0v9ljgyYySwROHdZDEq9B1KSdtrQ3Gp/k+TsDL/gwsyTuQaBHu1fIXTozMz
EH2FZfvEO+GT6Azvs2/iBlZbsAy2jKeE3WohdD6kRhoiv98/6rFZCQCar55c5jiywMaM7o3g+nPm
1fep273hvNqsSLTKqAkSZs/kaj6bWGvZBlvamXe4Kppg8wsEN66kDr5OqbPQmi7PvQVWJB0c8pMz
3vBb3kanFXLdVYaQLCo5mAEv1/dJl5CtNLoA5i1AN9Jkw92KudmvrJQQuZ67EE7A2UXOD8wYveG3
nP4bm9wfOi6C8mbOnIGfdTqbgq8SeL2UgZDHH6n38TXjoCVSmR+Yf8qcmQ1tKjTDOKWgiTK31pvl
QEwO0oHyTCARivUqytEO8vfu5zoCdVOTHKV3U6hEgN+FgZWvS8tI81+wJsjfKj+3QFs7MQEOEtUp
Vk14gWEuO4cAg9N5DrNWJZOoDtPKo+9whtss8qtzOC2FM88n5cbdZ2ja+DmUmepOWzwyZajzDyvu
v55I1Evx6bMQVM9PwCiJMXBgDqN9vJEX0G7dLwb7bPTo3Fhqoc46u6iBAEx0PhZKpkbxe9xWKccG
19UlGI/q2P7O9gDQVArVyIdlT4qVuxkvFKuwxD01f0aylEut5uMQOupWoPd8BeEBbzS7cO5949OJ
j6zN+qXhAUSnUVdBMIxKpPSxbqBTADFSI1EisoqiU/UL55VQ4ETT4FhcudreWQIvKOZQL2N30WrH
8blMjrRGGgSOd4q50lPpbdkf1RHgdqg5iHpCQYcHhew3iK6bMgfnyP0f8yiXBtchFs3aYvEUhhcb
+d937ai+tFM2GiLBrejtheM3zyR8NdA9G9tkpSCqIk6ZkrgQviYA2ld15eYgJjS/2HHcU57OztfU
mAcOT/cMALUp6vwYxs3/R3FGKViOmVZxUHAZ/OHxtZdFdXowNI8jrJDIPcdVX+SF5/cfH5aPB6Jt
UBgtt4qEjZ/CoKdkhcpsVKS5nuGWbFW4/qA0l6Z97iOhc4u7+z+bnks/XzQ+JBBZ0m0t/NkyOOhX
T9r3LZUoFkJ/3TsOY6fPf2R0O/XdKdACc2+TlbakRCmJScwMCAIBXoHxgIzGUmb+pnz3eAkb4fuM
6Ibq6iV+IsWQwUHvurnNpx0L2sb0BDwhqsQdtzg6sz7/vMCmgaWgVKWvFZPMtEwDsbfbKZ23hIKz
kXNpz5mgijCiFaQqjdPLGX40z7LJHhT/VuL5qQ5R+tZl/0nsNb5egA8P1uxJkM06yjSEYCGkO4K3
6NUC338KtOXzGRs2NtBITrtR39NJgDUNlblDlmdpB6BXhJf36gJ5RLseH89CxnNpm3Sl0JBN4xVl
Xn8V5R0U1HOrS+9o66sbEWYBzPsVi6VyoY6UrNP10eUvEcgxdTzwqBfwQEpcQmAo4Mb8KJPoOdFA
rKIl4XtSY/dZa0wn6FHYku5EaXHQvrKj1dLXIlDRW1bKBz6eeakH5woqAdxFP4Q/FnXrbw7j7hIc
DfFKErHLUewoX2Xn452B/+GI2kMoVMwcTMETvq0sB2SqbZrwdZmRsNnWw5MbBgnMA8hfmoyX7bRu
LS684X4Jgd6eMGsFaicsCTemnVPstMEx86HBTYWcI7uqtmsU8VA7gEsq8qiyoiNlNWtVoa3/uj3C
LxhtOJv4KfXJFKmuMJcgtbtn9Yg7kJzI3G0NcQR6PEK+SvtHvj+gLTkBg1PD+UoyqmGvCbI9eH7M
TZ+tPAmwNDt5+bImaHf7FrwA0j1hba+FD0MOSm2qtgvkqAtSm/RmuU2tf/n7yPZm3CFRjwSvRKar
FA70Hmv3BWyg0V2XxsiCCcZJJyiG7kHazAWCQ2E8DN+8PlzA6Jz96aWFswgEqochKM78OxhypXG7
GQXIZySMIU0DsT0i5dHJ0MCjhCV7yIs4oehL7qOa5qmj4JpFxxpBLTMuY2JnNTRSJA8MD/ASxe3k
h3s1Mxi1McPsx4Hq0iiuJroT7/4bJopejQpsCcYvLWmAjNaWxbdCq33DUmFPkwB0427BIVQsQNZy
/CfuQa0r0wy4h3DcTneDEvu32xl92LyOX2NJXs1rZrp6WbFOMlSeoCzPmFFqLEc7h/a6aA0KNRGh
5q7bfyQzZinGmISn36AHnN0Y4RS+Tp9XF0xFxHxe0Pd625M+vQXlFQg1L3WO76nYjOEoRO9AEf0K
8vU9NFGuqQDEB9pNwAtvE9pF1x3/io0nTkTPbQehW5IoOL0hVhTvrNeu/ZArsUHSyES0O++rk/HU
A1xDsVppuFNu01vKQvUclnw/uNJP45tt8hJInhHnQYt/Ok9/juM0LN/ly+3SXrIVjEQEhEfuKLww
a2uMHHaJ/ofS9U/tAZ7ASVcwh0mHUVF1yeNiLK3RIHNW8x1yvzygK2eOBb5Bsd8Udz3ThIQAXkDh
2uAjVgfxLRv1asSsDBC7ZUQsBppP4ZTIczffooPOXTqkm/7aQh0JIYVOH2jP/3p1R/GeGpalIU9X
G/PsgL0jsuMibfZJFVAhCeV2CcBtmX44fUet+L4rr92SF796e3IWS+js24kpJzukCFlNzezJ5fPv
L3pOiSOr5lj5BcY6I0RD2TrfzE0vQgFABAoE1T+XKpBcfQwbX57hJsFm/Ly/k48hY/UiNUzfLfZx
1Z2L5ObnagW2KoaSUz4rZZ6p65VhPCjEzkGhsCM7OTi4VILd/ol2e1wPaANVl0Q6mD08xfWhe6ZU
hmhuIGo9VJ9vnJWj8S4LOXyIUyvdZtratQRStzEgILweqi6zOjKqo28Vq2PK/ZnkXRgRjYEd1CyV
sT039eyBbCAq1SALqQHg12/Xftjyp8waglJKv1tCdC9NyJkGYHwPfAJ3VZ4K/BWB0mO2/0pnNGEc
CoKI28SnrFScNRyvKPowggvPa09or7fFN8af9v/hn7AktZABbllivpyd2UohUbE2qQfnl/dbXjOM
oNQjbye9haXEZ6hokAZEia0Nvtz+m7r5bkeTUt1jwNtJU4C32PexJgeS4pA/xgCRAYZsFMSP3i7Q
EcgUJ1uhyFdJVbFMQ80kKQYJTUK7Uaim5XCQ5J1Zn/QALxTFB6QV2Tg8+bJWPrxxgNBA1/moHh9t
sjceWEaS2MJgnxvbj7O3TLGaUnmjroEOyeHdhIetRaiLzgTCU/w+GSVQQPjB21T1UAgGc9bdyKv5
CZu7ZrJmK2/WCYlZFc4Y3WCDjBFvhXOW6aqXNI/Wqi5wDu3fzfiOmERHJuv3AFCB3UbJJNMrD3fy
JNWY1U6yNKBkm3u1vJrpWhGt60tU0hy6YAWMmtW30Yxr3X0pDjtT7mpQXOJ16km+QQAyl0b+W6IL
NJl48el3vfgAVk5j010pDO6bFS2OaDSSiNBV3tAzXedEkVjoyQR1XcILilSRQY4lXxvMrrxB6h20
nFWx3Ye8bZAq+pMCKXUuAnXPQ5Lkle7/Ewjx3y1+LA5ibFhLQUxn0BVZWX1A4c2w3yBnPIPgq+YT
1fwgJBYFH6l87Y/HN5FWFcYTr0+Ushwf4jQRKSKQyxyx4m1dLNre2wArotpwmH1mxwaxeXI2Q2CV
RgI+YpT3nTwYJJ1GwDAseOWQlK94rKPCfAOem/zyQGN8FwznJWoE5tBJCPwjt2QvsjpJMcuXNX3l
JUV3jHI/4BuVnC6ImSDfKQQVV5y0H3SSo0mrUSHmAmb2q/bzzG/rfh4LwG57M/CgkVnVmCb65PzW
Q5g5+ZatA8dxoCiHLEMAOuzsXzv1sXzi6wvpuMjbMPUrGTb1mB1YK58dx0Tfsg1Eb1KjERgBCOzK
jEws1HIURPmRPG7yuM31bdtSc8Kfj84UZVBPmVJz6g7sBiBiU+jCZLfky1BXw/JG1ls2Hr/8qzfx
bqW2g9xXu6IH1MocaCc3jVRwtSYg8KBLk1mJTi0WhsWU+8mmDcVFv3OvMTjkn20as1BTx3dEdloC
IjS93hgFeOdmtTgonTZvS809wr8eWAuNEZeUBrUDl1NFUcOLcBO5Ma6Bisl3Se06sMbIUO7shmU6
QRMIkGWp3r1eCLb96T5KzK1GO+9cJEDU0E1ZQyZcqV9hlwQkfHNcwR0IQF/1IoPpEfpJ1NVQ1tjw
kdxg1ZzLTDBg1dKYzadVHzjD6Q3Ip1Dh5KT5sy3htao2s9TSZBJ7tTbWEnfQaTMeGaiKi2QI/vhd
U9/vLuxa2umZFlayOtkhK8oqAMmu61H0VHuGutg1M90KV5kSMudFfjvNTC6ZATstB5V+fE++lkOn
XPaEWKKK3XmWYJHjESMIPojpfiIeP5L5F1NTyc2R2ndFVNdZigxrzntxip1NNz2QHbVJatO+VIWA
ZcXeW7J0N7gNmx2sW3aaBvu4VoL1ml61UoPjjR2pRc5czMk+/nGfU1HdFcdxcRffVr2xDfyPPW5h
HRf6aVqzzP4VM0PQkk5eOHGTsCzeJLbQ091vaWBCpgaGHMlKodlB76gBYnerouV7w31p0VjCIXFy
Peba44mzLIQPAh4FyVIdUFSYMOKjxdWhvwZoS3hoz1wHQl1/u4I6ioimR6W/8C2vwKKqb866Qohp
J54cMlWulKXErQ80jKd33HKE/maBqAapEo3YcQCoyDARLsHzUY/XBAkBx3kx6BKzEHQY4Yaa9zho
1zcdvRWUJO5T4OGzHa+GitFVz5iAymMPj5+hwzwb0NRq3RS5jZaX93X7eT7lIBwNhlw809yFriRf
F4xZUaKHpTpdqOBkBXmu4JzUFQed6f0UQ6+KUxziUnqU1BWkfnMX2ovh5eEg7I9BdBn3D+RehRZM
Jd1eW16waxoVqPxKgwdBls28NfiZBeObYt3iSTCCnqwK3oL0c+2HAgYjaRi+xu4QnCf+7UeYiQYt
Dnzv+s9bBLX0Wk9pXnw7ofHIzrkoqp9T2QxWCiCjf9jOBlJaZal4Ld2vb+eMvnCemApGgNLPljkh
uYrVofutsIQb3gdj2CoaSZSb597woqI0we9wS/tnQki4MJMDOfBN41D5cxydW90onQg423x46kk+
DJ3GGvfDj6XyvfB270lo+n4NP40xJ2ueu1SnppjfHGjOta3LYrBKWGlNo8N7WBoyqpcXhYDZ6l0D
5oz5EHTioZfmzrbSpikO9AvOWzfq9lO7XGIcbCRR1Mfm8QQoWSrsW6fYsKYJKva6vOuhtMoJMyES
Lvz/tcfJZWhpr5sS3EajpgiBD+PwxIIMzWKshZE9TWHLeu5vp/5C1Xv71BbwdZKGk6BrouBS+VbJ
+kjXzlbiVWd7XtkwUgQjpJuYjwLZGfht2wmAZqIbG3DLE7KyLfN13AG9WByH18JrTYbAlyqP529X
dyJofpl+2PTeYrcdhUOXNC4SXojHCmvqi2Dz5wbsj9RpVkA1QtcxqMEPVuRRqVFm7gOuv9hKmwut
QWCLSpQ3X1gWD3jKsbD1rEJkDS3tHENcVr8KoqrJZu76zPX0JvQ/TW+yrw/5MJrR5+3ld3AJgxjj
2kGigYvkXsav15OgBc3vWfD6PE3mfbCRZgoI6mjYbK4qDHHV2dwjEoJqNu2QQMRI7HP/GaIenwP4
GGE8+BSXb3S9ZiOkWztjgMMVeuPG2oY2bV8iap3EHNH8ZcH1XIbQHcmX6yibW85dsxWfBRN1SHPD
EHYY6P4BI9fMefmIoq3SAoDLy49xkyfJlLQjpIB9V9yITM1xZRLWoGQ6IaLLv3uQhFb2P1PyB4BV
p+f2C5vTrw7PGH1uw/VrINUGAECxzzPunZJFsJNvwj/aiCgy6STBfV11K05YGeOE7+ifRm4Yobj/
j+4tzF02qT2/855LN2kcdMSPJHlraRvDQ1jIrWY69fk4nMcxpSpfIWjCNlFjg19zockIPl2wNOL5
Nrq35x+PiUSIR8fqw7DFjw0xSCbwQ1sSdruKcGFsX6i4tGZSCTD5XRboNiN29avzKxcMF7cpkS5W
iGLFpIUiSu0IU1OHVDrwLDyZorBGDTLemYejDNVQ9dh4gbIcONeVULr0pPH0W3F/t5q4BfEAoZlC
AVc0B6r42LIR7QQNjBAE/hT8BhChFFC2Ue2qfBOHJ+uWzOJXXY+ff/tijByhJGEIuRot1J6IUCX3
HNnaxm95A+8WUrxcHl356+I8m6dASoDQY61T1/6/0Rk13mBt3QxaoEmE4DyqUlha5o2IMgOaCcWZ
RUjS4qfA+LO+KBml3fOD9HHK2bLoj5yOKZxEMLOQBBxlfHP12IWtIISqiwODpkWH+jRvDAzfdMY9
A3OnB7aWUvpmN7ylEGQ2SQGiohXm+kfoaR7GOyCsI5SprpIJDo7EzurEeMeJaCdzg+ZL3UNIQaVP
uH6NNGAZCu5fRutdf14vytCEw+2U/0u7m6fQO+wHQ/tKo9UeTNwKsPyEvri7B2ZHhTtPzo6Dub94
kk716387/wmuNwoSZ5o2B87mQwmG8R9z/wnZf4ZOGwTp91JaPIK4HDJPS+ElIpWg1zVQ+oCo5t/K
FNCBgZKKKjTrE/rYL3c2dEhtlR2ikkCaRHV/CkQaoAwr7RZTgl1Kk67fYuSHQoHKA+8pVox6sMt2
P3wCisvx/nD0H9a6a4EzLBiTHuqpo/7Wi9dD6KpV+eybuqahrSaRCLcfTZr7JIohC4n8AZNj3AcH
hAvF9kkdoz+DmJPVv1Ncl0YRaYt9IfhwCkIib07g2/oNyAMx4UfuTabfOC7ep/UsrllZ+lzABPlZ
9BlCPjE+EKiV21578KcKtA+qinTkdkpXTh7Oh7sIQsTIaWdwybVle7DnUKSCy3iJGAW2Hgr51nJa
fqLE+lrFuuG+F1U/H0lIYvMrUvRBI34X81JT4eUmoS8flQqNSvztX+MUIyEKOJh8kUQEM0QK6zT8
S32pyVy2jNWUazRY1pMBwidakLYWxh243DupDEzyD8QEYj3o+Kiu0UvCy/gl9aaXE8QavQGNLp9t
hFpzIe1S0xwqHwARXbmeE4dZ6zu0ZMsySV9ACHlSyXiUVG4HthC2vC1zazwZpgMvKdZUfXP0PoXy
Uo0Oj67IPaLmhUNiD/fussGnd+qw7q+CEjQAzxuMDYREVLzQJ06HsEMiHN40mPxILqLt/Pu/vsRL
YcNTCANwo1iCoHwXOJcKZk/R1pmanPs3oV+rKP6TcNqrJbknJeeiTwXC4+qzQk7aBvKkO914Z5dS
GbrNtG3G//xg+wSSpSEjbtvjchdDR0dtN9GBiARFunaNjvtydJKjwJAyAu0cDKpYVaJTnxMM7HgE
FbUOKzZnDOrlQbIc9AKG2Dzr3o2WlZUFvobbGlmAHrYLK4BWplx1Bcn+5Ac09ZkRTdVxn29ny2on
t9J65/9Iv3+qLBv4Mam3I8Y/lmQ5JTVVSNm1Ir5oQZrPU8zE0SPIr3A4a9xAmijYh/mYNVqummsj
WbpdOfLb/jyXOcZLAxQqB4eiSdwLujhfs/4tf/GNvMSbeCLxdRTAHlfzYpFeyYq0vc7wNVxJs+P4
u18FLaLM7bF6CibSG9/l9RFc9GhBnF25DG5JQFYg0v2dnGMIpqzRaSoJWXwFhWBJGifJnCpTq+Kj
Z0VxeW0oNWSOluh+47Sbq0OpIXYxVsUj1t7yLhV+q0hUcF105YkCdidX3UMOReQLaGEHpJEMeOBr
XBH3rAX94nVYtWmU+NDJe4V9fi7nhaxPFIpL65wNo/7TkfIfmeeALjsFoy/yoPnkwaLv6kjn2Fog
nTgvXsnTttbfNx+CrEH5gnI2xV3SM2PbqFj+GX96MT/XBHdX7bj55Ss7nhxMk73vHMaN/Uoi39z3
+lpzv5evddGjQtWv5ZDuF/APkeXQw6LrrLVHUCydcaHd9gcKeS+d2M/R6fkJ8ofdxCsAFpQEgoHZ
oV1/l7oIknjoMjHE+kUaZhN8/KFk4U/UZz0lN3UEDG+RkCZVzsG5xys5Tm1slusQxmhFCSIjeyD2
tuoYoQy3haTKYvu9wowUDOUZ6wCT4m2uRyFG3OGIRG+U1RjQhN9eHKRstZitVMSOfjvWJjJkC+F2
5+ugrPvbCYV9PX/gDGai8TYOv8QwmCwqYku7/UOOCB8ttsgjKQGDOCTFqnUsPM3Aa830S/pK256T
K0Sf1IasgaBGMcaJBBs7v5qWPytNSRm4zp9l7Rt24bG1Ab0hb6+oKIHXJYuyvJKZDAmjNGIqT3hs
Rz2FoO+nstBAA/L2mVyYonf9zDR8ATMIlHmm5T6Laot0JveDI4xb5Kqz2qTnAQrpXr+sepJ8ffAD
sauPxP0lpyRucnfME+Me4CjgyXoGanRIST95DBDRTaYhFCoHrNiZPzjuD4MnAo3eyosb6PRX+Kow
ghJl1SqAZ72cQnzzOEL6B+2Dvwo3OvoIXA3qZZUhHvuJAMhEXHa9pQR+jdEt73BLVblvVW4T0SRe
fAXapIUoHqNQi75HothlF8z0i87UTW7WVrmlodHi1CergIKkQ4v58IbgYbY4ZWr28K3jW4qE5QY9
jMLH+aWSkT0YI1zG5mVwNcUtShD2wz4xlfwJQ4cl00AcXS4VXdFYqqYtkskCsiwVesopeHvN5WM9
wDeLS53r+Zt8Qsheqr4g0bupvtx4wNbIHCrBghZ5cWgqRl8j/flp6gOSvD859Oe3Ltm9uJIGgxhe
ii8D4eEwrpzo2RD924A8y5zVQQKIv58nugXe98PEd6YJoAuCwwi+wv3/dh+/BRFnYupqGTSLfxv8
5OkUOpliAvkYICIQMag9WSehNoVbXhALH9sti8GRDj9GE9eatcY3jeOopIsx/KxHN4ub3cip1Y7q
+uIvCc2SGV8OFqYXU2q7eSelye0RKLdcP9L1VKJvmMCPyCiMl8v+uhYSQzF1bzUFpZ24SSeLR+6w
WtaOdAe08rYcg/WNSzpAyrYpvVZnhL1y1KqOzPGp6P2Pe/FanLcD2vCsRac9urwDNfcyF8j9hOsr
CoqQJSXfGQ0u9rzo4l5+wyGdmQF/E7XRXaUbrqHHrzmtqWWvDL6Lx/IqAOyHtHlSQV05rX2RGuDw
e+lil3aA+x55m13dgSYddtknmWsZfkheFbCHb1WMfWPs7ZBikNhkTPE7BI9DczWa97N1kE2ic0R1
zBFMuQGj6vkALq2Nv1hsZsztDf4EnCzWEEQdiTslBB7JhCZGsdDJb8Qq/EvivH5NsTygBI5MvQcl
kDW8D2W/Jp6FwStYv1TiCUr3ym0ws7RqF/m3taOV7DWfXJcadCmnkdXoSMHYZRYHIKY64h5Z/y00
6NWsEOvv5nxJlK+9bLe9hng5DfkfxKFrGeUxYYaz9YLN5d8Ty2mzx4nyD/zMHhqyH9QcXFj2wDGS
5WFWmBn9lPhqjeiv454C7pU6ku3tmt58GvHmslqKWotbWAZF+PbH8YdKJC2guOrd8ZjMq5Krf6j2
aCb27GYucMiCGuCwGWNcYzyOLi9puDd0BYJOmZEG+Dzr5BxN7cVizSUGIGUYxnql1ev6u0yeOqxx
qr68dTjO7lqVOGIG6lHa7EIGFLsr01tKK3ZS8R6GCI0nJhdfVy3t0w0lcmFatGwkBev9aNO7EOKC
YC6CBZ/RAhfgVjJ+Fr7vjCf9NvKNklqBlAaMvibcT0+hs3B+ArhP2tNdjZd1RSzhD5wHeCMrUO7L
Dds33PvIAmlf2LwqiVjpgdrh+2OIVnljZ7qriXm3xsg7f7WZsJ1aK9TTDRoIMhbLGmU3DWL/XjrK
jKr+5LeI0B0FS2xOw/RTOsUDS8Duh5UxFsVf5Q83FX3hhUh8kOBR/l2pqoQQVJOXQxho57lokXb9
lDU3LIFtNHG7ehcX5isi9F/bUdM4tcDxKMaOmp8x2akQjKPKSFwPUfSy3HMQHq8TobdFu4CG+YW6
Kk97L5rsc2ipu/a0OUljwv9oq/iJXNzbl41We5seMuOh1xlG/EGs3bJLt8GVhFyac+vfLNSq5vqq
+UR32ZzdwlbpPOJ2Zb/y40y21yHGXUXa8llLHD9KnPm807zyCQZyJ/fo49D7j7ixSZydBUu/eQoN
TaE+wmROG5ofkcV2+4gWG2+5LeE/RiHK2UNKPrc99Vfjw0PFnnP3kPqZwAqXdfan3Pxe3ntIQlDS
yrAU2NF0qeTmqypimRh/0/mIY3tO2dIPCUmiW8/m2r1DkPpNZCSNhe1jkpq4AGf45I/kb3ZR7bqt
NmspiMqnMPfwe5fiF59ivQgOp9STrVLo7xteDqyf30h9PAMWPptZH3HMZGfkD/yfEL1KbO8zL36t
FYJ4ydYbGmjFLOW5PzeFw1Y5s1KTwp7LVhLxYPOOyxHDbCLrdrqDCWVzwbYV06Svy9OzoaklCSCB
flglNJyIwo1zHVlA4Ld8KPtE7LFNbLZ47tDVu8ZwDtvxQa/hgji0vukSvznZelVXLRKkHPqKsHPg
5Jgeh4jQS12vodgdQkF14yD1XotOL8aenecEJW7+4r6faO5gXdYOeaceNXKfAIVjfQigJ09MFNFm
hWrCc5FPODQi8TcYkPp873ZQzX7lQoEOchO9gbY3dVboznb1s4YF5RIxFL7br47o72UXB3p3vlqA
j+LbBHUo9yKTTpvHrq3EK3OSqT1+NmMSScumE1ugYiEGcs7/WYRPxRMVyq5JL8eLrQDO+ioKwyZM
/h2KpF+YfoOXvmWEfg4A+xhMjN9qY7V8vjlrxapS8XU9jdtRpLPe52Bt08xaOPdbbADcetoY6ChM
ijlu8cXkTjRRjpqOqnOa2k5e9VS+JFeE6ELkVrQiHAxR210S0RPh+Dk6N6L8yxa2BPKm6uiXTAuJ
Evdo85QCDWKpKu7MeXdmj0TDNFXRdOEdVJD2HLsQ5i03SK4CK0ueRpUBGYEIqFEHx4Y2O0gXUWTo
l1PNxI4ZJIZb93cNvBY0bquaTBo2SCcMH+qnaGd4jh2AtIlCZOE6UHe93J2XccpZCTIgLJg2CGng
oJ8rUeSOxw16rKViVWlKnhRoZr7v8f7Tl7RNFuQjf4V7JQST2Z/NFswupdguXkcvyn62rzZc2sk6
0SlfQCXtzdafjU3walj58GFbubissJtN6iCiHVsGTapxjjPo11zqeJCBlF0h+64lBpoJJ0JxYJCF
rik6rL8sTA3KQdP12vbmYFf+nJHLIJ/IOw3EIHFsu2WK+5KWrb1FJY6bj8ElhBUGZijMMHHAXano
wJPZ5t/TplWmT2/R98JpmKpdT78uhYhDYs+xs5n3EBKjYGLs2IdrqnMLK/QutFRWD+Wnc1mEVeTW
qmefIiiDDRSQ9V1BlZ7MnODwrQjar4jb93/QvYYQTBHoOLtvtuQyMDvLNuj+PEVQQqU8ztavuFnk
eYp6uoltkfRZhwzdIZe36JNl+UAIZbx466pkHg3IUd2km5544A/ekt77DIK4fxRUTRE+As9B7iOm
7njohyuv3Of27+G2VhlmVnlkLQamjs5XJj0EvEoa8UZL9uLaSwkWBm1V0inVRKrPgI9e2k12TSFS
xOUczfbxacQOT1Ipdxv9AorhxHCi1laJkA6xg6Y6b1ZDO4ojX9ftMtRudweVOLv35OVXC7hP94xK
7u4u+MJSH+DOjZiuq6UvVGmU8bDJfaOFPNor0Y1tsDRhVnUUinmjkm1K6tbkdDzh2M24bJnw9sMy
oIqOgRQA3B+Aecepzw6OeGI23EuNfjBBKjXKsV+wqVhChLwfuB1ovQtTDhP0MmpQpqykiC/PBAwh
L5VgpNVaoJaPUvanVh8vKXNBhoardNXRxOcB4gAPAPuKTC5qsknWgLLuEZzCkL/0u3WMB3tVztyB
uShx99RLw82WDqeLqw6p9Cd7F//XWWtAbuHQUjOqke7iBg4Uc1pSXchSFuPj70ZfWshTDfhz/4s/
A+D7LC9m3InhhrlVnU+OaBtLPSonQ4eOFx+F1LHDRGjXXKIWOxwv1nSnVxnSHYeedvX5/Tuz0CX4
jQDTd6NkuewDVJUCCdLZlDlktLVMlNezD1GH7oKyNfkXnfQGVEEI99qu4V6ceHx3Wi2kkqgM9UIX
Wi53pDU9SWt3gTNpV9cYCxdDOkoB+aMyp1GGJnvOw+wUFeOWDDYtakN/W+bya3jVmzsG4mwek6qe
v4jAkX1uSnVUDQIdYjjkVv6SCXoEqPc0ORLi1z8RzDnwTuDhTGGa5xBReZl8uf0Yrdkhj9lZk8jJ
0bAQ0QjhMkIx8fqBe/KqJEk2Gwr3ZWHH6Ak8oH0EPa/k5Yo/Rc+NGVMp73YP96GwYV4rm1I8Zc1W
GrBht/t7TlkdlvRGmMNZBf63TFo5QMf5helSr0p7wX4/xx1mt7IYBhFBkbckPLlo9pi2N4SajuZE
LAqJ7wtLtt5tqj2UsQ5xOUAbhgcpiYWAzdpL/IvuC385hMFTT2UURoirY8QQh/tOPB8gLP9Gjjhf
LAPmGJnUqHHyXePRJBZ4EBWT2NQCjGVhgF4itmaTdg9PSXX71XBApiCbKkRavPyLcubtNhskU9w0
8iTrYlxuI3e++yjnZhe0j+56HhngqtWVQdmSbxATRnK1Cz8d7jcpwVSH2JUSYb0U5WmVJDeTZ1l0
7RhWcKupvZVVAIP82Psikl2S9vY61KWvA12f6kx7VsofYl8iarHnuxl5SmJwDuxc8jXOU5pxr/g9
V9PqWVxF04+fhuIYUWeLZJJlc6y7r6VG2UD5Fr/5lPhreFWu/Vqjo9gXSOrSSMZuxgVGmVZSX1Tq
sK/rY5fn3j4/ntwmiMnOtAKHADKtMEgtgnbr47MYBH2MiPxeBcJDQ3h4M7FrhL8o2dEhYV+oun1/
Uq7aBJDl9KeuqdlgNNPwSvtWnUkm0DCRymWoDHzzrBm/uf1eXO5BkFKSBAx9DJy9MgtKtCXkWlJs
kbEMicdkq7u5CwexCbp47Fs31TaXbcL2S7LAD1/SXT+XQIUcpO49Upx6iFNUle9JyswXzOHUBTmJ
0J6Z9oWf9ajClJf3Muzi4ie3QkYH13rz/cb2CCGFvZXI07SFGPnKOFjlQVl3WLjgE9urP65N/Bpb
q+/y6dpFgean1fLXdoPxV0JfFBskkqOxrxhrs7ckUGWf/HWNwvK7GWQl9pYF/5gsiGZDdPMLIZa2
/lBNUWXYrg48g8lAnxk7Ljx9uo8lI2fp3MCJqlCplYA3at09tx8ea2uLCYt9mpX50XUEB4/lZTb2
dzAhs96gFmrXbKKeSpBYdoI24FllbXJoh7xXfJd53/EdCOf+q8aHpMWngTrQDIKpmIkkzwg+kZ/8
UZFnAxxhqx4f5Hrr0ZRIU4+2+fSZkbDsxHxldCNpXQU7V0Vm/I/xyxmgJpzJrsLD6yuira9bn50M
YU6uiVh1wImwoCXS4m1UTapW95Nj/8mobTp7JmvtAPfDQ0VdQXQgh+MexEFv/6oGRBpwtcHahGov
7c6EayeijCAY3ptdES155EcI+OHuUOceHwVej9JDZmoCcZRoFKnHmgJSix2i8ErVtgsrB5XZUaHy
QDEx96L9Jki8oHVf1XkSkEC9J31wwmyyd5G3mOeD6aE9LWxlYoW4uA5U/bepEdY/iNFQdZBjgDil
dbXUfCqBk2sWUCYY1xCPuG8VBGj9HLI+HODKRNa1TT6vQ5F0cQMOt+pmPFZvjN4N52FeSIy1fHj7
hDieg7qDUo9BzRvgrxHR8UgJyH3JP4Cp1lbtVU4Nmje8jQafsAdllJH4+Y/9g7SU6zA7K4F2fsVO
C8FCCloK7+AcgiYDVzaUdoUd0A5fHK3bERJRHCIy7UvRqfA67jsuPDfhItAosPtN8zDeh5HxqYzP
p924rQ8hPYYAMrJhpiYduby6Sb8eEITpQ0+cVDtTL/N0h1Kgq+9OUQuDs3O323iSXEC1Wr4AaieH
IdT56le1BK51nUADZC43vPtZ/qcqtNaTqZlhPYHcfd/YrKpTRQCekG1zult3XOB4Xj2jBmRWrGDc
UTVau4P1Fla5nN3M558eXsGAH8Tk2f6xmj75I06N6a2icS07nKtYOt71cRS+dA7LnYTG0ue3/Qf3
OSeFCYGfXxdNfpUm415BtDN7nlHEGAH2yzopUwe2iLCufVFdrnEfdgyjM5oiGy/4DNG+Jcl2ZE+3
ZGVKEVCLk8hCL+bFAu5H7uLB4WfEJlW+Eg3EiP0TwIkCw9S9cm/yPaieLx4zW0LetPaUcfF1iYjJ
mhotabrnmg/4HuwOy6vUN6mj1Rm6/yN7ygbrJuJOGmRXKwuMlgvwbbKgcQjNxnBHnpra6uGL2G20
UosZ3EfXu5Zk02zpIA7Ld2I34uuQL7RpaKUsVIwLLhP2OdDW2WUlVVJ4rl/D8uPC/3GMRfE1ZBxj
PsMUNEk+FdFcZnKxaz0WtOS9lI7TUI3PsIr6MFnZxYV1Rh8W5nwSDbqkngUrGvQQPPsX38cwy31p
+GqdPlwjzXob85hXZGtPE6ieIIe0sNvAoHsXVz4FW/LnKNZB9d30TivNEMYB1fjMagsifOoIw2yp
UefR5d/LjNKyyARKf+eCZLp6LkCsX6WLWKp3t7AkFtooNeC2CrliHqD7u+707eQfyGjkwGXO9KI9
AreD8t4pWpkDIByillwgQ4XVpxW+NUrHk9lmrvW0v4zJmeQ/pF+sHi2HxDQwF5ncfpVDhYJtw6rq
nfEhliF/5GeJirsfsCJtu1XxaJ+cmHYS0j+CXuGonGeeWHl5rR39GH9hNN5i7Mc43KpQor7s03Zd
BbNQzIruyC/+T8W5Nwd2bZixdUrgPCvfn3LT+BxPRx6Jq17JUG2ufVFGxEJV3oUmzz1lXS1g0SrZ
0ZCWj9HRE2jqDDgWLqlwPgLru6uxB/K+74/gGVXoyTYH0Z0z2TLdwF4+Wfc/0uS19MY8sT6GthnD
MfmPYOhnTp8SDgJp/uJ5lyDg6bT//++AXc+x2mXD+N25akYdbIsMNXQN0YlFd4fJy03yJEceiEsR
crDkUct9YXd7uZqIIVLvW44XYPj4RDDPcYVn5wsK+83/VkAadZXtQV7ntYWh1qNFiCgdRoOm+oKR
HbDY9cMwgqRER39ojcCiaMhqBmrV+1gzxkUzS/aBG6kiBu+5hoacjJ0sBoX7dEYXpbpUArVj6wS9
dMzS2gAiixofRhDv4ZZXqtPUZhxnhrOtPmQhAWRrWgIHyRETd9DKZKQ4AcpocPs6J3gO2hMziQaW
TKb2H6w9iXDCInpqfjXhyNQ00GlVhanbaYSIcCVgZpCY0wXV5AbaAu8Kj3yqTt44x3Q7ZgfWtmgv
TjWsp2hJwGMPE5EsHFT+sKQOzpslyrg9aqVSoxSKpkl1ORiMyJM6HKI4NmA0gD9+uAaIBa+qZQSw
6tavbFzpa0diRujMMpF3BCQ017zf36uPNRN0zmMnjvMWjjI/1ZMcIcsxg0cHYO2reZDfHAt/avGR
Z6NgSFbhumzYZUJ0jZGS2K7QshZh2KXYorkBsiXiwixFqEiDdvFht+6ra/OsyXuknsWUnOQsCjYV
blIqtsKTgFLu0EHvqfpdm+S5RI5bBAlPl1kB6QlPi9IN0cJt6Rn5QRat2g4OKjnf+UdPWuiVOeA6
fxQVrz4G1p9MzaeLQdjjWLQ6AII6PBfIsChjjgYjMlnMVpvfMZW0CJYhlw1ZK+QM76zCxB7F42QY
PClwLfN0A36eLDlNTjbaJ46ZzGGKOY0AFwsBowh/THwa5Y14lv7XmCko1po0QEfN3EMhrGZwzEDR
wbpi9kFE3xYsafyvWpHKM9cYyb4pPTzEXOUJr7EcFITunjy2UdPQaKyhzf1xrYwfV4GgZeHfCyEp
lhXJ1z2UUn0A1Haq1kjq7Bc/x1frFzjc5gi0mm5V5NN4HGUrUJRnOk4w3VPWvLvAbY34wVgzAH+W
EMcP1CzzNTwgIGSBrXl59SLmLVncG5xMeniTJ8NOLYUnWg/QJ9PZzPxK+A4K8evKZHRQkY27U7PI
ti5p3kBJVbKWeTvBv9o5hmu4G6AEAqlErWoZI+E+8Idr6OAOufCa12O0l9+wD96kB/ZvIedr6llI
JrtickpXv5VccOoszMnDUcL5zpYAp3828nFQ4lpmfD6BHmUcI7DA3rHyVGlaIt6WSEbMjIuf1wgC
qsd9LjHVfcOSekxV7Fny3VGEscIpMyeEIBoR3Iye2od3eqJcz0mI/2wL3X3O0nPeNQJwzAPG5x9R
q6M3xPH1NXdjgekpO9El6rL6XSo/8moysthtmy35Pc1gljWN9MPQ+LF4E9t0Do8V3TFfSvOWfk3y
rKeZ48wP4azLtqIjqmzn3+pu1AXIqDJXAA+icCbL7B9iilaIIzfoQggS19m7EYhvrNw0X8AZ91N8
Lx02UQAeETRYiTKUaHvkyp+/Y2jP6qvCyEZrdduXuRNhE+GHSN4B9lBv6EAKfT0k/dCJxvQ4ZkwS
kfPWY4WirrTDGMEcwywWvgXa3gvOolNS4Sex3gMx5mBoJfUAsyIuJyzyYlsypmXlDSqJmFD/bAWH
diGqN1CGGRZsAQrnv1Ca3Kyfp+yqp9JTzv2+hPlk/ZF78TjiU68eaO0h2jAxyu2eUXYS043NKvtb
Z7G/lgjtO1T3vAHyrMyOpPKlx4/6jbfJHxVFksy6spI5P+LxRP//adZfyBuMyzTVAwgepUuTgUjo
FhtkyI6icHZJxt/CpV1/Bp3U+LMbBBy1dloEIQWSWDDBP63DwcRjjIgVMROMidMuS3RqZ/U1nCsX
5dOxAQh8BLBUbUOTw59MpCkuJcy7+blaIWpAknl/MXHqZ0XMl8KhHngffCgKamjyrhAlW+Xv2wvG
PLroClMnePCyLtXo4pSFgdKF4TgLgicIuZieYpfXXSQXM0ftKq7zDnM9mnMTu1E+jYE9I7+2LeR8
vAarvXrDE8H0YCh567g6g9/cEKXvC9u42VvStaxDTQMg6PiMalu+WNOaZQ5Esu18Rt7hS6TpnQvN
LLiV8nDtZTvSu5oD1jpYypyvrpDTNv1hv/au6cZQLMoENQJUMdWJp5Bxj2W0z7kQJFWbUXM8g5Dp
l8XZ9BW3GwAMBh7A7frDUuzHrzonDS+tDdiusDAYR2Ivc+3ZsaHTVJ8cxTcPxAAjusC9v2w+9PGU
eAtY5vSUDI2tW4tkpd80tGbtzKu38t/cn0iDAISX42ptHjl6kD8BeIUR3WIcNKsBSB1AcqZhq8Bn
NqU731bGmsdgQxHajc39aT3ArA/zFEpxQqISaOcDlh0wJfftxSSEwCCwoQMGkWvaK3T91AWTJHrQ
M+CtUDdYQ0kr+15ium6kYOyBO5W1uIQe4rpma0mrH8kxRl1zCUyzNh5IevUjM9BY4tOZ8vfXs23Y
bFAkmyl8iBNlZviJ1RGNWWyafQHDOjBcUJG506HVKy4PYNNh7bS5C7HOYRTRoTIauS2J3Z3o4/3/
8SF3wgGPvxROVg70nom3/WfIc5/z/jGDSZ5ELTk82Xa7zKEwdi4Zx8MIC0i3ae30EiTrJ5aJXHuT
sT1F03pNIXfWXpIiQMh1kkKdfWmfN/5uvI9lCDrO2CQrb5bh5IgiMyHuxAzM815mnqPX3p2sPgFh
FSB/fUiw0M9bD64eTX48k4X93PTUCTNrHkxTNtHJOMaSJa+RS6EWBsRjdfRCFR6vh71IrE7UeJBK
/Jpq9a65td+if8KdQwLj9AIlv3o5cS7JXU7mY9LFb9ypsAYANtGmTcsg4uXutl1g6NcGubgsrxfl
QegdSphXu5gVP0flkDWMtv99SMvhPn7/K4kHwWzRsqqaR4ceLT65jR2XFax7cki3FbcTQOhQs3lt
kskxB0DljDoWwH/O4OwpXHkJXgfNd8+8QR9f3vZTVOhGRoSLaSll1Sw+5brHxAM+gHvKTwbtaQct
2cKRGBHyxhlFBMP4XN5vO8CukvomeZJ24WloZMBBPGK+09qRKZk0K6s80V8tpTOpxucrr6xCDMHr
mIvHX3IlFwF/sBsjsjTGZw4m+oqr8QLfOmlbqScwAM3B2Hblu3BtRD6BsPLq+Fv4+gTV8Jx91fp/
/R4+j/zFzGg6SgRZS6CB/rTRyj73ImvZKF4K2Rx3Mz5d5d0oUBchbO674bvwXwGMz2TnHHKSdHfF
qIjImr8qos4Ri27lh9ubEGYKDdldY14LToIbeUJfy71N5vXCe6iVdMBECzESlMUE+UFSbk0gyI4B
Mbttusi3zwgi0zZ68Zix7TFtmqMlFsym0bau0JWMsk6Fnd9GigYoQV04GtGRpN1XQCMoYaE2SViG
pNs4Q3MG0NmTy+HHQ0dlL79NFwCYiQrRbtUizcBAdWyIhT7n96n7WRrj2E5lkEwnPihSsgn/4EVj
CJELKds4fyhwJzXzTmfqL5Dm17cRWJ/sJOHkkNM8wmZJ2mI6K7h4yT1tbPMmCZP7Nrt71UTmjbgZ
8UcY0cEYxmyI8Tmq4N30S97KKSuvxnnEHo04g0KCwg4aja18xqMjk0H+Bin0s6sdmYGrxRvp490h
yQNJK7bMBAM3VVX7k9gFA7Ipi7bToW/lMgX6r4ZKVDcVc3OFdZqGk4e+JTjPnaavn8Ey59l7w0eD
crFOVj6/nWwL9LYWOZruQD3Y/jxKs6PDIHDsMGJqCzC2vF5nPgPV9vz5BwvrtzEzpoh17INVt+d3
0AhzWk2fvl+SowfrnEgyqGzs3WgnzkQFTO/agb98aeHM0uP5cZc0v5Uob7WAor+nDD+Dx2SvaGyz
GP6tvO/eTTWb12VWZsgxoj/Sl1XQHzmbb+vPeAV1qyRjRDgtUOS0+owaiWTZ2vhqBCkpkLyr5ep6
rq862uRGj4JEtyV84ZojELTARHUAUwB7SZu4NSJ8o5w1i6iTJOHqpkd20jOKI7KEnWXXdnZVLd2Z
B5OsepgWgjydf3hdhpJBxS+ADkuF8ECL4idggd/FyovHV8yDbILLUE7c10weTGm8TWzWMYpb8c61
u+zRXGDVAQgY6O6eDnGHyyom7MNA1h4NVgf9n92KG3jtJMM5doeFjPKsB+6sLEQ8wRvW8hLbd3n5
LUgpu6349uirX05lRzu4XNzYPm2IGnoQJPGl3FM/Ht8CRp17HS9CfdT6WDt4WkhZfqbJNsLL78QA
laPPUCvfjnj6clmabbJXUB+PyTGbLAAogiF/676rVl2ifk89PA+P2xn3Gi8C9F2y+J/SJrJaMFVd
bX1anPjKiFvCefy9jrffJKe4D4CPpm7+HFcQXT7Oh6gfcUsduYRMaBxEDwn0/Ugn7bfJ9Ss7/2HM
AdaxvESe9/7OQt7Il5CLL0BpYUrnlhs65V8uABaI7TbSE8BBH2ee/61gcAdaT7Q450ahCnvyIt2a
s1ARkLw5BiWfNok+1O1FP8bLncJGBDGr4w3GfujekLfUOK+VtBPNz5aZwOVJgxdbi1hm+BPwbpLk
PtDKFtoKqEoA2TOzdgMITHtR2bx+Ux3yz7732NbOZS/Hp+QzP7tOzmI6NKYNySLSPGra5D+59AHq
PrYoi+U5UJwsqGzXukGMTzkweHNBkBQOdINW/1ARwRopAJfBUX0eBEHix+4i6J/CYgduL/vdrcvx
89ySTL2TUShNHET/hu/YvefZ2C56UwTFlaX2B8xqIhul16BkapbCVooK9Atf4dRJHOZuco7ZOgc3
XJTSKYBMdOHpbY8czXtLgVYQaZqkmbLy9rB+7JGAZWfJY61rUxUaZhbOiYV0c4jxuijBnsqehRM8
zfe9tcu3mzzFQvWZ5+bYHG0G53Rflx9ylpcPgvSCIzMcOJnOOZKjpU/kqy6Gf/zc1Aim10AhMo/b
6JMmKN0dwGitysnZChlbn1LgXjuWcZ44W/IjdaYhPtqJY0S5ym0eA599lhuzG0hQ0+Na92Z2rtKK
4GmSxImLXh3Hop8J92OXASn70Ow68YrSZC8vWxQQ/Fr5EQGWBTwf40Ke3bL//TJM0b3C00e/p8hg
YArk32tLrrZ8/fOO4zKar4buQMxF+nvvTsPcE5RXdlR8GS9DCZqmOs7GdXMu/YiJ86u1Vux6mqL7
q9zfkBERkNOvde/aEdFYQHTLRtkVXWLUi52vjBsRpwZrOsI2sDdLtg/OgjIobGL5gPp672yoIkcq
ERvVpu2NzyOCQbpH2btmwio+xFuuzrdxZzNQ+uCMkzMvqmubNOoxMvqKUJ+gp7uLOevoyjaJW1PT
IbqCqzXkR5EyofpLZhemT0qwlUe03bmJsANBGglX6TH/3KHC4igKBQQI0m0IRN84WjGYYJIffZcN
1+vmmAlTVHGQi03w9fHlNXaG7PBxCpbzCt165+64P8A8wtabWML2ACdLgq8E9cLYsm5UeKfLPWFn
unNb1pgf2EuAcmkiUoUVRyvo3mKkVs7TOnly5IVB987rzPc32Ge/Ujmg1VCWof9PEEfVqZ5BlF9j
dsyCuTgJLcZMteml4LNo6JjZFyZRo4rpuYj6oy+3YzecCHzjSFUixFeF+Yz0tnfuMPbvCdMJMKuK
d/uUhhCGbqKRCY2FFMHp19e8PxFLSr5EALZsdoHmQzPe1PoLNc96Ho2wdDVU6jZwdl/aRzM5Fhtt
074kUS5/OLzVYtmgYkbLRgab9YiiUH0ozTSw2aLIQ1mR3cGX114fNAArn/nfjaRxTg30tISV5qbu
dUBPqpmwaQOhwQCLiF1JL5THZrESIKpARLGsTENp6maCs9kUrd2iVYvP1ef0upkhUqpzTA6NvIFc
UBQmv9oGJ+mce8//NKBtCWcQXgfnluBzJh1btXkZ5LC5cIvpm1KW/5JFQmCkiXYDGnEpAslgLymW
Phwi48UgXbXX/s/7Edvc6YwXO+VSxkbyTknDOHQ+RFSUqOfdeErqh7G4Vs61/J95/1j2rZis8VvO
0/GqVbNER+yA7+f4bn6oWsKuIpcT8nsYiUleOBlRf2iXjcpAZPd7Ge1GXL7M8IPImI+i3JTpa2jY
8WWUbXunhYJVyezMg8wRp8FWicC8Ae6+B0IDACP5/I31i59B+oejnFXuhp9r8a/IFecDl0Fckjmn
HFdGUV19rcrfJZibu20Seax2invvDnhEU6HdbWlqBrRtYcyYdivwCa5zM+05GjxFUyJlIBdWm5iH
HgQpzaCAGdSh3lw5Fs60REz3grQ1vLp4RznHHAfNj2z4ry+hFHtqZJzUX5ne1MjH9VjUWRDPosQ7
CxZkoselmC42S3kuBSFmDNzpfQ3nxAOB0HEVfycE2yftHf66zTu4xtpqVRRd6l3b+pn4qoGwNgzb
+WYyCH7o29PTBJ9OZy0LwRR6NI6E7IIz5dCHxczgp4YZEIbI+2GFNrFEPcAPM5A2+fooMFbOCAcB
tLxEs5hAygrkf/FNdaVkRG0ho0qiRIAoeUyxUtMAfICDTpaEHlaZH19ssXiCt+USo2WVPKCldXcz
sRJWuQavL4an8K3LMX+Tv38HAYMZIB6BuveNPdOyxTabs2mVl4c2unxkiUPQBRGfBbiyL4pha8kN
kP3IRY+Rcv1CZr6AYRUyfWyv89shwtytJOJKlXntndmVutpbDIRtHVUMsg3jTVB5j9nLT50YM7Ca
bYrifyAjRNzgUiPhEC7ph0pjd7lzkS8lHiYcd/5EIVFjIVP29IrNcG8mW4wCZOwfLn3HYavMBmDN
sEiISew4OZV67mgUCQw1OVykasorfan2v+9fTbQzoNoiM/lTexSoqvzM6jE70h9UOZF1UwI0bitU
EOJlnVivYPwtoYncp/wIoSQsIOJjJhSX4Sipc/70YS82cTVtXFE3fInjQO5rdjZLLjl7P6KvR2x3
p2isXzEm/KgGc5RM4IxHJnLMUU8JmMxxg7U9NkfwmEPQ7Fp3MPppq6/asWYHVVuqHVQ5D9t1VQWu
k1TT35EyBP0TDLO7LP8Y1OhoY+AppbFQ1mTb+qd2zBc1HnEFrqC2FMQ5BP0zzza9tHyjp/h2xm4d
GoDHgz9xrjbYDs0YiV1uhMoNf96xnfgJ0Rfi2tBSm7ZuDuLKpcT3RjHB13gcggNhEj5mw53NLZe3
BG+s3i1aICTOcdMi9AXKdd3TO5eogP6gGhvp2ejNBVgLCUsNbaiTOUuTbSmCnawEynDK0fj5LYNw
vd4QwSVpvBLuCk7pFVVCjZ1rmeQ4pvsN5TcPlrme+roqV1QDJcUj8yL+acbpBvfu/3WGjqvQzbMN
NqHV0akGnPFOVBENsr60WmU+1RJZPmGSAVM8ASdk+pD9t5NVEIS5ImGD1UbudV5rg2nm3Omwo2zK
hsycGhT44RFqkkTiqhtEjaA08ejhsuL2snMEZ1OzAcyxpbYsChiE+2baJOFSVGGQBFNxuzrOXX6/
u1AEi34VP+rxqtfAc4Ncn+N+BgylxEe1Z4T91c7Oy7tIY9KHXu5pYvD9X/MaD9sOH7s0bQH4hu9O
NzyjqYXswGP8Pz8puqrqcRsyp53zOxHhZGmvxXGtRa4qBwELupXmkI77d7ZWbBlj2d4/fFG4+3y7
6oPMgwjkzp9RP/ZaHEUiS3PMGgQv/D/pl8VT/yWTCaC/BqxDFDTeqQV49z5EhQXBISGXeCqhJXh3
u/uYg5FA+KgFbHNebLWuVvU2ByDpCA6QFWgLpYAZDi2HJVIsAKlVqZsDbYz1/bt18HIZSnin+zLL
j9vnUimAL5fpBVlsvSn3BWie10O9nIP5VgWtM5m7wXELTbs9kzLgk6MwA0PQez/Y5xqWm+ODt4/A
4rajHwvnrmp/n3V3ad4JI4wEcYOsP3yo1kqv3/k2RSH6jiT/NmJY4+7aS3oFs1Muu+s3JFBSF2fo
smookmllXCVCyi7y1nsBbrWyyq/rVAMZtpGHowAPmkiWwtV3ikDZ45k1QuT0Rwzx/Wqu/GIY4aQX
hPG4lCyN+gkMTLGfToVG4jp8qKpjL0FD01YI9CCQvGYakZ7TZjYZ9ysAzSGIj7FRANYBhaPh61IT
GSaScti2I64BOIagNSJcSvzha8H8eVAlkOCd7xWqM/CrIGpQVIYaEtdo1Vs4W3RY6Jl2cV45SkEd
SUk9+OO4cG110Syl+nwfdvohIyBE5cjjzQIpbUbcyhx5wDnaPAVxNp94EeyU4cVlkU65zjUBi8Mc
OzAYhlgHn7R6wm/4WbN+R3yRdm6N1zmr1+C12wsenMy5RQNwhnC+hRMCtzrLxb/Z971s+mbnjycG
5RLfSZVuROzgyQ+BssRlarZ/OAah6AlBFcSv1ffpBluz/m++NmFQkYfoOTgJX7KUgwRAMoFbsQ4O
fmU6nc0aTFjhRkd+p3IYjihUlXsAypx545Yz91nO/MKF7f1o32U7T5uoRquPLiKq/r0PwFmNkr2A
lzDJhHeCveKgiwjF0FgDFhSJU52sAHbn0v9qe4Jh32yc3X8xb2v9rkf8R61aRn8L/c0LZSgoPNfk
2o/n5GfUZ9gE5uKe44kn7n28XMIappUsDSZZO+hfGf8jlUHX/GW5ryB5Zc9FzQ3WFznnJOKXRkEB
tPbpvWeLEWnCSBpT+3JOnGUmTV6yO7XInEWhBQi++BiHY3Qs4a76xoSZyPe+OtN/CBJgfH1f6mAG
XBcVoTtuAzH4tEUeqOhxxSg/L0qF8cBViWdyJ4z2GJVZXpZ3M1zGD83roTzQZ6bu3THNx4Ecy+dU
77iUs7gC8o7rZIXTmCmcgqlQbicFwYPnWUf9DaAYhaVaYCWPrKl4xiE47PTMzLe3Z5ClovCxSa1C
ZLe+oFLGSSuZrV8T6dpIU6pn9iLUpGoMEGZYIexpKKR1Tj5bG4CjL0SJAD34Tb5KL0uAF4E6VgW3
ssRqCHO+DYnd1Zj0IJEAarWSGHYOxvLwUVnyt1gRs+P3fdrI7E1g9wBVLAez+suixN/ECOgUnW4I
03HlOTBp9DX4vCvnbt1AzaV4yqt9oS3nIAd/rekzRrrDvacwiA2IUGyphPVz4AUVXQ5IePftsUYC
g+vDk/oTzCsZhgy5l6NSi0N+6jrcRO8zUYMWJhoh81e6ATx/NdsJEtRBnnahGpZTlXGjXFNWJR7h
taCb24gSpYd1e9hCYEdhj/CCgsAg20cJNA/RobedZ9oefAQwKb32fQYeHuUdH6pBEpdkTxs8uj9D
5FGNPCo806jIKwUZwjRtaRtscSEE+qas4DjDnUhMwjU0Z+OPgzrfjocp4KTDe6MUitVle2fxcv5v
n2ohRSduh9Yp4KniYqBjBKqQRDg9sYZdCWrUo9OOq43caiSAbJiCh/BM7kUzUCXR1415CJwJvmuq
LxRPZ1vKCGwI9bwlocyT9Sc80/U2GYA2JfjlNaIBVKutX+HSa3VwMBcptNaLymY6/x7LaqfaqjgO
VgqRq09uAi5wjw7myw7W6fPuLnhCMk4XKi1Ugtw4nS000s2n/m1bp+e4UDDL8V78yUEooPnmkO7l
HzGK1/F4kCTbOsntTnX0PA5J/1p6idmPLnsZepfBG9Fw5l2/1A53lfEG0VyPBTby+sG0dRuh2CQr
xe/oWRc6kYC8gGrhPZKAjkltOcR5zIiPhFMnyWY8o4Y0TVIXGEiEIYtwhCYDEJ3VlzIXJpxzETq+
eNar4s3A+eOXojPRm1DBie4RVF9bJIMqTvM5dWw7USn6Bxi1UbKWOd8u0xCPqy9eCosmRZAVeLD+
hHg1M/ov+Q7a3RSAtM6+Z1WHxxSk6MR5hVWlqtjhcjhGOQ8Hvq+gTYAipPaexHLy64Y7rnQsbNdM
vuk+hmAeTdR4o12sPjIzG5XLqe5Ba4Qy4Ckj/o7urif9atUQQWi+h4VX6pZHSY6bRvKpRGQmJopr
IXPopQ3QoAHRFbpqBxsyTl9cQw1jGMkgdp4cpVCPpq3/H21eNXRzhM2fC4+NR0dWVypirqoi9IYL
36NYWufMofQvO8UIk0j0FmmRwzFuUetfnyfBtAd4IwnSpjOTpaUFpvVIgi/ErmLb4/nZYL31CqO4
aQ8YoaW4w9Np4Fv+jKVCYHEiz+rxcWKB17Jsmm3v93VBdgtvRvd64cn508nkWGi9QWuv58BDwUbW
BiPu5n98X6nuUWTqhfCuWPLCuF5WUdW+w4563tLDvbnBYCdJezW7JAtDeDPUN2u4q2EiiIjDhMXa
dAvn6/Tt+ko1kDopI5Dk0/VWWOFqm7qSnBwJWgAj/7eQi1KFy4x/enS60JC/Iz/LT39H9Y01peCQ
gq4yS3vsiU8O1CYsboEuHr/JI2IwKxA694l/qn8jv7KBznGKKgd5D5NG3TIAAINrRCWm2SjKjbr8
t1YqvnUHodx1sCWkhjvqTRv57815QBHtJ7Wl/DehKH0tiXhhlgUclKHSPW9jMBFZfZvKlTyiehBz
GlpCXFG96dFDeSSyL0PQgYtSdB8+3bUcJRoteSbyR2HBOWrZTnASLEkyhuvs3bJS1OXVeBhbwVy6
/VVKHrykhDrxOhN1lvk18yIRIuthJoBF11WY+XRJR2Uqe4cHX9DskUHtKHA2+bHk01k/gL8+ZLXP
vDSe78yaPqEO6EYq689KUdvijfH6bPmtVxjkOmuu60pxnAKqFzGaEcDztbzEVjh8glJzgj7RhNXX
BoR3qPwVNMgf+oq8xySiLzTlXapatOgsR39OPF7RhP2HwbziraP+hOXxdSpAgxT5jEk6DfbB0UCQ
3Zq0VcQzE4z/cvqlKkbh0/1Yw+p2SZ/BsNtXEI+aDa56Oq9UfWvgXRq2vkM4riOBgvcWEXd4dBot
0g9ECpn830cCu9fALtVnjuJeLW6WmZr1UttQaMAXgX0SxURWlRSarK8zvrBzahSWzT5jieQ01RPg
/6d50cYYh7CogFgQbv+PbozqwH2qZWhVeg1JRwwA6R3wMLODBe/ecYheEqSv9bg76bHj5AxFPvo2
fbJfjG7PAq43Zd6xHpLHyeSSfbCVx8UNR2KCpTnuTYRy9sYUaS1EH+7Kl3ztWZU8kwifrLP52HjW
H/FX7Q0xyCQlUyA5HrTM065dUfLHpmLtZPST8q6gDGTf8/5eJuzeyn/HIzi2/9yRHHPR6Ha1J2RI
dF9SRORbdfaz3TWcyIwhLpkopb1hyRLfpctaY3umYzC65W1OiNzUBYU+odI4itMH2Ws+tnr2SzWv
/DYiX/DlvIEPfijkrWZ+eBh8EA+4VPSMOykOjiTtDqSo6YevMmnTIW6Uru8iVdSuiraZaP9LJg2o
Qg/XKaA0fh3OQl5lnmN2xeJ4NITdot++B9ShHhXE+T7t8SL3HEuHMpc6d816/kPI2c6n3vQjeBmE
5X4rENOUbfXInKtOd7TZ02lx4O4y/eqBhnKsDF76O9jS0QON8Jy7hU3O+iWlAYONppVm90cYATA6
jgxLntB+ICUsmx2nVwmSLVgeTidbf0Ve+wMXUMGnrp5/XGod/F8LFYi9kUh0fyd6JLhJKHjrIhq0
Q/NeIJdEq2r2kQuj0Z1f2LF3LzsV4gldxH18YpvAq+6/UluOMhmMrcYWz5kJlr1h/Z495pJ9MkIn
yF2DXfyl+xU01E66g/5oX5PtQeicqSHoZFLS6awFrizmIe2sza4EnTIxm+120DD37js9XvlZCg5y
/ghSpaQ4N/7MPQloHcwxLdbmcGEAJY0JpVReWlRqv4AhGZx1bcV8d53wuQ9LrpEQSgCn1/xeDXQf
lEB6/3qfg1a3EexAy01ghr//66Ky6ZxK6MbkbaBcZZfwxADhdLF/zbBQ7zEQS+YaizY16FTe+5UK
glhox4kMJ9N9rwF2W8n+YpHgD3PDnj6V1jAgXUab5Wjt8dtkwwv4XNnY8A9IwX2X6tT/odSGu8z0
tNhSXu0stJaPyx4+dq+VSzAs/jDKMxyPr2cnbXNkcV9AjT8ljONWcAyGUdnOrLyMoCCjFcfywpyX
493ClLh1MUtLadNMnXF1fx73P8a+FjdDmTg+2Hf24NBuTwaJzmPG/CaCOO6m3AMKGQ6wzjv6BCPZ
3AFzc2XMBn4QEOC+wPZW4wJKS1Gim6WQnJ55Ikn1P4ge+CfsIELi2Lz9h5FSciF9PBaAT1/S9cjB
cIIa+4K4dp1+XoLIdI+pNu+WpT9wxUFoJna9XgIJOeKXtjM/4H9SuTo+/DNKBnLQDR5zX9w2DPMt
3sWznWbZ3vb6NAZPEhpJ7ct8TAcN3T7Z5VlpGTyQXYaYAIkCaFJpCADF2l5I4MB3BVCfJ1Nm1+eI
Ct5QPlCIJaHTx3pGCrtMTvrORO7BnC+pPvwxwvE58sxUr6B+Ew2F5By7kn26viVPMCF6VMEQ9aEH
lJKtg1LtGtzQnlKSzedcJ3t2zM5r/zly6qG9AqYyBBQ9FM1t1ert/yFV56oShpYZjKZvatprSXG0
q9onFp2QXFcJM3x8yWB/Uivqb88sbsFwRgsR/wWO+q9AC1lAcyHm6ZeCmKG/00hB1gFXdRpabSuY
aJO4Zi2hmVLaf6LZ5OMuYBJ6kMp9Y8+huHZocjRFD4RRlkr7MkKBpDuIRyfFVxmvQ7xdq07XJOYn
qpmMN7JaF16Zpmw8VbutkAeFxFzRiWqLvmmeriaK3OlrOgBOQIA/RntrAMlDlThvau8iVzMQJ3Kt
r8lGqTKRDfIccnonyvVSVyFL2VEnU8oR9gld6WzwCiAu3+KsW3105r1BnQJnx4/XHSL+WrKZnQpE
a7FU1lcR3XY/ZJIJ0ZQPsqdJz7ovhA0Rargq/+aWApAZa1BLjMukj8CIbGQh3MgYdg8SlzGp5QpM
/uiVVjJjbcBZAkk02QeKaA2T9lgbMXKPKrWoqmaAu7HSkbQvHICibts9gRY6uSUujjuGyefvb5H4
WeSGQSXHRniLfHsCjm6HzNjf+cA9mmI+W+OmTgQdDsIWfDMILNXhYbn5GM4gwWcdoetXGDuyzfPL
z13we8X4xeUQSaglcCsrgiWYV2Ei1ghK5hE4N1AdL6jYKn+aOG679eImREreLz8C/56YFuY5IXWn
D4uOO4sR/Se1Br0DJC9gkCuG+tOa92LnxrLYbMFdv3WA3bhTSBI0R3gIwLuFwVsrHDL7fEFtjbRH
kMmbjE5q0zujAhpMYMW4GJd8gaZ/hNlFhWXYPvMg5ehG6xFt4ppTmB4lqwY8Fhy+EDyVnq/rDqUV
0dLevMoezr1UsUISlW9G9AMBAWuJ+Gq4m1VcJIgX8lyActZlFFqcGyROMVoVuSYnsH1Z5126f51D
9fGUjeJtEiJcsxlMl+SzxuhAoDTEO3Xz235u8yh+HAbo/KV9etY9ISg3LD9BID6MgOABi5r71sc2
il0VZVw/f3PmB/VXT3I1+fLzsFZAYe0TpsDrYQKhCKzyjEJyYBLXUNzK11XOTuQX+ymBIbQ8jFKi
+jinIZfIm9Fs5hpIh4bOC98xLxRShRrmS3inRkA+9Rih9rCdbdoRrcmwoPpXChbgyQAqG8eV+ZOU
ucaTbeJSLSFEMC+tBca++xyB1m+JGKWGYrX1e5JDtzY8+cwxD34VcjXVcwUCw7nPVlBaEnEBZMEk
AskoNWaptwGMo3YaMZBhOM8pcp2cBtqLD90Ufk3XMKd+nCgRg194pZZVhtNaSfkRXjZtyWGwaaX9
/k/9ADM05JrfB8T7ZlsILPkyrIuW4Hob5zPp4dJmVIp9NnIFhbm3NpkFVoee2ZIinsvrmaoUCWPS
xUX8jQ3IEkLmAHwHLCwPkZKOR3N4OesdbbzSNZmUZlwuaepjtOTrHZkcTPl0SLpNY6C1b2UtEndj
CeWlMsq6ki5nbQk7INQlq+FU5h7whxpxXHiEdXhaJCuy+nkegoI1B6tG8U9yXb1cGjeM7Z8h8/vx
j37fT89UYtlEmZplCi6Dc+XAL4FKqKNYBLfsszn2qDXfWG3Ocb+wTSoJkdp7AXb21Ul0vX39UgAS
ayXfLyZThacHYGd2q0RTYnE+n3IcPm46zVD5Act1vldCNx570OcbbkFDmT/1IF7owiqxXv4FyGBC
LinuEFcGjTI/bHvCu3LPQo8e7BywWzkbu5qfmbwFgHg6QntApAArdM4I8YkNvBmpuyDkNq73OBrz
QsA71/4kiAvDc5yplJMpTPr4XbIKGOa1UjrQjwz3/q2BDlBF+ngEVcBEU00Cu2k5lSYcP66Mcqx1
BlkYu8xYFcAN6lAl6sz3N2yV/sPHfXwDavZz0bCjyiHQJGYldXIOy8zuhzhtLRlojFqwMRX9aBXG
KVgHmA1BiccQnm5WeFUIMqIo++588LaVDGTI2yBz+QcnLadcXpGt3f8XC1rAnl9kti4ZDQD1YHmo
HFXtURAOCMcXzQiASA0y33NE3pYv9RHUnT5CXPm+SUKX1RjqmRgJAVNFsu/8sktEkFq+WBHezbny
ygdFeEJ3pFRtKKVy60JnaIUOQ5l0ZX5H+IYikAazmtU7g621znvWeCdngCWJVRDj4XUJnNweeKax
CeHSURhfIKfQFXogjz/5vK1rEg0v/KOcBZBWLqonznwYE1XrJd9kar4iqVlnV0AYT5gWRzolqzOH
6CT00RGmOinkMZ0I/JdAqmw7msbD7ytkD0eD061jldIWh9aY8jYwZbTUhIOzs+ggFjoYJ1MqJG6H
22Nx2mfhCmbh3jaE7NVXTIBK+mFSZowpPicUw4HNGabr54954/WOe4vNhjY9vlxdKBaeIbHJhE4L
nNjWvMUMQ8MaGT71bNZWkvah450F/1+QV7DF4TOcAMgXLyG/iCViGt42v6dtQJ3zni/kXEdzxAA6
fnaaRfUaSpBWLcaGoq+8aKBIjfC3HKMNtjpGGXiyrTHv0+MuGc6A2zVOtT+Vwka59rygGPJZvHbM
ytxDkqYfcKJVD3QODQMlZzvwDIrVvxYQgPuJxoYB32xNoyeehN74wNxGYMKimLEzsM09qlArbpRz
tR/V9Qb0QhQWIPeLk1qBvMc5zLxcJWDbEdfZ+B4f/VDpAQj6QYVxJd1yGFWvDJOKtrldhJEx5DR/
WKllONYEvYg3angP89LpLUwFcn60y1oE7rpbCJZKFb16Sqg5eIVYjX34Q6Tf6mmvURMXR0oYgy7a
JbDrOZ4VfOTDANc306AuoL82RXYbHSIe0FkeLV0wahoxiH1wNq5lCXWNigQZP4nfdcAwsvAU0T32
yt8uRRqdrzzBb037AHakm+pSK9iXXAsDz/wUiSSttQpDXjn23ChAIXuHkFbAMviqLbsfKeYf7g7K
drLoKp0oKg5BSHgW98c0zgrWhLd99DQ1+Ho5ZOgiGDZR6if9ZR9Jmi8roH6QsVWqjyqQ5qQnnkAQ
igLYv1nVtaFeRk0ay2vHyQI78UrkqReTgorCy8t071ieKjv0+DUIDllwRTPqsJvfBEKYFscTcUfQ
fOfXtSgxNe1TqTj+Dv6JLMAQHwiE2Riczujest39wYRMYMgF2JrCQTLNQ1Mjd4RG8wLKFxM/GfR/
Q1hJ3/wDvseLk4cmiOgMO8yEGg+iHiEBgJA089zlcLHN0waSq16tU0CR3NCzVUpFeWZ5Q9oRGy/5
BwJH1UcfHEm05Tixr81UCRSpbdFo94B7tLI0efRvvRSsiv9UWyxllLTpLkWDDGI7EFQlItduVa4P
8dtYpkq0YcR45yU3ZJpIFi4++86KvStYSUmNtSOHzOmWowhodGXRIDe6UgmIx4DGz0Rb5DRP0lsG
KU14T1K1JDXhQK6ZMGh5Inp6w0X/aYRyGKVEATnSxGnrNJ0Rhekq6K2qbm7c6ThLhf2MxZ3ES1B4
UCDjuKAYobKiuRzcSsF5NAK4FcfsKh038m3RqdM9+nd8xMU/0tEJ/T9OLG0FIMe6mKwZjN8ck5cU
9chw5YHYLv6IzSQHIIwnEAV5rfEZQ0U8NF0bpeD8qc/VanVOij8ki+XRURb+hRDLRKtXl0U5OYem
c5IYkA8c4w+miAtAyTPV+9bPhfiqc+yFTnFGhPKuqX0l8eJBWTHfR9E4FZ087tT4D006G0y/WN6c
C/8s0IAkLrCwzFlclPaF7NjKZoqt3DKYe/d8kBUHecgEpFvSHiwV2vU/Bri7w3AKMEQdppbwYjsY
QIN2jr52TbdpElO28DmJYKJyeGA2HH1grV8sx1mwVS3/wryK8t1+tgmZTvbCivNj5ruHZHumpFns
b5gcxfaBYhahCq0LnSbdCZdhGwqB/OGVlQJEApgAdWTDZlPlODVtFwpWKu6TTVNdchU3MKKZE6kK
f4MNwVRtL+dQOJ3h4+5VVjDWrYrekkyt2cRY8aK63dDeRj5ry2Rzv2YzS8/3SonIjkToCjdVO+nm
kfnh43ATHKJYKr+TVaonk1cMimH+FrZ4F+Xc79cFWEFmj1Ri4GTwsr/YtgGq4va1B3xbtsCDvX6W
kKHyvc4JVBpG6NTPvJWfivJQx3Ym+BYjxWJFfb4qZCjdWReVySruev4wN49T4VC8SO7ByspUSeKP
QYZAD4hhaSGAbtTLf2Ay85pUD0dxa0DJQwTovKUdSYLjY2pOhh/BArBI+206EVKGnLfWY1M+ZwPY
RuJ2b3rMJErFJOjedzRDM2v5BkvbmnjeoXvHUOjd+6xbr0lDaAtgzyMj2IotqM/K9B9A5lPH5dD1
gnezlwftXkqaGvSrbFFhOBfOJsIgaQR51zEmkkY+c24d8WeNJM+s8h02k3UGnua/1cfGx548bJFf
kPqbT2Y2SE+vgz0NQd2t5m4TyRhp3Dh2SSXdcaejD5rjqJ2K20O7Re2w5Z9t3jAm1vPv0PutKpn7
V2solQDAN8ctljH1ejh3Wb9BQiMws2LaIhL0f+zKxshpS7QAKfK2oCuqQTeXx3uis3vsjG9K9w1U
LkTyWwuPmT6AaNIPI6HZtxYhvz6vPnHhia+CgMfXz6kpFxb6rWuNB2PUFKM4D/rUnBCgtOoEzMUy
VHFGNLrMX9ricIDhFGdmYDf84F1uzPFTcwigIGZIN1P6maLUNoQlg4x4puDOcaQF2R5Y6wXxmrqc
lJFIS+XdTNimxy4bGb6ny3qc88PzbSBCVafeOLlhVXkzDWBzHts8S+9qmHjitmqI2ISLspt5RUoB
cJkU5RsqRtsdpu06BV446veSUPRO9xOD7AW0SS5KjPqzp5JMoz/CPGUOsk1npOiHMXBKO93AQ5yc
FR6f5FANf8uVRJXvS+ui9yVN7T123e028BSgaFkkEnZyTKZON4/YxJ69+tRx1jH7+3m2H5pSFDp/
pNuxjvmJzS6QYFFqpEVZQ691iaBHVJmdOqAeFuaLfm5Dqol0p6i5FG6W97nMhqx47wSf7AwOBL5s
DcKMygCvCqvSefq8kI42A7ud9+mCcva+PCWYuzV7dxiv1rBMo6jGWIZRTFIAim9/kZA2I/jD6yml
aN0T54LLQgkdyvhrVxGzoB/C1nx7QreEJik5HwEVNRXJ2PqJA5VsFJL/uCqJKbvYf1A9gcE4iE5d
XbwLufLDoZByMfALDgP9JLuPp2RRCckkjH9jVMk6M6AYt3FuuGT2MCl9Ypm4sktR00vA3tPENou0
Fjs7TklK+OXlv3dY3n0b1QXWGjn88uBme0hSJaoD0bEgf/Waa6N3vw8A6b4HEOh5JHAv3vubdWt0
h6icGKYtPLe89QlNfCzhCJHtYg8ev3IuyTi5jId286XNjzsD2jQGjeDX/bb6vs3ycvlx9HW0qB+O
WjogVjIvBt5xqMSq/xqIQEY3J3UsxcMVbFH+NSXdHLzpFM2lCpkyTKTLwsoiVtz6yad7gq1/fyfn
XOPghusWVTPSwiJMKWElPkISBdNCKFdyLPF1AxbiB//pbEroc6b9Ega6Ia1+nCBTdtNLG3AFVjas
ZLMlUJMYWe8yuHvBKHvHvneWNFCSOz2ONQlJbx/4trbkHvPTkPLtyNbRk/ZQhC4TBvTqLu7eRxPi
tu9IHNGM4ZIjcv4zUOIHmRTVPBxmEEua2FVIhPfp3aPEQrHBIIXFbouFzsF8vcQUDLdmcDicszSU
G6K+wkfciYI1PEfNCV6P9YnWLmamwuh5M5seIHbFBayqX8mrts8Qr6mgCgq1ZrLNEGesU79W7uof
rZF580u1H+6RPcZotWqwKbX+w7Xy2vkGXM2pItXgvScsAZnE398CQm7jwR8+124nzrsYn+yxO/DM
XiTrma8/54ZPHp1yHt9gDq8dFTQSJDj36bYXXUxS7aFwRd1fubN1Xiut0r5yTYwtKHWbv+MXweH0
vLFegguoT57xH3zjohXL+0WVD5YWUOrLdXpub2/x20MqSEPIzj9OaJYxQnDFnFSpA/Cce6XfpLrF
ExIRiYb5ZaPpep8O4KttLzAR3aNdiIGT3UZGDUuur/0NqBA9YmIHOKrvRaxxVeICzns8skGYLUXG
/aUQIaEuyt44R0tFYkTx1jkM3fERWQqveFq0l1C+Ia9mwLN1XKXMPOmNOOARbb6ine0fynan8CDf
Gtg6SDDNSeRx8KDkcliXQbkPuvA95ew3+UfJyz1YxOTJ9kuO0iFx1+3qFVbzIbZnQ13ISc4dM80k
lddcwwohmipnTf0tnpZcz4lVybtobxLpC+POOHB9eb/JHM8hNxp5sqV5sfuFjjqKM0WR+RTeTXnf
3nkw1ND+45tC5Sd9ps5vqtAQYWJmKrJdenTlUiUU5qi4i2b5O/eGBppoxBSQgHKaWr2IFSR/sm9U
jhJVkiWJhIa6LHJn4cOZSm/lvMOh+bt7yBPN2N6TtLIedzzUQqrzhK7RRofGXueru8QZmr/HFKQo
MIi8tK9g3K42yenLRYUvChDGqbpGQOmaltNFIpL8cOEM+b/iVryRiCETC63qOzkz2+Lth/OKScdM
MC+bKRJnEZ/zjnGFfMtLVDHiB+grMP3FrwwadnIkSafReoYPkcYH4AazZWEsfMqYo3X5GL02/3iO
wvMunzDo7BgwkXqzPzEhumZ1WV6JGoAj+ceqqIoGi4Izi174YhS4E51AmfRRYbykn9gKbbBHddHj
SZNyvd4Y2bJs45h7V4gv42C3DTtzK5aQTjoSTVBRmcL1nGaALlt94jIF3HjYhLvuTZ1CLjn28ylP
zuoungUX5tq3DBym6RHvxYNBfjrGwf+Epbf1VM9pOEiSXAZX0Pf1TURLY6AAQpIE+6SbzF1Riiqi
0UtK6hMj9FQoxp2W8PsnSbFWJIg5aGi2os7YqaeONonAwPf2yTHGsobBitVW7M9uc0eDiJL5yktG
qpo/0G5pcDRi5v2QJHtprOLizF9a7ylpquHsk/1KvAEs8UWVwgYQzhG/eW8Lavs+udiZvroe66Vc
76FdqlceCub0i7ue4ZIi01WUgTW7HZQC73+ou23/Mq4m1oiE+fXJj3xR/+Rx4I7tMw1YLyACqg7U
L/2f2vCrboFM7UmYWgKu1tshIcmeLAtw8Vdni46otRtH8mmepgzsIB885fX4PkFnxzIzz+jaX27a
mGT3I70KpEdCM2QYC8KMhj+PKKpFUgGSSNXkMUYMLDq7zVsXEwlogGUkXv9Kydcgv6iNPIFgsUb4
OAQgSHBXQ5NIw8e1juHqrYe8LWFZEnTJGCfTURta16ld1XT/5Hlnw0ix3pnS4t7eW/kIprKkMWnq
atUC82C+MH1G2g7+xIaWKzYUqHMJKfnTo1PPWSeo5mpOK5VaCAvU+pLIaULiFcv5avgySUqLEY+3
/LcR2ryXSkAjMOrH7aXgytzkj1cgFJBgTSaxIjp1fS6Z1KQvIOk5sZKV/LzLrcYA4s2UF14+jyV4
ISQfpM6+buYLhzV9/RJuCcNoo4HJDoxx4TlmTXdDHf0Vabt8iASqkXdvfYlpT1XfR8Zaticd4kDZ
80b3kJAJ9TA/aSEfHc6L5uH9plfzMNh/ETJJPtLFc3nQ5XWNExXnQDBi8r2XR5NHd76i1Hj6Snlb
q28co+5OXly63KayitAGpCMwyb850ucX+heeuMc2o9SYPyBRgPNF6uEPtardnjCULYhy8k2qcdyI
Jhb+MJVUG5tyuLTP8PlpF7yCgFNOWOKjXvSzX7BOlqNIuBiqGwKloTBvd1vZehL9yC7fpC/K0AD0
K9tP5NlfRky32ayCkxjNmfd/3VTjOkBuS7Bdcz1gSAXDQGi5IwjhSg9/W+V0Fkwnxfnzx9v9402i
9bu5oIPTMaf1If2NVBbHVjiQGPEmeaPtRcrT2aqhjWJeRV7J3Y4BNlRvmIKGgZj1XUCiOjnBYFAu
diH7/FBVtxtL1MG/243ZPPwpiJSEP+UwgGAts3PxvQ0NoeWOvX34tnR0We3kpYtHb+B5zUwcrkdj
OMlgzqRV5b5z+setuIzJMl1w9Y4rFVBOsXl+UuIKBF8hrG8pjumhfvGDtke7s2yNgnn+DIeljzxY
oRocjFNjIVrDaXNm0Y3FhCCfaUXXF9boVH5Z5dIrsCe5K3/EcM4qtukVJ3JaP4ZcSR5+ru9n90AZ
vxG+A0PH0j4e61A5qcb2e2omCB2Q865oDLBGbmiesCos66KaP+FwBJjB0oXQSiWO5KAWdv0wbQjh
QaiMFxunM5z9zfjs78andBh/tewI78nqcLN6DGD1uaj+Mbd+VSJ4msW/MTHJc7YWoIbPGNHkxMhz
8VV8oDW3nwQUNqMvxrZNKp5G0BfnqD+MOsrxTiRKQXf9DYTyWZosvvZKzUduubTe7cay6QSSA29h
Xn+QrszH5E3Z5MJjcdShg37qaJZyyqbTnUP4bl2Y4cVtAwrrMw+221pB7UFRzT/b65OR11HOPTAH
sDpo3VsMos8GCeLffhwLRThBZUc9fNXRlFdyfaLurPX7KzkFkqpxkyXHaYWX9CfhjqGgWsuvXSXm
I93NK64vJWrZiJNUJIjfTXmd4h3VpQv7TI08DM9AdoZmJ96LPfmqddu2daH9hbJ+qjdlOsLYmEEX
xYVrdbIriD9+D5Cz2ubNuo0smKBA4hDP2xVTwiGwMtLrYyS6EivXBHJPq5UkeJPzS9Ll3rK+FXJA
vJnonhowOZyByjUjKb50xvs7JtAvBifaK47FemmF1bYSarQ4OSKO6CdmngQfZT56dzD1qfcvXDgf
g255bMs6dWIf52nE+z5Zjk8zbE1XKnIjpclh+koFI68iyfjsWs+CbY6of6/9wqJBKWxC35ibR4OI
zPTT760fo0MFm7zQ8YsxHVy3iWCQrRzD5FJgWIoz0T9SCuJzxtTB5jbv0HnQn/sNa5WyGPtKeAJh
mzcbmVUK3v4uimcQjUmdt6cjLY4S+QhlHBTRt8SN72+jGZS56+LujPRWeqdiERqVjUoc9sOFbi7G
jlv2sF6ZR5kIx20glHsNDM8U0RrhqNYdQ4xm/TF/zCL7ULKd8kLBA37QqwKazqaBWFOCEulVAUQ5
eOCgeYkOD763eGMrev+u6bZTpLMfsCgwaM0minSk82XbXUdvtFPLa/rODwB7QDhy3Y9kB1L5xWUE
6sAdkQcAaOt+JLPnZ7tRLkiCVw+TDTAp+0Jp3o1rNf0i1O7kz5af3aCD8JpVoHZEKIkmdTEmK7W1
yDgYAH+drIHH7x0iTVncfY/xEF0N2KobIqS6pDHeBFdQIkiADFaMfIcV1Zn3EHg/csaT6goy80JA
XHNAIaOaixpv+SrYHUAZdHLdh3GIara8ICx98sgXzCQc51xRqukJo9nVQrwGiJap+J5Q+jEYKDNR
tu1tM1ikTpj42+OM3d1+/V0yYDVzAcJlxETkJ6r4/Nvc98qY4qzfbpBecFIQspm2Y66BTT2gRall
AVRS1cC/Rl6b/BkPGZVbx8f2ON2HJAlDio2LTY5f5yoh3PUxbLcsmOaLs1a9KMjzi7Z0E5Wt4QEW
3Lw19VKG9mzVSjXoMZpy2f9gzfnzCO7Qv9F7sl3bqyi7RzLIahoak3KXGGQ1/PTXas2QO2vLtMd3
2yWNeHnfuDlsw966uWpqIbDdHtOVIY2wv21lwBET44zsNc0IToLaBuBqKye5AHbAWO2E5oY0UhEf
ZXsG3dMqFdgNsaYowzQO7M6vfxV2exVWy4HzIdxvZ35+/eHJu/SfnFdiE+jSVWm1c5fl1UA7rNRo
hKX3lgwMFj7KH3o18Alwt0MSc8IV+KdPN5w4WOQgNlTTTWHAI6zo+Lr2V+n7VZWpevCVxPB63xRu
GpY1RZRa+qCHQqElbsPlz0NZ5XZhsxc7DQWru2dBu7/nNkmOSLoYfEi+GuOCXW+1n6Y+x8xjqYpn
9qtAeGigthl1mJocCLkqMMscqrYX3Q78hNlCODCoipc45mlAHHSP/59BJ5ulu0yubhBtAyXEdLUG
aL1UuBA9mI3Oim2bqi5uqPd+oxcxa+SUdR9SwjjJccsnFvzWjXNvyLqWQ54Mk1kGU2PzbzXgcwtz
8gdhmqz1jvCicASbha8zDZVqlAXsPMeR2M/cjMwdPtQrZix3202ynYDP4l7bDUt0dYXANEPjB8j1
wlT0XJsrUgofkeyB7an+YGHwsvbORE1DWUYoexkwI5kG8xx7PNZq+0OEAd0OyfGl/0Ja7BfhLYEm
HVsZ4keZQqf4OAtt1kYJbxZz2rxpuygv2f54jKiQEjhRMKcJtAnvqI5s0s+dJh6LdDPyJuCcAIfW
/RfN7Go4JDr6ysGYK1b7zK+BLJ2/jCfjSaQbZ0theRFl91SpZrdbomqsMcTsDvlvoe6jIYOTsbCs
+7pKbmxI/i8euh6Oi5sslw5aWz89W8YnwhJTTgmBwKwEsBSpvCIEwVL1CYHq/EPupsHz51Lo4XlL
CKevRWlNmkHCwHc3bGCDGkilruPY2LXkgKe7p5yHXBS/8Te1oGzdllS2ms9u2qGcVr9juLvuQe2Q
SXI+JMKUWfvXT0TBjamiygpQR8LQtBnqCz1VdrDTerCLP2NeRnNJ//KhtiWYYL3WbF3MsPuLOHfK
dZLplpMsrxuT/ie4aJEwnYS/DPlZ6qOTnwmurieaKjqwjR7x1efsCJUkegu35MOsx6Pek4oEC1ph
Cg2D9vKjWO+6NExr3jvwKpLOI0DljwODApcEM9ViAtRO2iZkH6JsUEPyBCWiQxqq7dq/8LEIFNnO
98SIO6F82PUZJ4Yl2TDoWFxZ66iMfHK6cvCSh+0jZ3xgiz7J2URYytTs7vgOnqpj7KRHMK5ryakN
O3BBNAa1GjyF95Gtq6l8XEbyQ9RPjbg9oREJS+MydNbmpCBpSTnZzikyGEO4B6w9lKRL6XSnoLsQ
95TRJeQ4ddm72J1p38ZekAybM8aaTZtcyq8SqP1pidGA12iKi/qEzcOfnKIKdEDrocf4gwDSWDMd
AYdGkUvNr8ijMK/JpvmcFDzgcS7DZCOy8j/4VpiIdlX2XkzF+S9d+LW4N9OazmHfh6QG1T8rAjBR
BUd8ud4cVaPvWs4it2u17nS8HMcwSKjNBMtAovfkCSkfJdJ7TZ8bugOhQd7nuU/Us1V9xoLBCryK
WU3Cl+qpR1XIa4wlehhWJ3inHof4SS6OURtqYpOipufOElSUm4K6NKWDYK7AYn9wPFyH9QlLztdf
CcrLh/a22FYJ/boiXwm0Xg4limaEac2F7P2EGzwOoFynEOfAgzI/lzo+E8Hejvy1FDBdMcd7iU+w
J4oXZ+D+5b4WFbrOUgXc7iaCnhKTmKkiF4AOcLJ2IvYRSBHXsYOcze2d6h/hHxZPDomoVhxSfdwl
x913Su32aiHqv0pf0aYK7j2Qhn5QbmLe/qqHTOqy+PyK/OS/8EUtO8iAP+wP6KG/3b3K77a/gq4i
IEwNDlpgMAv7O5bcNCKvYJQUlFXsH0NvgSezINkUmGvDUj8eaHPx/vqpDBUyu6hbl7xtFCGBowz5
fIpP7tPN6MdE5/XZqZR3Dslf+fUsak06EUH+8MBGt2R+9Wgl6g0P/6GhwEWykLAN3Z+I2pPSt2pW
GH6x4e67PoAGjbxuVCSWS0vsLNXH+INZwEfTmhIPB14Ul6bXTsTh5+FeJwhnZSlXnC9IPT+/K/A5
7QFXOW1EtLpUD5UM0ERRbY+mZJSQFpBFiROa7helT8AeKp5QJQbb4vuNJhCkFyQDIITLUJQl2Nz8
kPll4geT7AYh3TFvUHxNQ0Uubn+QVGH3rSosmN0W5t8m0vvw6ANxMHp6V7pM6zi9D3JUbMXgcBK9
vVTtq5Qm3eVKBEq5/kUDWBErhXykEcv8ii1lOb1tmdUG/uo+XNDzS8oKJ14tX39uwXhvBgVDBx7t
lPm77QquyjGozHfRCsrTJ/T5Xs/MVcK3itG9BfQF0VOheKnBBmrTqec6vatPuZZk7/TDC6MYNMvC
scVHdCkYS9Yvr6YLjQP1P2+oLzC2uxV2Ho0A0w/jFpf4l8JvGkUu35EJ8UfU07yfo+JhomC44UuT
dcWAcFswXAR25QRK3E7AKmXKeNH0QjFWhJTYCzGogXA0Op4YEAmuaHkavnIqys2oLTfrs+F32VPp
GMQ/K1qOEfHgOAi6CTVQJCrFz6TNVyn+Qz6+5scngODiGGJPHvJc+/5XrZ8mOX1gXixu4iqZOi7b
NSnkLhP4m+iwr/MalRqYwHb8+tDjNq+VeZmIvTTfZp/BPbMjUzDzvczwhnKYJrDKWdMQ8ijoxdGU
BlJRZwbZGX92wxkkDstiOaezctTQBT/0LKiSHnLV2bIeMnwdJAGbFlD3rdoJ8yjIyY9hhH+NPgr5
7bDW5sW4dn76zbbzthMYELuf2w68LR3bULbMmrzna+omLNUVUcx+PzRX+Pt3yxqA5QsAi+KwFFwR
TQgZuLlIqtKo9NsGT3aTAPLiopTP+Kuaj/oBjiu3wGkMhnriadee7jtfESrwcdWbhlj38zApiZyM
PlOqwjQts/P3hhrRvbC2uBeUvZx5eUQwT6t/lGCxFJ7xVcQhA00jkRv63pJDLL3hCWRLqxDz0Cpm
jDD3l5/u4N3gKwTuSWCu6XVKs7b+lDk72F69Gi5QyJ7Hdx/zPqoeuLwWUdcr25jRulQMk26BdPb0
CpgEGwWPleHb4JY0Zf1igjfc9+VAKzVKrFWErP68qAT403/k8AfCynrbYNMiabM9XeoD1YKLYmb2
xgQYHyJV4gyJK3x7o8fvuclDXC1IbiQqY4jWpPjtRdEl8B2Bvzh5jBeAHI/IpawiBaUYiqK3hJB6
ZEPVkQ6w/e4rKsqiZw3LxcJYwBxmY6GPXAPer9XAL9Cmc2qgGDWqj1wA7zCUDwITOHUV6cJ0LMiw
Foelk3ZmziB50T2P8bIyI59zFjcHtM87wcX6f2iAL3b9hLSF7OP+JQOOML1qOBIFkE665vP4mkst
WbXTQkpgg7Ssrco59gOARe9TYH2LuV8+JEsNTblXng7s7PHmRS1bdRRTZZ63zDGnRXIHTOhWLjHe
Uqgtyu5I3xIiTGIaFjvk+ux2luz+Lrvpw8aXN2cUbiZnqF+d+85yjD7VCMVOdiHHT7DC8KDikiMd
f6ttg/9Dp1M5XAKLx3V1MCpRd0vD2Xi5jSCLl9M3UTgfXseJOybsbwGLD5FykZWFi34RCUQfAms4
CdkQ+rTM7gVKfNurP6OfCE2bVu5OP3eiAc8RJtCCsEcZbsjft1yA9uTgUus5DZjQAIzAjpyk0mk/
XQczi4sQAzssF55W4LjBH2f8RYvsersUcZIbmVImmBUx/gS/MThi6AAzDBaTdBeCZ6rMmC6lzxam
vQL2W30bwZ2A0Q+oxhVOJiE/xUftrP+kroDZjMxu2vGmrVyR/kwOIT9Ix8cfiirQUW1hEwPekudn
fJVPLsf/xOAfYbwaMyLyXB7rq0R7bLsLzRKZ7Rc0SYUYbsyF0Zw7fYx3Rxu6dOST54Hhoegi0vP1
5y00E+mzEthIF3O2/eiDxSUI77c9h91LdWQhnpPZgZNKZ/NsUJn4xXlPLkFWZ8/OkJCgfiRJPQ93
7D5fp6C/xOFQlhjnmdm8bgb1ebwppUZE7/4ZM8/OolYr3w2JVpHvbI8oZ4OjchlUEpQkXtYNGRm0
JoLnlBFMPStGiKvSVffG6XSBYiyOSHMFFKp9sXQ1pT3R02PPf6NiEHS0F5woWbfOBadN5ybTKPFE
MsT6gDrDzTFjK8im0Kk9VQ4vwAl1v8rbIGa+uY1JiwX2u4cnHxy/z2sCYgOGbX/02Pfq6nueDHig
HtXYnrOch03Z4kXGBGeNresqfLCOsiqegm0wR2uwPRdWVI2Ifv6aYWwxcMe0mFk2FU/Mmy8C35lR
wYh/SdU3lh+UfjMU81F6LRYQb2E4K8xW/BePTkWTLmdmQjwxpotrxwnXhe+Nhmy2raw16nIsrlBZ
FmPzJEXA9KnprKPESxmAoSUeFjYB7IvpB6VS5eEkaJXAUJlsw0p1BK68vDskQbc+kcAS9S68SUnW
rAQHla2RMVjltkS/sToK9PpEqWAXBSoW6HVzG9nD1psHAeM0VKAuf37ZgNlzVuron1KFCG7Z4Ndw
y+ZsPskNkfpccDVubrd7hdt5mj03asbZfRfuHO7yY4nb3ZsMmFNTfvmPfrwwoYKCrRLpuXE1aNsh
IX7j2FuuP+REnjiIk0DAX1M3qeGruO0TCaRcY+CWtgC9Kpgh6H4tilYnpBXKbbAzjsEVQxDRIeMc
QUWBaspoztvaFKKpgDuuPNZjuPvWv5TBxA2TkX+rg+CQq3ElCxF6OQqh8lUlnS/p25F86Myd5Fxm
AFj1v7r3gR2niiErNJTRXqpEDIHjQ4I+NcBqhm1KscHhEHo46LdECZeJiz8aLFSKa5hO9k8zaB/N
xKY+mngVTJb4gdhcG+hXWzlKdhfSANJbpAqPM0CrTUmYBlTWINUIAP+NQ0xEC9UAFpP8iljymnTN
wPxq1ikAxuEw6Ae84p4E//v1dOzPP/LxxJuYl+AWZ1QXOWEaTwiGkTFCbQJ+NEysQTSamBWDcjQd
l22qUz5ivTi4czU8i2UEC9pPXvWS1qGVFlJCILZfnBrlnFAMf+wOIk7luSwUFDXmv09QbxY+rvWq
l2Jm84OBqKAkrtuhIzd2D1/hMMc5xLJ8MQz717yqe9vsfEpbXC48qPNwrhcvouG5k5B4v76H2Ft4
v7Rfzq4bZLDKG4FILadlkHD+V29Mmw/uD1hhB5ZMhf+hjk/sHqylOSqFQIvMRn+9d0A4sMDH/FfR
m3gVujNKjNQjya2pdxxP8BJ3g8kl3z0fHNwVxQSIqIW/IsMkDROJK4Z14ws9NDXVBN9oF2Kg6r8K
omPtouaB3ffVxcBjq8aVnu488puST+L2yu3fZzUuI9lqQi+6YBR86IdWRvTTqbn6lNiHcrl+7pN4
ZorWEQ4EF1Y4DutQBSTb0GEXSHZUqyTobbK50wGsyrmYd6UYg7AsPGqhe6Rwt4uLFYWvWCESg5pg
4sLSfa8b9pR6rQrbqzenXN36YDY59envqVLSkHpI1dAN+khj5H9D9Lyy6Tw6aSgtclkyr2Cmz1VX
IaIj1tJWI8/tqJkO5v+6aTRY14by8Xym1YGOlrUDRuGe0bri+Zyvx1sFEGwAUsnhdqiOIw+XiWTE
wYvpvCT5AFHOxRvuPPCN3yp+Siu7Nu+ZsctbMzqPDDutctR5OScCczty+tl9lPK1GmsWcJiRerKu
VGOAiFmpQ2EBDh45x2n0x17W+fSTG/WnJMDvDOjICBi2T2zgS3hNQiATsR1HArVfSCTWnmXxLNVs
5bqpcV2igS/+nGvMt7kt0cg+v6hoEzYl3YPY8vk08+p3ORIgKGJrfpRm9zhQqdwjm7eXZcE2YUW2
+msN+IVlvG2jJEI3wR5SsOOXi/L44q9qyXm3Gf0REcpTyrGOvV/1UKFIDnC9c1VW/PzjomMh++9B
+vAFDzkAN5HL0uE33beX2DGrc9yCtLG43qyWTjEuoEKhEeQ96KUMK29tkovUyHnaNuOlV26oKiRD
LpPwwTgo/4Y+Fcwx2DSyKrghI+BoMA2LGR8YatKViih81F2XrmQUO4JdWIGLsZpiZXoa8gcu0lfz
sgT0ZYCxvfZ2PzT2ZuHxa0qlNdvi5wiscsA5Jlltkbn8aBnzfIXB3tbSwk/ShDQPhdB1lBoWdMZ6
HBEzYsKkaHenVn3k97nz4d+VUwo+hx8ckUF6fO3ZV+7b3i43gP8aa6WceiAyr0xgyIf2PyjTcLhr
OxDGqt/AtyAppYf+eUifPTCujeKmXSD23G1I50pr2Akt50gNvUGDtzitOqkXSB8TdHtRyBM3uAh3
abyhs3W5PFGL1f9qEeSCBTrYjy7SzcFlUvvjvxOzq/o+ZJVAYr5A5i3gEqu5AZMVWjwmOP1OUP0O
fnv4CLboe+/Dekv8oxd3Xsfh2oUXrqI20xXgRY8NLFhe1mIbvUPDOdl3d6AuWsIKjjHLo5Ea/dJa
j/FZd/O8IWkuOESOB+XwmD3a+sRrvr3+634kZBgSsAbrKD3KV/nEb9lz/F1dVrpqbZ873qBv9dJl
At4VA3kh+TOKpsW/BIvffjbhYXp28nYRIcwH08P3deTYDS58u1302JwDpAPAnC14R8OqvOl9o/mX
34rDlVFdbBYBO9kfpWodp4uzI4Ahr0Vkei/OLYMyWYL+dklLYic5GVqEV+7Z0K9vw+GM0oyYUwC6
mkDUVsIkT7SBGH/QUpE+a3XzdAo2y/Uc4QjXCTDJeLSokYCclv9RWfTz4PHBiIPpMLMfZjhN8vQl
9XZLBMcLCNmYh1hDSlp3b9AxwMlWEHo7dvRUBl2RBiskzEQsE+AuJ8uh6W3YBli4qWS4i15ZEO0m
tftW11/hhrpyqJNoBZBGd6BIyeH8o6X9wcgQexT3uwWGjCFhLIloZehlF2Z3RxDnNeWazZOQntG8
l7/QboBqymRLgiO8Y3fI66WETX9sCf/PR7wKtzo0V6uG43HXVm5ka/Hs8RXgIFUyYWpASP3e4f72
ovEEt11K9OfGF8HqjVyqa1AL2ptYDHWaf5OuimuJeNQe/eXLYLI0jpJrXbhBdSGmubxQqbENurju
+4g6gqozmm2dmgsQRTi6GDoS08epOsxGXYjjpz3YbGcng/8OyKzBXx62bCsxlMyHtiho4+fs/5wS
wvK97fr+PaFkTknXCbHlD8Nr603HIe02dNhQA565RkFmyMPFpD9IjNUfJrazANu5fUhOTtyRzgmB
mewzrBKwyFOJk5atQVi814+3pf+Dkv4xqB3nbaqvImUUlac0MZRBbVpWyppKqIqVfHz2EArREtiu
+McQHEw5gRIgoNeYxDTlA3iW1P3Se+MiTHD/vjfc2qE13HcQkRMso92RPd4UCcx9eV6oEevKtYSF
oNOfbfv+0fj/kQz4G7dD7jd7pep6AQv6Clk7ZtAxkw3fG2xMVSA29OS6hJgROiSIKNHpdbVWxKkX
tRO5nVGGxxGvIVlJJEzTEzD+JTO9jevJPjy/MEDMEliB2NLqMfWyx/EfLExMd8/kEUZEd+JPlGs/
ViaTeBAz64D1g7oKMYDliPsCqwIDsQm+rN6ULcB4HFu9LmEth1C77Y7thXIHPON46HGoBLN2awAT
OzVe5nH3VIseUvd44ARtMDmPEP79IZ/b00YToU2QFJaXLWow5xihcdE8criAAB5riwR8l7JPfqYn
TsZF+THzNCQtijXhgT7y8KDiknT5dCbMD6jgDyKlXn38d44ksZUQGTAqJ9jWkTbhsMPUXY2xEnS3
crJ6N+1OPUtWVpgvP80RIDXFCdIeidisOEpPGUSHU1VTcZMkxsbS++hZua24DoymrQNTAPe3BWrL
gY64FV2muxJT07/V822JDHK58GH73lPGqgteH+08ZzuJHeaq6lzvAM4vuvOn+rWcFAuY8Q2qAi5G
GM3XIIf1L9ug+XcRs0ZJNuy8jsAg5LzJbqnKMtv7ZIbZVabIQ5789iqjReD9rpj0LTflnokcpX5L
IsaGBag2fSyRnDosuVUmbTYpQ0nW5mkOpzBaaGLyyMuqjN5CptwSPBB6re9I+J3rkM4dd7t5od3I
NjOTt5h5WD7oMWSzDDTCvIEp9dXIFmpQSyTG7y2AOVNI3JWzc96+czBxuYJimOunfiya58Kn601u
rWMj1x7e/NrUcilvAIoKszl9GyZv7nG+134aV7sO9DpnufUf7fbdn3OrOtQ3slWuOEFZTIAwcpTN
uttD6OnHRNGKkhDOzzhKVTO8orc1J/Ny2+GQKu6rk+zhz3zwfFNc6BE5Xum8cbbXhvtuPG4Ig3e0
DJ1JyiTzHaGoH1AnL2fJ8xTFb1J+gzjAFreeSqiIoelupQ0m1Hk5DBEQnGXDDiUk4SNBJ2rs8v4X
UHifyaXHmjfVB7BXSXOKo+TeXhej0ptIGgGnEpWxdiib5aR7owxfqsYrPNlx1+1NLpaeNYO760JA
XDUJPY5utu2IVhhSnFKYa7+YIlQ5WpfNmeqZyhVnNspCdKMjV44aaQ7OYa75pj97JT+mIRM5fPsl
aCqYGBAetktp9SHgb5xwQYEapQ3cw+stfchhAn1eyDD+Yxx1Cf6ciAYqwrTa/XfiHGf2kmSF18nQ
7SPK8mFjiaZJvS/huxkDaXK8YyenSSr6cR/I5uEc3N2qoX5djlXquEm/mY754eFONcdON5Tb9P2a
33kyWP5yeLCQYYIjKN4ukO+TodXBrJNz6mvu4UEOvduJG8kVTvXSSLUbffECoTTpT1e69i/UHoNR
Xbh2njGDfpiXJTBKSJNYp6zvt3TFDH0E7E6lOYZncaBo2YatCKHemqczw6Xw5MGT73M14rd+fUZ+
qqme8Q2KxEYIDhNioIfyLCQKwt9J6CqhH7Xq38+IPmnhSxWijbg5WtU+pEaCMs2VBfxZVc3ogBY/
PAdyI1EJPmjshVZgjXd8MG+MFmHBCccTmFcx0BR2FD/ATxq9hkqX2iFxjwEbf0H0IHSSqwX8LHG4
fNF1rIwy44CdcWuUot4oJgTwT7RT0uZoE38Diyt522jY6fYWCi90WvcKfEG9UxWdEARpeYMTzijP
Ye/XcVOz+YIDrtGxU78vtpG8Iiryot71zNaQwDdV6EqFVwb1rgacjVj/tnudhYf/Ru/t0eUuQ9Pl
q0R0kZ8Pxmxk4rR0rXDVKM03M97VXnLxS2Sm41uuGnYHeuAxru1tXNDIQbStcWtNOAQCqsIICaYb
TIDEnRWAKcBiLfJvE0TXkNfAgWCv14B0Y5h09dyj4ihW0O4qkrAZjdbKSx1jSrcRQxl7Q6FKYG7j
muNCzjtJtLxaFpEzjVZd/k5dIY3ygevyA8bQLA1528QJIGoq04v46IkL9usw3aZJej9ug1lVHXKM
eoKNqnGCgZ4dOfl7lor01RjjWecPKu1DLVKd2Af7jFSE8x0P91KjyI7Kulc+5Y46352d35IJ1MJ+
e7zVlgIjEH+cSra24upvJx8yYGxUIVYoghPX4ZhAbDmBoPvePhChPD5+lenxcu0+EJQmZJK2f0od
1WFo4E1aim4mdBWRbg2/Am1OK9Uap9Z2OdYdzXPpM1+7y15jrjBNG+yOznY/0PaalBdVvs4qEKZw
gop8sTs3WiWNnYCS1hqaWlR6Znx4QQxTFNTyOFgSmyyJ97kwMr9TSj5d8ik76mqILqFnC0VtJASP
y3Yq8jAveYncfN1moPcGzdMFn02qn7Nb2xg4X+8pd6KqD/Gt91yAArJzbG8zFEl21ckd67YwE6Hn
vr3pf+oz32Z/Ta3c3H8H+tAhXqXjWoqq6kZHXrbC9zedTbW3E7FkXvmySxuPAJlperwrQInEYw7r
vP5HPOlbJpPrHlgX2zH/W8v1DSy36PBGy+s07yDtdpLacjMB6WU3xbsfnd3eGle11HWDQUjkjT2y
JFKa+P0WwzuuXXsRQtL7YyyYvRbR0umfDkEYbXY3xKn7Wbpzl3LZLiYuD2S26ldF5AykVfzUDM29
WDT73CJSc3x8Zj+m1JEf3cFxekOF9VmNwlqU8S1yieDirOOI0mYGSEM/oW3ooBDZ1ZuMAEbtQanV
FdFL8oSvQ5rNeg3sdyW0xWLFRc+NE/PfLn2UmDbT+kk6gwukOTTBKck0wKrAmqOeQjMyiw7zV5tJ
RTMElK8IRlwqVez04EyQWmWSnBzYBuw+afMIaU8m8+O2wwV2p8dKsUQNskMITXuf1LerQh/5Nnc0
N67jPudkqL386GDEUSBJ0dj+a5VkOpBBS53+Qm+ZvLG11VCBOGq1Qlt3W0Gd7MDACcffceUzcJT6
K4B2pAB6MV+SqKPCNfjxphlFht38F6NWQ+RJRjSTwVtXYfXdhjkU+X3hOrK8Ly+dao9dXpjy+koc
aeaQokYsUxWpMsnIhNNcK0mvcdYKWBYaDbPseveplCHB811fVQRVTnJrVfgExo/zGRn4xABpUaDV
zxw3o9O8yDrQzC2v/4NarikxJp6XnJWm5WX7G88fsLBhUKNU/JabmhpETB7fIj5ZdNccf43Q9B0l
eiD4YbkfLSq904FhL683kGhFq96FlQxFU7gpiFAjuhS0GNqDi5N1IolSnG4S5uZPgwsH4SWQe3/J
heVIwcqy52qAhJ577jjVLOZVXQAlI65b6DAFPpVf9dn7Dz1QFLU+kN5Ke/1QZ5hzaNU2crKBBm3x
6A44CBvrKuP1hcpuay8h1uS0mYM71NlGc+km6K4xHbLZt6BEbgh5DU0/r3KIaoml1Y6zE7nmN7PA
JTqzJ/ggOjGT3mafXAhfj54fVK+AewooOuCX6HPdIcR4g4ObG/Ywhu9UYxHAst1D8PpnDm/bHwLv
yC7z9tM1g1uSvZBqv7hMdayTW1uG9ciVxjdUZM6LsVAbKFLxANdggldUV4rq60VV0h+85hq1o5hR
CluNdfyhGfo1eI2sLFsLZp0Rg3M9a6MfAPZn2Mt9Kdm6VO2Hag670eBiHV+f7Xprz/6TcW1UGQTp
vhLOy4bJ5QlfZ82m/X2BADBxHFYuDRWcoFtV24Xuf3JcmJZv8WDP+7m/rR2wPQ95bQBH1cI5zEJ+
Db1IyKHg5YIN2yUrS/GgIjhFIG8GelOEUS5Ww1XHISvBC95v82sF2hX7QjgTD0OobuAnB3Aakand
AQOS4DiaZazVNOpYc0DW6V7FwnYUxWnCku3AGXBrDevHPk6xbNRMb7KDaXq5RDYjSjD9dZ+EEPUv
p3e0Qt0PgB1+KOCI2FUXeyFMGPBioh1spIxnq5w8wJUdjvEwQG08FCKEcN29rNlg5X1bk7M1WaX2
BUydWYfk5rerMJyYt7zB8xthO5NXffqZU4BUGwkkLcCX/4iRLAVMSV6dIeDGcUYKS/U/JKuUMQZI
4zLwn8dHVClWgncSbI0VHt4M/lfSCYfxeH+7Q2E6SteYwvqBgJUHFAINvBfGmSvzjd/JlXIpAn4i
NVjdZpIedLq5nEHwjrmYh92xdnjUxpSAkKwNwNKQPBr4ATwmiAnstUVcIbn9f/utKczX+1tGITmN
nA+G5IhosNyY6xUPWHWOXTc1wgE6QVtGMLejoQ/oIvmKBg0J/OfKuurd8k8+ZfAL3pX67w7evZm2
6HLD/oCJ+LBG59KQLj6zHtiOAygQPNuWqjx1U06yD2N/pSGergjlqyrFltJ1ZUJLLg2jBWM6JAmo
aRR6xrnJy5FQuj5B63z1Euw8uv0jRTKecIEFDYj1JL/Vw/OwYqTYTyp/hg4xx0PEBFpDvYw9yhmN
SjV9CMs9uLfkALCxKBIyYZa84aMFFqL86fqSBD976Y9UtwbDLIuZ6Lp2BW6TEYAOO881UBpMaGRK
+8CIl8RV6o7f2u3c9FubyrJZL1AuelGOSCb2zGG2ZeUnYtZUOVyd4w2ZNYVgZrcP/MxjSnC/WQrC
KWP70ZmFwmKJupfoGR87Ur3bnME+s3nLIIkNpB2AUy5S5t9sa0oGMVCpfZoe5poa8qWwiK2BDa/u
S5yoq1I3GGXoxNGSDfOwcaoTXWqskxEDENxyjJO/Eu8BEHlvMEEJU2Yt7yCg0tx5YrSa9E/GnTaY
jfxIusQm6iYo6rWXXxQNmG28/4LRY8V4gDMLyPbhAd3WQH5qfCzCHyAXi0QU8TwpRpR0jwZPB7BJ
nLv64cCkV7ZeWOnCxudt2K6757I5hHNQUVH5dh+zMP8gALK9mWI+DPTrcFYJXv6BfBxV+7ccTx/u
J1YezbwNSQ52wEQFYV1ldhDqZm7BOnt5m4JVFo6nVzmjhbWVmkjICa1n2Z28eFwYraIoVJw84aK9
mRfAFqD/A2WHpQrny+s+wFd5O9OH78KNAFZf0olznNPqYbfhmJiCpGn32R73lgygXO7KjBjMCrgi
bNYsIG4bFU7mOGovMjBzwDv9E0G85S5FK7qwzwB9NlpRBs7pAOeZ7mhnGi4/yULC35f54k/Yt3JT
6+MIT1ygcYfoRQ/GGwU6HUm2RerQNsyR6RYDah7jIEvqLcsTZwnF8TqFUfAloqsXyty1UITqZpgb
gxErz8OhkDNxKTu8VHTl1JCRJCFsXHopMT/RPUnuEgeHiagamAIcEWmyS9ddjPbcMtRJ1ZXukmbM
+qIWKnsvqynH14LkrTacRB+orueDAkHhNN/PJ00cV25kfW28FZgryjzaU2zBCUQ4bJgg2r+jcEi5
k3rthCdvSL7/PfIQCzS2gdTDU0FMDaXXDx9/VtqlHiF3N8lQpyARxm0ePDeU4ti9XFTx6vQElNOV
M3lyBVkyGuWCQlfHMUZ3EpACA+Ljv3Un3eICVhwCo+wzrNFqKPwPJWfU3GkL0gTZxLclSQDIjsuc
FoYWd3kzFe9bJO9WAuIYI657mAfpTdCSS/ACd+HJbRZtpuwaLr7S6lGdpbaJp/gATpSVsiRqKpFT
35pngxy3M5R9v9QK/5bdN2EMwchTu/D1j+tSp1QKx2yc60Ep9CEip1Mu+PZ2jY/4x/DjjeR2/1lG
5Liob8xStmjy7awDK9CzlDLluNlmOA7dtlPHwSi0uyV0fNGajgCLePlTrWtmaEyD6PrDVrB4ddlW
6shIyqdGC8rAV6APoyZ3+WFp3ZJQxaQxAzNhZpiQAptlmNRaygbBRa/yYp1ky72GnEq8SJyPQBTM
3cfka2xvcayyFpAu1GVFoKNoCOt1lIPNvt/p1y6n2L+HAPcv4DzCrqsBRPqNa8LvLDmItxgGOIzY
QQhQ9DfvfyHfNkjOox1EWbMwI66t40+TKkfohr8K5U/xllwK4JRjIy7p8d3WCeOaf2mQh4GeZdov
guIXfK7BWLFeZXI1Tjq0h+KRi5tlp/r/mSG1XFnNo2WaNStTkSCLfx/dzvg1c51SUCAc728c5/th
BbQg/LqDZ/y3zFMUxKArYPnb137HCn0mHWf7mvnboxsEZ3xg+Rb9pM+/wwkuVedmcWo9bN5kosYs
AtIOc8coUKb7kAwInv4Ect7o171mpTMaaLJeS3ZC9pjmOqL5lekV+GRl5WrU2/4n/w8TZStvzxCq
7N4PHEpkR77dyi1Qqi4jBXyiaMecaCpS3bHafP1vteYZ11/P8oZI7QMmPajdIa+eZt665Et0W9qp
QDFhpwjy19pqlGcewwCyJOFhaZ6yIzaWyho41zUulZsDu6Qcr7mxul50sVm9TOGHzUwvh/dPgWtC
v6sGvX3yGhVvdQCLczPKGHMbbO/MNDX8MHybo6Y6faJq3XM2FxgfvFhOHmLcX5yYMXXQvv48MYno
PyaFAtaOQvESIMtkdQ8KnZTa019akaQAapm71nIEl/WoOPkc3dTsSa7VEMZClmWdPhvI8cwPPeK8
b0b0fF+u1oj+T7J52+RYVJozDaMsnRhSVSQlb/qtZqbz6A5XMIt48djM0lRuB6TlGXRUky+eM6vD
gNXpQ8IxLbAsmwGmAqd1kFbEIOLruOF9BfgggCyhubs8fEaRxoYRj6Zov2KTzj+V5fDxw4Gk/nmy
3YbkgzCpF2DQLNnSgLsLjAliZbkCtxQYn6iUq4GT3P8MV+08bB4frr90J2RqTj0thvdu3xP/xDpT
C+LI2odnp8wwF9euLeEC9trKiMKj0ewJKefGBWgoIyzo9uX9GXPsm4OCuRlOse5fjrHqcHqfGV8y
ahntG2MAlV+Ji7VYWsIsaoFlsiu5/j5lxGoakeZBh7/AlXC6q20pZKL3pxKbDHx6XSvlnUCL6996
2s3uVdRxNL3D8ywRjpFi6a4hF6UuTEc+tJ9N5BeXXCyvYxuw/ZWwTTtNQQxv8UyekCscmM7jFiz5
D17xI595crN7QlTiRUnX5i1+aWpf8J8n50BcxjuN8xNe+Dwnbsw5NZfm4q+qoi0rZrS5kP0Egcji
VxpLqsVqT4q1o4pnDUXiZLVX01UyENcZu3LytsvAhtXYwswl8walJKeOZpKMGnfo0lftY+HK9YvC
is0Tkbg4enjEb3Wxb0lXxEdmVNR05I02Arhevb/li6cZbjmgktJU/bKL9eG0qoewvnXSNchswvHV
K0NVuhTMLamP5ofueApDV965CiBmvbc9VWluAcpIL3bz0IB8Ar3r3LIxsVUm+w5BBWXQax1Ndiwe
Hc/JeN/6D0RPdm3Fz+rs08LfqiNIxFw0hJuevbAoBJjE3U2XVB87BQWiovVMPflv90c5e4ul5HdN
kDrMC0dv/zyuJ+uH0AaBJ10gwiKaqxdZGwTuR0fD/mJ3VxcxsVUXI0MwzZIIgumWMONJgejbQN01
pfSN80mQzG1CNBhDHdSfND1Dkq47TzFwV0QKToX954cl1YJJQ5LXV8RaH6+zbqKrful7Qh6+AtHl
DElOrpPQMAl/fT3K+9BT303LiFIWIzgXUa0LJHolIaCYP6hoLBwCcwcVyiByCj81ic0EJcWceS8H
dDnDh2blCCJCbVWUA8nS+Xw1TsIHP2iHzMoeQj77u6wzUuO82oNzWmBltz767j4celnnGLbGih0T
LHgTvZk1upDztdf8i1pHdsdZD8a+ZLjNf7a/VtT9y+d74kEPsJKSiUV5jJiz3KcHPywKs6ZVRzCp
Ay6E9uRC5P3iRuAfTTugCOS2VaK3rdrgbI5ChjFFPPIYQXLSiJxRVPzfDOXTjT4ubmS3Oq8l1sfB
P2OGvj6+SdO4dbkvrHqWwKInEJ8vWsmej0WWwD0gqusg08nfi6ofZWYKrMJpxCqSVTI5MqD9ntnp
O1ucFCv/8AUHNRbj0Pv56F6DRQ/CVKqct7WvK7qK7GIgTkMXXuoeu3Z3Rd6hhMf86a1MOJneqMtZ
06vno8ljZY4/1p95MA2ZnKmjyOnh5WXf4iT6ONQr65B7rnQ4gRE030CUP0edmST7qXHebcTuqBjv
k0jhigxxr4DtdvHoMdqhOU6vVunzlDuKZhpr03+N8c6GqG1QL9olUEfU1AnZnGJ4O2v8foeyKL+S
djTLy8JeHJfvyimNH/18xR9OLnN60Ex7sTBbOZKiMUJF3sMFnOW1ysqEK1zF04ZXX5MvuNnvBLd5
YOC9p+kqn1wa/ga6d8S5rHsrgUdsZ2m9qVJDW4vn0P60CSW5FMXydCTp4Y0edtYoBgL1WCHakIYe
DfYD60kj2NkZbYp8sV3bQl+t7gFEcabNeE/aBDwIKsAqm9Hh/qTdauaVtJwzOb3zYUsn1Ob++v86
nsDxkjL5nXYJpowpFdQPe3lJwOFtrkQgpnWL2EofNEmQu0MtPD+iALEGEl+cJ3i7dh7cDGmVfiAY
gWYBJC2ZienNnegA4iK5Zfkoox920cQuClAddzpSwq7e/+gbvO8ehgMeztWVJQXfybWkmDTg7w+k
ylZJ4aNagIMoeyBb6COj56WoYKYnfsqC8cBfDfLrEjUu+Gq8C/chlUdAs4PETZWufzLK7w6Q85Qs
8GZ+S/hU0l8cm3ppzUnYQI5lNxgVJ+gfckVWWVYD0tqbKnR99QQJ4mKiwEPMr8UJXmscWvj31pEb
IsUkr8NBbEufyemBfL1C8njdXORIIzvdAd5mwNe1zVcAH6ymvQBznxCU2bRmaGl6UJ5xJ4wys09F
ulnEL7DuNWUO8yAGhVK977lcAebrmXutU0e5RcxEfTnwsKaDHunGOvpSFGpuPI9f0hJCb34kJJZ+
oXXpLflVfnCKVc3pZDomZyTyvpUOzYOpwVG7PE5deDrAL4eLjYNWEhguQcUfgnUqD5g9LlD3omK8
kKsIHxZ5dEzXjUlqJoB/L5sLER80nk88r2EyI/EqpXaWCnfc55AuQk9ZDKeHPl4T6ILr5kUdAHFd
O2OhFZhWLHN5x1cfzm6LRGWAdj2Hp1frddmd7nbouZUGL8r+0DBHfMqYfPJQ5rp+/wgWSh6bJGbR
8uxdqHjLaA1amOp3fZPClLPCBG3QJwf3H/Jio2APFHHtzFh95l8yOaMzmXjRNbYvCS7n797I+StY
eSt+R9gMkzqYV4O5dZEZIFVG1+qldxhFpXy118xzDBHtRu7RfqOkPeNyX+R+9PLIUnMkjnL8oZeh
pdowYP6FElLOqOjBpmH6GKfJcQd3Bw+PMCADNk4Ix+MIjrebZP8V0TenTnAPVs2CwBpsx+LRUnrM
asO1D0miemhi6cKcbOSNiSsOFmUNmwR3GVnU2e1Impj4b3dVRX2DHmd9lhvCpdXwyU8S6TqdAf3e
05TSPltP34Zxj1nJHDK+/7fC6T8E24vF0cAgS5KNsKCL5Tnw4nTA/GAs2VXZNk0qSpC8lPRP1ryC
WXS1nCC2nC4yq3DPDIz0/MAvjVnv7fMBorMQgQV5F/NfVMlABebN9MTdlSOd8pFtjPRQI1LYTMT3
W1Ttt8UqwN1Q/zv3QZHOiiMO+OtzdVsyrEvf0NMHXB96UG4vkQOCid53hmNpKhe0NSCCUn2yvXMJ
+cmcVSDNDM7K71TOiDo/m8gPFvA8YJmIMTdLR7YrRqygm/hxoyev6PQC+8wDM+oq6/gJiuOvty2N
6+GtY8qOou3jXLn1hg4EdaxKTDqkHPmZvJhSOcZ7AxQRrPCnRK0B+2hZkx9ll5p2GvZ+DEALOlM/
aE+0rEsRMCuyoGo+8+GFGCCTN7h7a5WAFzjKsmD/tH2m06+kaW3BvMVbp/uJhVUmAnKIiNCEaZsS
eqOO2aA+KZW/lawm/1l5MTpocPBV217eqOQjQglJnpUGf5Mdny3Wut4GaimYLWpx/FFl75HtlgC9
EyOOnph8Vxtu3nwlEL2TTvCwUmZn8dTk3jqnr8L/R+uTBnM4qGXlsoS7kp0UV45dW7qRA7eUCTrX
/e2g3uPctcM6MfbAC83Rng+cBX0EqJyMHnOpj7l1t/JD1/wzOg96NWkyRsWhC/M2r+HX52j4PTUW
hvXDsNXJPFpoLBcMaSq/OBqG1A5ukI8o6zf+niglhfFoJR8IT9onfaGKJhuspQiLf5xhWg8jg2UN
Ka198KoSoKAbXoncUWoI4+2964ndwY3x/3u32uYWoNjVNQsPKqIU9G1YTX6GpKLZx4cHMenAGskI
P6rCTOlIjsB650DoPAFRHzI/+rF9kK5lRRa+YUHz84U44b5pAB14o3LIxdYj7XHtLNz3T4cKICj7
FL77Bty2RCZa6KdDw/hdWF4XlE02hikadLhWlVW3vXMJCmrDl63BVX3qY1OWk50AxJ3YH60QMBgA
nFwOgWDkPKlWpIoriLxDsitf8HIf6U0b9/3LrK472p9Pcpjlu9IU+sf8WidC6ky5D2DLTLL5qqi5
iCp4Zu/wpOWdONRH2DYj4c2YJO2XLCWesViNj1wrpxK932t9Ux/1HsWmfBQuBFLIsBm+DdJ10LFz
1jwOxo5p48s+BtLKXIMmqs5FWBpErEtLJ+sjTbHZTobi5wRjvCt7arrD/5RcIS2YUac/Z1zh/Rot
JUc1S5GUOcCoRe+rmkAZAU6mxBpbM63mVGF1Gdu6dNPhHk4+nBQqWAO0t8ffno6FkmzNduteKdH/
NBQ20MApg650t/vxnuLiLs/T5dC+JFviCcPabM+6AF1thR1GEIEjjzlkaDXDD+2j6hDMRAfcMb8C
m6nVNS5HF626jG9BeWjyYZLuGL1gbVGh17WbkVeh0TscRqHJGSI1s+qXgKS6PYvZL+4IgAboKKNU
u4taV+CMzER4NMJCxY4+KHSh/SeTSiDhXJD55lJ9emO8oSq94lvDcMlqxbGvcWfb3TS91jbqndnr
BPzWfD9QF+7JpccNBR8RWwt9wb9Lv584F4Q4Gq0Ph+1OFKfXGULBACeJG9gtEB0pu9M6kqKjlxui
yx3ufDGBy2klBaE9t/KEKYYRhQbuId9ox1TmHDuFoSFWNsJvNM4lgM3kgzo5q6kRJfpWfMVLztAa
+f0wh/9ytOOtwhSPdkOjMwqONFWfydWOetxu892/rKXghfWwZXv7YgVUB2uGvAnrpXXgruGGtvVN
XmWer+L9wtPxEsdgM1G3QJ1duLTJuD3jzGMOgFSshDLpPsH+3M5XfgOgwm63G2OHUBeevtHtss8t
d1WG0arzTwgrLhq5hwcyiYVzfRn+DP2mG8c+z7vW1FzFTKJUobq1zXfyRYdxar26B+WwhwGPxs6y
iWhZ63DcMHBmD0cWt8W4KpvRl2/x1AYycGLt3OFh7L1uPoB1DbnNJijgz62WdrnU3dch84cjKfOQ
3CnoLmT5lua0az3hiTXOnHfX9RtLgFnW9dP+Mn1BNtawW3Wi8eUQhLaInAo/USeX/bQ/C73g3Mzf
cmu+EE/skEfEDWilpu3X3urxPEwmxtUPwWfA0bzXioRofUs3d+Dzhnacq+xQrwMH3hVESawMuUbM
paa24KMz58G+yvrWcco0G2LJDdBY7CcTlIGdLBTpRKTNm4Kz//M7o6ZS71nvcmjZHR6jCxwThzDC
DNlY4UK8p9i8ujoBnizoAV6y3HMHGI0IyWvYwnkFkluRSuFEg1AeAhlior98CGOvI/Dtklq81KV1
aLLUFclh3Jeh6GCAm4O1lDFpsxGzjMZ7myNRviDpvBRQ4lQEqSOeuZXf4EaVj/pIQMubas+Btg+n
ZnTWGBbsLruiye0wzTzgOLNfV6JYN676ofDbbG7V9M/eY24Tk3e8c8fV3ka/uepfJBnioiNFLUDh
e8cpfWHx4Va/rS1eVX10XWu7nhKtGxQ7u4fw6tGmPpvAKiJ/oNUOgZmarsSMFRg6NSkuaylT1NwV
N0uJgfORSONBvprgQEgwaF2MXSEnlEyvwL36uPnPlXOEnYrGe5X8YVMc6bhFw9tXTJlNfWLY8l2s
ZZbgCIDygVtNgPek4V1HyhhvZUV3I9xk7rVbbrNq8T4M6g/Ws6hxRs0OPslfVkUQIFshnU5NL4Dy
DhPiUjmt03rSaTBJ8uaP7IFRsAbkS6q+nhGNM/Gc3X+jSe+54ye0yj26Q4bwgZrpVrf4J9Jro3dd
qTvcrXHbKnbsAtwNar0s3Btz1WBwavGlBeZselxMyCyAk74LQiO2g2PEZ8Jc/S9CREeqDaPDi4TN
sbmVoRZxWpFy+LSK5q3MUXwDsz4Xml8xp8FPRcfdCRkE9IhPpZByiJvtHhhKZwZn9HDbCGdYujkd
ULL31YpRp44revSS28Xu9MFtFNeAkH9qdvigDZLA2IuKwCaN4sNM9zNvDfYEbe2HWq34+Dat6m64
xtv3mz0shOAunLQgdLCEmn2O96OTcwz7wIgtWsOQpDjrLIKGA8ORGttMtjRnyGeaxv4viPrxN0y1
RZ76H0UISsdde1za99arnR71kuaZvWvNjNEJegxnkK35mTUBNDQeYrBWFDcSAoQhX3vD/csReJzH
S9VUZFKwHv/bXQ845fvq5KKe8UcC8EaGt2xwuMS/gsZx+njZdlqmqPeDWBWOAlMRFQi9/tyLHoyC
J8g7lOO4Z6lTF5Syg42zdvjok4qFQWoEMSk4p7f80niZGEXzWOCWlN7GOs+tSS6LueehVCQ1xzOp
gGCd8eyvchoSIaSXmz/FD2KJ2db5EN5/6Nx0ZOFUB/6cvGdEkEJ/GwDlOCf4gKgzstnre2feSASK
T19vdFVm9cF0SsBPOXos8mNk3q6k/+yajeKwqvFU1dzXMM3jh+e5oD2Gkthyzt50Pg9UEP0UqOca
sgOMYLuJwPOxbw/hms3tMBUS6Nkjo83xSE2omSKmk5iudymbIe7iR6Z/ucYK641q1CDQ6i56U1tP
P/1ars86D0GNglE4CiL7YeNpGSWg7aChU88p+TSwJuV7pb80xF0Q7THG/UrdEZJvMFQ9jUwxM2Mg
XoB5SuIQ0Bvx7fphSSOMjU4EpK5jFITKh0l+NyjAKGUS5uO7rJwD5IxAJrjgFg4oqKjpj0VgYF9x
FOR9X1GWsdhQ0MRLHx8YqEGBVXWP8Mc3XP7TItd0QKlLfqwDxF66bkPD4NGdUd+p4EQODn+mGc8c
CXzqSUb6zCd9x+ePbl+MtBQI+RI4OlhjO8OGQcQlZi8J4lH3W1bsiDNezMzPJHvjBFTv9dEH2MYy
2j/C2md7tsvlkg6ImTtpgNkf8qANAn+ajS1prP4ZvpOUrs3F+1dN1ie9GTl78pnKBAWW8GisCRVn
GTOND6QnxIFBzoRJHhjbZwdseGICu6VCVpDlZnCf8EnEFUffTvLjgfw4Ug3r/mo+7KuZvgp1OOil
gH245tfw4WDDd/vLdtEzb0+3LakuaKvRtqXA5FoaVIL+ti7dftzVV/zCP2a2yxlTTNrNhMbKUnTn
xmq5ZTer+WqTM2ylgC2s9WEzMV01TFQKEa+nw6DRqD0UqH1vqQX82BcOzb0o8Z8H+k7Qre0bp84Q
dcPOTZx8SVKAWxVJn9lanTKNfyg2sTWxYVffv7ckREzFQk6KhwZZDqJB6tZ5C5vMS4w7dVhjiCLq
BaYcJMRK5lEGPlyDPiafy30Wo+ZugIOCLpJ25LMNVLUuhSMeYYXQO6zh67CBdqCy1XDgtATD8Hle
NbHzcaNbGcdlSrKlR78bP7FMnbfiYvlKr3yXbBS9WXIkDiCQzqx3RhAOwiBIsu8Akb/ZkqhINvNo
9H5oPvVEUpzvTFv9AwgS8Wze0sBjm7oCaCgVuun88GgCfMqLh4750QIBnnY0NjrF+kr8rPxH2TtH
KGmo+Q6HEHVU0QqyS8rYsuA2CxdXtqpYCW4hRlPebH+EOavqdIoQIL6YikkmraPnQpuOVPiZS1p0
6AwYRqOadpFMRr96th86CM7gKDG9+K3dp0N5RITRHS4ps/88KVcWWou3iVaL4pLKjbe0ikH3bfYh
rybl+OiYTQ2iCya8uF+uff+WXN3vsqjS0JoLuAcv4eHsNmwE+heKY2zMQjdgkkIKHpjOBZHOp3xf
28RTrF2Pul9FCM9A9wqxlVv3SvWcSyqQOZJ/YOiDCKvS0HMRmI1+Xolod+ym5bV9OPLwV5gKBd86
qf0qnbkz55KeuMYncBcxtAc+ZqxoeEHj8pIARZ+JdcDqLwbZFplSEsl7MJ7x6Nv9NVxPnaTsbMQs
uUZLJzNcQE0+rLF+2pY8QngAikMLq4OwaqEHtRAvTb9iU9WstlVyGDSOqoBCsbxLTKIvglHUd23/
4rpNwemlkSf/NdhhkyM7I6Uue8PdrjOaQWRMHBJVzZxdtDAebQ2GJz12p1fTViQJe/46tRxF/lhZ
sMXLCN6aE5I01ekqyx4flTj4cVNrBw8BLwPuHjoEHvMvwaxkYDCmNOjWxH6+7zOsMIeR+x2LUhOl
EfddmvEBae9/7B/++jrXkRvOD0a/cVibVbMt++DZnhlS0JTCtxyUakEWAWhIspulGnm5T2OCKHOy
K/R//0BqnSftKNVjiDrxp3+Rn+cDU1YJxrQKAajODyljjp5uXaB9u7WBpfBngEd7St4Nd7a8vplW
kjEoHmoOnuKuAsQCXEXD1aQ8z0sC+tUA+1N1NfsrSJeGoj19HmfQp3+b1Vr41HXNJ7Tau52wTFLB
SWO1DhFKtACqMAOPwKodPJr3tRtj9JWXAvjjoRgbizLaZrGEHvIx8UZNjxtKrEwkV6CXtgO6Hvrw
FgUX+AsrStqbYM5yWZv5ewsfE3LzTUDqxQlFhtc7m6V6to0IxoYl1pKFzmvR0ZBQkuGubylnvBsB
ig3nSo+F5Y9RMykH6akkFmuHcnzDAweyPFfnustS1uGzhJVydh+LtPDshwKFPyEU159KJQ3LAFnY
srhAhjn1mSUvYNkmQtoR5m5hut4AryOH2E8qK/V1mBxIcfa/ns/5xd5/yMes+M9nHRmS3gtc083K
A12fR1ZH5PpFbZ7d5JxyCEJ1H8D1/L08kzi0hkO57XjFgwqe8Y51ntdWjNXS5t9xPumqNMTcCRJY
6DgY1aeKMGvHrJy4cg3sTsmw0DnwfLPUKnF6LFW77Eq00YTeydQQ+mDT/tMYu4JKM+pDycNHft5L
aur6XWftfirEHkkbKOcQxvRVOlwxuW5b1eXK1O/B03VQIB8xKl/CevbeQIQurTG5+uYoEV2aDvqw
BPi2+oIMv/CuxGA5Pma4R4t9lSFU9DrX8IogN3NC5Y4bIFPaB2AahkauKf6it6jgze8MGJtQ2V9y
4cvDT2NCPv9JhgwUGg6Vt57iqz7i02iDE103j4R3Q/9PFVJWugtR9nrI11dtGy476TFqSwZwnfDy
YOU+InQkZLo98Evfe74+1dUhFkbaTiDYZ5lSPR9hA7DxLOlTBniMXjKc0O+5AkQ1bKLOzAVOJo/s
Xk166RCZ0ATLQXUVlDcfMeU4yKqd65HkXwQwedwCGwAmLYfJCYyJztpNWRQf4fXQc4fgVfx1SDuq
EQFAJoCOgVofOSbVvhSw1E9BV8FhfXx7b5tniD4zpjXAY+hCdkwUvu9OU6idpno6oR4ulAMI9YP4
0FEDdLvqkA0XTRdLvQYIXPlALL1MKrbdpGHbbYqD/KmM0ST4PM4mYfdeLsVQyl0/LnZbPdx9tRFz
ydQuie9d14scHec9D0qjEYAQW/gcGl/q7ym9lgqLakZiRJW/cAe8s23l9NfNt7sGZOKCEu+SXQTL
CrVb/z1Emg4s1M7WxngEjncuiSSpFB/2BDtwXQ3W1vYi7PNGWAIoH394fqyjkEfuv5hU6LyonK7F
E3QIoZlhD7WhETcVpFDZHc3sUIM3GnHGbC9n3ywiKPPuMLUW3q4Gsm9+HFs8IrxqkP5021/S0bSN
Z+5hKvvxHiC1E12mStyZ4H59e0jEkJy4sSxYkSO+ax66KTgqCHFgNILS4kwO+A3wNbgDwDTdB9Ps
WmZFBOH2deD6Uk1kyw1oLZ1Dxp4jed0XLpGKk9tzW4X03oVCS6WWrrFpO/BFIb+EytGmi3qtCnGD
VDnABw7aLYGAg0ANLch0Bk6VlX5+S7a/6lblFtxZMoIC4e9svZQzqW4r1/VhtyUzdbDvSfINkFHs
t+ZBADlisIKNYhVau1RbfQgUwsC32UbG+vjQkgb9bTT7Ny1GAuFURb1V2KJ2wtFZtj2/KHwTAfXy
5tSKqcsCr3QDiR7+vVYLEMglF9+XKPqp3nvE0KIYbarF4vDXvOdvSy11yelqJcCmW5/lSG4dMWVI
oG+S9sK8n8GhQUEqezmra5PlMWJgZFYjKQeXYU50F0vvu/zUYLa0C+62XVBz5WLXUp4ovPem/zhv
M2e2nJ4YaYG7j0BWpJyUP16CBIMAcmfHf2yqQeNUbXblPzIoXXc9LpsJ/xj6I3cnkvk/TMwe8Kw1
Yj7gA3oik/JGELaSkkQBioHSizLdx0Mk66BGeSn8aKpFDQJIOiW65uJNf6P4B7jXop26apfXM0Ft
snQFiBC0VmyzgW06TcP3eQSpKl/4KBNhVlD7tayMdY6BpWIaBHYpObzVUy/Lw6SM1P6POi1tVCdE
XI6zsqf3tI68yyR6/XxTE27yNrAhP1kIaNoqUbiqdN2IkciUlk/TBq8GB3yW7Hvw13qygMPSBcuj
iY+PWxvlDL6BEDt5LzQH5fTepri97igbnVchiMJbCJsGaEcPM0xlfM/8U82xJ9TgfXWAqYCkoAgq
aEbSKyzPLFeORHwf45vfnJQguyFLr+nFggmOC/w5eI6UFixylM5AgrV1K4JRa0xNKxu3JiMSjxdK
bR37EkbK58uciSl372Y507e2iXxQLi4R5veA5xLoPvgXQwzmn6wsHmHPFiKJYtk44Bn+6khWltIu
zL7JOxHu3ff3W9XVlFZBqWuNOvqn5f3e+YhMWtvCQRMt/GolDyXo63YUvHATMo+VqrC6LZ2657f8
eQfGd4C6Y7a363gaKOYWQrQHHSShGvEWytBGt8c9Lxr48RrD4NYENMhDvDmPABeXk3m9FSPnRSta
LLsLbpUrh44ImT3p4sS7PJWOkTSaVlJ24ZZIV2V3O7DDAoNGf1C3MzVGt09nm2iFTmmRZH0+flqd
WVtRoHf0NU2i284NWfO3obfHvoc9PmSfesKJUHJ8u9sPohiV+bEGi3P94nSWsNzJZQr4QbChrqLM
tQwRSBubmJX9MRMK3zEkiTbGSzF4Pjw1C8FJqLltO13p2hASqmnPEUOTVQoqwhjE7wUnkVbseDPl
aTFQT0R9zeQXwaxlyKYWgeB8FFUtJVoj0alQ4+wm9pA5AMqPla8tdDVVFBKmFOnfG4c+/7o51Vv0
/BA4082bnG9173TZteVGN5DV/DcQxtGBYMp9UoKQMZNVw5FM7QJBWIJDSnWimXUsXjapCDMHKTV4
SmTCiNM3NYB03PZTGD1l85kg2S7YsuHCZBCXSZ/WBLXOKPs5ORgZFwNmdNpyc5t7bXUFp0B2v3Q4
jMp51Bc1pZIDikuaRblAcdJRkOb1BNk0kVUKRlXileVoBj9Cs9yc/T6Mmf0Lb+b8E+yqhowsWBFt
sZ40SwXnxclnzeMhr1B+LxIRnp4BdHiBoxWPNb4wwmnWGw3GOplYG7s/GT0EVnPco3NorFTqXcI0
cVZCIvrijj4jqJBJl9RVtzAWcbt+F4SZlxA9qQ4tQ3hb/MJ9eTijD1+KV3kIihk+U3UoPZppWXFz
SN/+F8/MgFIDg7yKvIFIxlJK1qsnWLFtZTReNDlJE7NE+qRSyn42BDfadJtPAur6dqshQGt+0XWv
qs47ixs3kD0cpl8ITizYA3KECLIckIPc9eLdc9oSOPgAkhiK8koW4GZbX1yNBpaYC9mf2zljNUhJ
/RtuD8ganw2VA7NBxrpnSV0y3ekzidiey3zvUngFQ6Hp77iENWGrNJMCbkIN4BO/lQF4jlgZWwWm
6CCIaItC3Bm5acp6BIZxPM5PTFUV4Zij/izOMuvBQmvTYeyEdj8k0oYlCdPtKyWs0uXE/ihXMzZb
djKPoR3KE38eV1vJgiIzbacVvZOVarRtTGvoSz913AcosD81pxkulHP14UVjvMGqi0xw0YzUtaxr
oxzYveuR3dv1eWKHr1ZKFNWr2juG2nT78INXYeDGuXbrQ6jC58lK/pRY2yWOS+KGNPCOwFX6oSC2
ekf5yoIGcue9jsrieVA+AIB+v7PgF4KQAhG1PkuvFjmQo6CTt50bhoTsHQYAWV60yYxzrWNOIYoj
xHN0gRl7Ql4hVa8kEa2yZY1DFgeel8tHpwF+3SPa7ytbjBvvneJB+0msurwuMp5NyB7xBCj4bRoh
nmtAj19oSfWeL84un2J0HylkNuxp8Vb/8kkO+fxjAObTsAHP2zniqsCb4iwJ+rmII6TbLnIedmar
dg2h6QIt4ijGmCpHiMd3oftcBYkP/b7DcVgiJV0kRjZ66h9+InXAupDN0G+Vvkpv3qTqKSNUdBYQ
jZ729lL3DdyEboYpS401tQdKpPsDyov62KF7mKeZ2iOGeZbk5VNL7hLpiE8fcXtDe9lAGc9g6Q0y
Kmrgy3j7SDbXwZ0U+edFS5a5HjJmfD48H/Pebfg/yckQ/EQHEzjmGg3AsmsHa6158c8Q+dl9tvzY
dbfFWAJv+heABsJrNczKTGyBpUnqwM16p5HbhRd18VDIOR43hgoOCOnP/P/KwaxHQghpQUIXxRSp
DGRTF1zLtzTEeBHR5w9K3AKDz4Y9Cn5s0moMpLxrwLlGGQYPVlwZQjWBNxz+SepEmyS73CWsDS5x
ZRbqim72Krx+w+G6A7OyNs0ktnP7gs3XGRJZKDd3KGrRH3l7O87hyHhIg4dR3VRs3KoImlKUgLYs
dEVO/TKphORqMUJImisH1R33BtWfmib6SUZYHzbAiIKfTVtTi6VYC504gBWZEvdE8mkrw7uXfdko
Ow6xr9b6ayFsHoL56OvZ9oodqVSR0bLcLJOZihRVahSyfHNGDJjAZkfFHRGVZ+kQv/Y5HhtsmR3s
1Qymuil/wARQyL9DGhpKgQpEkuAZjnMjhIQg3iU+IQgwDVj3JIrm7AMmkQqHoLz4+8RVCCBUbmxu
r/CO9frxQDpLYpZdnJ0Bd1WT6cuOP/c/grP8vif2vBaEf3aEyQ9USFLIr/lXUY25tnQtM7J4mcMJ
iWQuljowSALhoYckeGyTXPmWGuA6QLrSYMz2bO/ZvgCXrdJv6HYTedfV6jdwEaUi+LJaTjeY1Z9Z
Ic9vFNuDxK/cqd7m5pxw2KnIBnz1HFQWnc9bq69N5hK46sq3faQF1G61Jejd/hkXqCH35sJSDo8M
+bu38KkY8490JhdcPO6wNmae7vFYSmqQwkzrYsKHDTJpC3eeoz6HRXx5Gp1aX9YjPD2oZkUjRkdZ
xNYKqgJhSI6GqfkSBXTpjnAnxPc4LxujhqU68rfz01qIV4FRcu9Y54eCU7NRYdio5xu2h3mYxgnD
oK36EOUT3AkX0sBlBYenQ//rL/ThBGziqGjtbY7aAwkCLqeqnKyaOeB7GgCcgyI15gGDApMuGpQW
dijRO68p24WcMD+UN9GevHh0H2RwbvJRgQt7YVy+DZfduh4e8v1kgC0EE+hkl/htzrXY66xV2Wuh
+s16HLDcnUT3wn3BTKIV+zu3lWeuFbVE9wxt7DzHhNUFfcwXUKuUQx31OatZvedPxUZGZySdpKKD
T6oOqiHTvyr9gscHci6vtKlMELG4BTuOd/q4tULsNRKwfiMar09RFccqgIwFEdw49cPpAI0pACrE
s+lu+HppGmiSFxKLT+FN58hbrYkEmURKi8BubyFOdP9UvEWQ4tG8PZhJB8c2kA44ZkEWJDwASIAT
QvD/lN4QIENYqu2DOd2YTVJQKT6xgS+tS+G49VlFWCo2HehKFq7Os2l1u7f7T8RMc7Jt7X9KtcKG
ZSFSrn4mkpyMSsvZtIungksLR0/AchUBNdayw1FacSrjWwnWJdGZkSDSjCkz98ggD+MR7CPdjUJ3
8bOO3Q6dWIzt7OBo768OpwOfaUqYqJPXJZIfm8owJNbql8F6CcUuOt8vxPpuDEDzH75zezWGAIDQ
almIYHu1B9HRYMNCpsfTjR2L9krj1kZEdQOIc5t58tn0ctEqxGxtOM7yWf7noKxx4Il36IcXca6r
+WD3EaHkeCgrPH6T6vIojzw5H97j9WYCX2MQae3JJrFW67gtOOjvngQ/lzZHcLb8MNEObOn4OYLl
e52pp11hMgaSJHdyupgYAjATKboSmbaRAYwbhDIZTA7tAZjc+HKEuhXnRHfPk2oSEzI19jiuRPmz
FJTdbaiLsXoz9UpOttiXTMKQAPVz11XDT6uveHlNjQBMYuG72HkQNbezuCqs+SalT6OiqSAf54gB
CDnzP1zql1C+kxM/EDLpA1dFEzo7IVT7xBuzMCVq4/s8FE1hdZkeI7JTHg3X3OEkDGF2qVW8ulD0
ZSzQ6eq/vCI7fWpjpPdhiFQ8kzcT2aUWSEEIO4j0ZUfnKxZfI8N+l9ZAJnVj4LFUwAch47ZhtJ2m
dilBPJkUfFpibkVI16biikNXCmuLP/CumJSQa+9fBz0OLiFJoa4g2voLErVk3j3qDCy6kAOddVXr
MoaHYnhMMSyRzO1C9QTx54s6j81XxHraGdsaTKXchboD9tnj282ioxRs6c1TxYDW29kRhwI2G9ix
gweYCiI/SUL1c2Thm5hxJh1pUDOfai02fjUtMDk/+pvQeF1yYvjRMzpR7qofdsAdvsjEFcu3fnlq
4hkmBE/0Z0xBBGfEIxO0ah+BvqpmECMSerC6wUO1GQAVf8QrGM/8UyOd16akWKhPfOV8mn8Akt+I
7QEDLTk03lsind6tN0ntrGBEFFGA7WiQW2Mv53EAHGlb8AfBPoClWI/cPqtT1f4A1flNsb85lD7C
RkG9CARckLVYDYOHNRQ6DJABa3MCb53ErM3BxtrA8i/ilXlJEszQBc+iTRrM0lez6sZqXuRzYZWq
Lk1Bk3oR3BESYVcOePGWI5gm+L0dQFbXgeTriz4rawN5oj4sL8IarIAv/t1lHjYQ9kWSOFnIe15u
qLe7mQ4NMwuKpoxyDRf9u1PmjPUBrR6jNGjPdyu7UE2ZcRWV25FFRJDjn1A4Cn0QYINSQ/39p0+O
Ij8KHR4oLzMNwV3WiwdE/3sIDhKvf7qkKImwPLm3eitH/XZxsUKSO+aqIXNPSmx6VohkRiyDfsxv
TQy9G/B9psPEXWC+9HqW9zo2P1rcFl0fV2AtB32yL9VtQJnstSOoYXZe8sNTtAm4LWUQQGMRX9HU
rRfHowj5+GGO3FexDBE/07gR1yMghxhW5xt9J7Si30lp9B5Lf1HK7pt+cYKUQAGQQbeIMNfzoblc
9CsD0JR1WU31pMv3dnSit9eIOYd0WOOp8GIVTIM6/mUTMPtNwSRkuj/29kyZYNUiwMN3Gmks6GI+
psGlp5EbkvCRDHqplMEsbAcX0SpOFR6Czm52Sl01UIDFonzn2cQ2KdqMRFrb6eMPS4yxkG/Npwcd
dDQeXEu7TEz0UBZc9iPRpFd8Wz/wqELp4V9LIvx65mqdi9H5mugd/OTyqox7/dH0xTMtyzwnKGCo
6WH54Mprx0ER2hjv8qh8BJychwpjrFL8VVhzjCVniSTEbqwGc2yzToSvv3Zpg6gIXSn8av0WVWW1
wCZ7CLYM8C4PQPMbPphJ2gQtFQGAk4XonTA7E6qor2dyMpnfF6fsYUbZu2JY6VUzWBgGfKhIuJVA
yQw4LJRh185eg+VXAny6dLcl6wWfLriJzL+SHNFOgM8vlpbRyfLiWhQLMIvIpe9fNm0SASvau7J/
7QQSqj2vAM6PPhHa05MExUcgoF3oNKva/dDeAa+Fyi5Zw8DVHk+B1wzfXKdv/jHkzsC/Zlkp0H/6
0dZ0DvrFoH8aEZrDXZdG9vy24Oj7kOdJMUqkVsDeFMweH/fBjokPbFzUix2Bj8u5eloDTZY/VEiJ
B0NDHcImDd5+PHncdBGbKoYpizuiKVwNS2GnG7zBvp+XAHncZp9Gg8j7C0xoy/aTYppnJfkVHuCN
cznEjt9KunJD6yz1AHFxoF4HkOZcEfRZcwhy8RzGbG6q6MZwkQ83Lo7/gep2kl9ysuNOB7CMGqH8
vAyAOnCwee9Dzlu/i+Gjg7LYptFubZ5DysX8IjVJN7BbyNFjWKu15YSt4/uJPmHj4p2exnoYoYAt
pilBGFGICRHRMbkqX+wh+f20PtHNmt24VrWpYSf5IbIjGRpIMBHxiFfP6oomXCv9pHCJ68th5RTB
xUvRYvqauJD7CnO5VJdQKTr4Fu3WN+tFmEZesR9RhYxIfdfGyEqj4RlcvmeOV9SHqZIbGTS2cRpn
ByJrimDoyiohLfc7VqtQqcKL2I0HSlLDrWwLg+MQmgNfcXmYNLjifJYI63mmhZRdL8e3vKQXFgiG
TZeBgxA9s4vWfavI2cIZEOBljuHGyFS19lo5PZm9ThkNucibGPgkMU7lfNYk2f32GWlJLmyqI/eh
boTxnOWLl/EghMwYg+dIYPkPz5w0FQHgRjc1LF8D3FYzBJeShq9jhKkeWOXtWa5A2FsyG2qYcqD5
E5lcopy4iTWAZGdsGdqhTBrdkqqVxKjqKBhNhEianffvyfWlLmBCa5rktNGZAbAP8Lt3nWr1Lr3F
19806wQgfHm5H21kgeHjIsjzlZjlCVwAncdLCHJkApwryhhHbJi910yDdyQyjzqoGN3oLTdORblD
Yo8/X38nK261rGefffFQ5nDTfSFM9h8cnFpT/2fYUnSaHe+w+IceUKbYQ6wktuY4tdeV2QalBBI3
qohegbCer8ItRzkRRKVMwQ8ICvdRcmuFw8j2jSbeUeDWpC65xJIushxQpo86p5uvLnlPgVd2vKTn
xKo97mT2bkrkKXLeFFsKLEgulSs+Bx6o9VbGokjgUUKFMzPYoRjfgW9u0or0p+OMOwhdFXfMPhXT
iPKqko4MFJo3/idDjeCsdrh/zlLL41wP7e49UfL/UQc9aya9fFGsog87e5QTrtTpcAN7GVAxKDlo
2YcFssDO03f9Rjg7JI1vYZE/3PuSAD0hzkBz7as8RzC0zmVUY69X1gAM5sPO4MFgSn1a4Ly6URtz
c/NTW4gxCdhDwFT+JiObBQF1j3je9+ueLEz2E3ARcd7phfryT+bftIhqjnG+Mc9GPHbGc8br82j8
/fVAKsHVbxBFtaRGCc78QUWAHqbqD1JcWxJxC3DGAt+wQT7Fu1eu7n5x9glQBf3cebmlkayjS/4r
cY85kjWa9VHpS9ljMV9d9vBpQ9YuXrdeF/DMzo+5/TP4Kglj1eSls1JPAEBM/utDCminUWAWQTLV
1wf//JUNxPB65AWe6tXr3cwJ0e0F4O22C1qRfbJUTz/eTgBHzrzqkQXqmie5Ydxp/Kuox9QLBUaz
j8SFl8uIW1kMb4d3HOka5vzJkZiplkt3xYMN2sbz1GXfa7hKHPeHe2bMRX/akL2lSsR3D3hWLg+f
o3BgdjDmcT3cphyrtDwZ7E2BpXA5M56rL89MhlVzrMetsY3HoK30/i7AVfAQp72yC+0GBBTIkES8
DOuJC+vOt09lhY7Bj9BKI7MeT513kZ+D6N+pHmFmJN9lisaHQha09DX0sgQ1TAVhN2LLOLtupzOM
lc0xArbCxKMs8h+k68VI6qnzjdYjd2zJIU61xa0SEN4mndZkcEZSRSIt86cDUm5umLZzLuURvyPT
jxPN4LR47BTT+Rj9A3SQ2F01Uk8HHmSIBmafdMfkjUP60zwIpgDb3UKkwWq3kIPqKd7b154RvduL
k0YQKBk/6tD9h2yo7daQcU3oy41iNHcP9cjBVVLWbZK8LeCx0UVDV9uL8ysGZpEVemdUb+JN8+G6
bLjxKSj4OXhPAhi1+Er1gzSWeo+So1GfYykxb79UTk0Awkdkzr5k4Du/7WNhk0R6DdPCoNeCrYcd
xPNk9rTAcqvDW+UPMUArr2Rjg/l/VW8pxN26wR2HBhfoJYIIu0XcLG1UBCDQTyYy9ugibseRdWib
qgKRHrbeIoy5d0/Sf2wCm8aNR+fm6h2yOvCtmLwZFM++Xwkhajw+zUkulVtHGQtjHDDNUiri48F4
yl2srdg+AeCGSRog/f+kasz1Fi66IwaSRTs+VZLU5hW74B0rlCmruAyllbDdv8vXNUYgK3nIAsRq
ZivGp6ZZ7DFP7JBBzcvf0qtDE6D2d1TAZ2BIHNTpILCFdfMZ3rJfIt0fdc4QmBWiSNnKfDI4wFFD
7lIkXSp1JS8EovpmnxGu+aCjft+XI/FOETULNlV8Wwr6B0nGpkYqBXH0EzS1DA1b1jWYWXJhXb6R
+VMtguvpSjCRFUm5f8oBomA+7NtIQsbLphbRww0AUYAvhPJUCa4xFkSoWa+Gcmjw64RZpkWTOSxG
jb07cjB0BE5cKBwoqH9kwcYx9KJnw33d4sRU1OV7zqRmk04W9Roa4mgKFqBUmJD1OHIKrVvG/Pxv
dQb6dDjvSpvMeMnZoJr3t6IIHqqWZRiDKtDsFaYmQiVck2h9MV8Xsyu6bIy0kfhBndXzhuKsj2+M
IdtsC5t17rq06nGmHSe9HajlnDv6eP7ozGnmJCzcx6wQ5JytfiZ0lHMu7zT8ngrF4XmngKAbSsCd
bXMjVC5tbYCb90XaM6POj+nkr5+umHg/sHmVSVdezBD9kmVNIomehKVvg1xuCTQJZe+Ijd0AR9vw
Y1Yz/rp/sLyZ8KUKbUtYGb4T4clTai4f4kziLkAXXLAefBxTlifRA0FGqP5Pgu3j+rHjrGvtKTav
mGPkX0kGIMWYeLJ7IZ597+mGgO/ti1XnYK0Ez2NNjVezMwd4BezQXaBNUYPmAASz2AQJ//2ZaVb3
MIdjrQ4+X/K3T2aMpV8uUOTF9HdRhxNc/4o50RXfloMxBkK046iHmXNDvECKnQJjwxgB+vXgAiBi
UlFDGlErbDTKift8MSGXKMTHFE02x7JyvCnVGVpA/QUrUHjHp83icPZDMyRTzdi5o2zPufvH5C2Z
nIhgFOo7qKfLiZ68CZ/YYh5/qAT5RY753D0RRsaLC6pNAAxD4RRAqQfClzRF7lZJ0wV0UWHlGwme
cga++IBwmvc05BMVeKR70AKgzkUJaXI2rDjyJiwXBDbd1YBiOEGKekJscIgT9ctDuJhBB3oPyzk8
FaiDF9bIUd3aCaVAfzIeumXQCtwrD66U54tPJdFBORv7t1b+jJw03k16CUx7zaCIx+v20VE6X6Yu
1BcF3pKJ+L8Sfw0wR7LheKj2UxleR71jQTThc+V8DYIHouAIn24+6T1tiIiWbuW6TOyiPkfvPGoX
xTMW/v0UbL3iJWLY6WABo2kovs21ZJXgTo3F4akgU2Ou4xhqbNg+VQLQyW1ZRh5Ksce4sRTZsMxK
CR/4T5Lbo7XqqBIos0Ccv7jDWudWIY3F4XFSCK35rhntrps1t2gS2QNLFpV6OQ336qM6XFWLnP8L
hvWOXaG3ZKIGbTvMvJVmP4rcE1OZGGRMmon4GPVZ/F4xygHGBPOZtMUQa4C9YY/CpzOjFjuOl6VF
VwD0AqR2HA50zWcd60X0U+6Nx5hwY2GpZ5H0q4lwQWwu+SoZ6GPGtYCeqqEmnR2Tk1pK7rgg1l6A
p/egtU/0rqQYXnuYhyDVOxLwpx+Ib4pNJZ4x04lReCltdp/bAOThgquDV2UG8LCDcTKsOdk3bH2L
DNw6KXey/2jubfYRn6udR1lElWIQDdcMyhFcKHEI7z7IP+UjTTDhB0EH75ihHdkojcEw6lmMizI8
zvwkjLIo10r7Kellt5c9Hcq9G6qjeOvMDzUEoTmAyisWI9rXUtE5Ih2yVdD1FXrPFRyTTuGUzlJa
RCZ9oQ9bf+0zaOn+RzdBGnc2dbYgxDqIMxqfgCLU64r4ND8cvTBLdJt7Clph2ciU0M/xZPNTBtn4
uG7Vv6KlLUcUj0xq+yc/tRnp+ISStUrMAJzsLFyARuzE4qSRwVifjfJgBmX1MOT8GA/buma6kbvy
P83rtDh1b0S87IbSqH1w9Wq0mf8sg21JBAqMaf4mTxi2OkKKoOEM5KRm8Mbxn4ra6PXq87KBeoUO
EyHAOh1INPHT0q0ZVGfc1CyH16yT2EJlV1FYefIU7FJOvEF4Dedx8De6jd3hXjiKHpGBDi5DKcIC
jJaRZsLswoRzAa0vGpEcFbHu+bdQO9JcsEHBwI13QutU0Rkbrdngebu/a+FZNavkof3zvCAywoJh
p1tH26XK0Iuf+P0W4pyjsOT5LMyFO+PalxzCDAo7Ydj8bNDNnvqD5JHVsbLnDCfKZuBxUijbsmYp
EkrSsGdU4P79Td6xZOE06WrBzxYRCZRqICitn/D6mWx6lznmyWO0tNpO58K39mwTd8X2lXnbj/F2
A0EkMAUEuR5Y+uXugfb2GuBFGhDmRGhTQ0J0D8IVRulmvP7YUjLohYMRgE5Cv/V90Zj+W2545kJZ
PkdC5Sq0kysPsIEofzg4KXKweTfDNG+vRIW2bdvi/HdO086VI5kzlbQBBujGHO3QUR/K5tB+F4bo
0xAXt6+UL2d8PcmyZjwRb5OOcj0UdnAMPtqeGUsWiyFO2GGvcXKl56IYKO8Q1HAlzfOZEFSc5uqS
TH07KN3ryUI23m0bQWxsmXpWez6qWfWINuwS/fweLUANBS2kYukQKzhKHFDf39s6WMTddLoE7fhq
V6I1d8hKd+uNsWQgZzmSD34icYQmvzyBk9y9xkFBMmUesYuIndKeyy36gpJNxCVn8P/sfa8m1XCT
wisv5xZkITsSlymuj6cWgg10yWZKFvhBRY4B1zt+M7MZpAzYp7OfSptBx38VynDADgPMOMR/xz+p
vmBRVnD285UWku1JM3DXOiCAqtYL4rfx2P47yiFyVIbCNazc6OXHj48IaKDvZS2A0rP67m1MyaIK
CUIdu2zR9g/78sLpQ3paXAw+5ip9uAfEGYCUwSZFgR3B1XMN5MZQKhWBfJVLBHuYgV8kHiCsW4ss
35PBWZlfrPBPaWcPR+J3IncS4YyTAmfNH8B5r4SwlIhB+wfWYpLAzvhaONB28DXwa2BVe/c0rrJo
rrKWCkIIbbZO8nvN8gCWjN8ZWXc3XldmnRcpD5PNIkl7SLBunq1j+SQcBeVNhBKUkPpg1B4FauYt
k3qa1VWfYzwLGmaWmxDtDtn3PYSGgCEgNvgciJZ1YZm95uFdqj1G44O22d7HnKy/LrL42CHRMvnp
JCAQVQ8GUt/njQfM6l2XiKGJpbEfASt+ihft3w5qL7PaUG8LRcyl4lDwCd+4YEoIn3Kp9rcuHZZN
wLnxAA/rkOsdKndK01W6OTN8ZndIWCV8AlHZF3aZzVJEr/coTMGcyvjn555MhU2gvUdODTDSqX3l
fOZesk0uq0O9BrOxnq7Tv+MgiIYGG4lSXMqlZYanqef5RsS9lA1iAtekkAjn3wvl8I27SZ9Gfn8c
emqtSiDirnwSl30YAaPNJJgd+9FqV45apygVMmi463MFuMCAeMxOC+esKifAuYw1P+f1nc7GzNaN
f7+9YGNQyrBKk1X4fH2st0CvPGnoWcHWXfbJOV0/LccebfT+YYbOOnq34FHKTrEJXHyTPWPBmMLR
zJNOrmPXhnR9NP+H+mZxD+AEJPA4YtZ+ZIFcfdyY0Frw7vFhq5iUSfhY/a6HOIA/Ay9rQT3rbl32
LxoFMGjxrAPV6Ygmf3WKUYXeZD7FvKW4AvPDsCPqK2VsuH5KyGbZ7meFUozQ4Jx1xv03jo/GfNnD
rsvcRv/Rb9XSL6C2S+3bKr4Lu58xx2XHEDnamq42GE1Qk9Wq1aj6A+aoKeDICenLWNnw8mAJwCDb
TeNxgDov2MEkIXxptCr15X1c8dkgNfLDWkhH37NYcxdURSy2PL4oJnHhVu98NESlCjEjpMgn6d38
phjgC9tmPKWTDka4bYEJG3ToqKG+KTH4b04L0gge7S425ZFDkWJZ/nFudW8ME5lkg4UEF9lw4X4l
UTxjT12kgRHKIbT5JE3A7XrVpRoemxHvL6Oo2RTGL/mqwI2hEMgRXrHwiIAzGEAry9HBJYdWb8ty
2mBPxvNWVUKZmFE2A7KLGp648zRmDDDaMQaX1MClvdqCZDwMs5/oFNYwLU9w5kS4sxHVwbQWD0pQ
GNC1LKPLbe0YAa9VRMyipxGGVfHgy/t6tFFECa/mNR7KrqIyNYKavX3MkXUddOCU6Hv9TGLZYtfp
H1Nc3X++mQi+2d6TPkAni3TKDTJ807PgClrFnfxx7ARPc5TYyHDU6arFuaVQ05tx9dW1DjEeRT2R
305fZakWTjbPrpg0DrvbVoeRb6wDPvWS3v3mjL4hNR7VLBBspsfFT9Nlg8McqP8bJVP+Z61ndxq/
QfT0i27BqOACYmahHhNnVrSaulVj43h3I/h/DdpFEsi+R+6yT+kLHG2xqIiUMV5N8M/BV3cJL9+W
00IIqchjGPiyHBVUiyZtIDK9qds8zyUlIgBm1kbkghCD4HvOf2KZSeNR2YLsjTIKtpEOOcOdrDiz
uztR+oEEIu5Upl9PTCQr+EkDGaGP7521SXH30FV7KN4A6OlaCNjhn1YUsA5t4GJsJ+gW6F2/Szu4
i01O2ulNIwX/LkK13riE7TJ4eUtK1+IztMdZOsmIwTik5iEBVecJlvfaLy60mp68FLsNvEbwy6nI
2P4CnIPhQ+CFJkX8eGgBHf0rmFwEVchtIoNv/tHOCu63m6CWmFH1g2MyFiqtPVgsx4QokDrIdLxN
gLl2ISsFLt2QIcR069kA08PyMtFHjDOvJloisl3aC+JcJl7DnMk9Q3q4EPFgjJ0/omXnhVf0gHbx
AbCwflE+q7N4E7pUwigCjU6iKC66qiZx3SZv5/5KTaX1uMBApg+7vx1/9uqhBrxXcE9YzrDddhio
4K2a2kjnKkI9lHl5+XHefVBnfeAvf+Ij8Owr6u09nYp6WN999DPQA1pVMgyQpX8i+4hfqm/EEPMz
Ry3nnzzr6XOHrYBEYC1h1WGWXoPBICBK3TNA3R629pz6MWACTjobEsZesiSt4rXfUp9GQaLlmY2b
Mkn4hpPMLLFgo5W4fCkMZJun4p7WRK8muDZgvEUmJbiTGHaEyeMH0WByDqzNPSnZCma92u9tZgLN
TL+UuXCer3Ng5rSuIWRsJZ85KXrnXDL5y6P7onUMhXN0Tub9bHBbDiy4PTVlSYxKwr0VlPqdhvFd
aTCXMRnF9eL5AaC61iNbtbXhIr+S6e9es0VRU5E1HASeLk2VsnTqlvDs+MyauXr4S61G2btK27ES
D37scFMcwb+jwRQ6c7Vb6n3DGPmA+mYPVgeMO5jznKRWmKdqzLes7o8dY8pucjBJF45Eu2awOspw
Yl5GzfKuEcNQs6LaXuG2TNLpFyyhecxesqifHGicZzkN9IvCmnL7Rr/i0GNYXJ+2J6REMcnvRHPf
j3TXr2Aabj5g83mJuuQkCIExcHbbtP9n33dlQOlV8PpT5qHeJEcfARIi/bUbNp+RoaB/q9vaGst7
v6EjdDI0bLD0oAGfYrJkGaD6YrO35NfV7M5YF2zyLNj1l0pvO4v6LpcvA5qODKFcEq9DzCFgfBwF
WWI7IOw34kYx/D9ySE11MRvsGTUFB6JZm0OXUxyHghXgZcRK+xurWhFn40sYuMkhr5IVJMYrf0vZ
9hSoEEBz+mnayosFwXWjc5qV30yRUy+HmAbII17Cv37zga2ZUkSFnv0SHJ/QsFET8xcGfXolA/Dn
MfGK3y1OGCa3Ze1kWxQUeldt5ii88zGq17GIeuwHA1GhMkq8CSXenRusPv7zvCri/B4xh82ZO/eo
MB5Sis0ZW4wvddFCn+wzIwoZed4t4ByE8ZEHH3K9NV+mWyfeY3lz7emgLcZRTzjdAmYrnCbpZ96h
anPAC9OVN078kpenyO74abqlHvOTdFdgmP2hkBk6RlwMFXm7am/EZGH4aVJXFlL/DqEN7IUBOHIA
MFab5XFrOayHyNlql0sREiTnklB2Pe/ISYPMtAQFFeHcarjNZ71UAX+YSBhS5bu+hzILs9GhpQbi
RZhQTTC8o5zTxCKmxl6Ye51A0LgOM4z2vn47Fiuqu+7V7X+X5EFuihre7OyMSfTSwnkRV9gJjdCG
rPOXSLcx6ZUsGAKdBgu871W+mVxzqja/zc6Hl3PQJ+/WC9ymMFv78lyvnOa/yW03JXKpaq+jjISp
TOMGJnlpWwANmSyrK6FNb3td+AWdC63jmrAunHC9XwKuCKxuRZgKTmMQtP+urm/uybk8f4oQ/GHX
mdeDqS0lMmNoon/OikLmCYifl8oLI5rflmHFsnNmgTAD2Ijmyt0XmB8QW6T/hpLh6zGENEDmc6wi
ORMusLlc1rjuenYXCdCRj2dLV+QFjsEtOTjZW1ZjdkL+YWiuoXI9vUweJgPAuXpffbXBWnAV0Mul
nhcgxJHCFFAvZ+iXYD5DAGsDr3JwtjxWAJJbj9T90BGisI/YALnCvZaArOvzVJTeKfRd6EhAlCBP
jHC9PzE4y/AtYZrcb14N1ZiOJJLahGkoC90zVQGbIXfj7OP1bQqwcwI0fdQls15wj35THouN7FmX
3RxgwRBuWFkTkAfx6DfAXqnbpUbIBZqHy8AkxHANAZYpaZJ5mkdReM/ehpuvH2O56X3+3FEVxl0f
C8JSgyEYhmpiVIs3iKJ5g4b9N/ywmoNCrSW60srC6WbpLTIpQwY9tcqyJ5ZPtZuFbk2EHh8ovV4E
GD+drYk1lN8fqRqZ+zUdODyh+T+6uBubo0sop8zHfIHlAXB/+JOq48GUwRjXhemaWuZTLpVPvggA
rc/BDYD42kIUbEdkW8eKTl8UrkdqIux3smA3PBP8wvvQUtEIOYQlEvrMHwCmmUqWp2NYA1YWiTa7
srqd1YOEBwmMS4fnn0243aVBL3i7p/y6teBk3503F/mBJ/LXqGMEcnOugM9zeWmxytDcp4DD1BP8
Moj7cjVbWJ6qCwR4a0m8zRrlnyOJZEUoxWF7MDxjZb7+zIdczuS5fBRMPE9glvWE7QDNwe3K9OxJ
PFGDbhzPGJ82lHsyAvyukMOWpefOQ+ptDUYzs8y+tByhJuLBklLgw7GYRCsJtzdr5MBouMano0zu
7i7WBoxeyk5pQj2i/Zpiv7MJnQkYiHSyIw46SjfmaJlaWhqNownlk5Owg0mPhJm3xCpeOv6+zIP5
vncTYlzOuUG5YNFe3YmzeU2fTOCBWsMKB+MoRegUBYAk2lStU53Q9MJPBLFOdCgFCCdIXotV2vAM
qvPGZPHTFN02RstcHYIcILlVM04nvVxnQxsQG6igQP+pqiYjDfc+qPDxfnFzGE1uPqBEZTO6gjhm
Lq3JXErHIkUg7pbpsJvxiQvf83wPHh97MAIwc81mrn4vzUKcrzWZX869YT5WjyqOwIceBigbg8CU
7ZwgrD9TC7GARYeJ2wxjp+3CwoG8La0Xgms+Cj/7LqOUzj1akK8wxrEmbB9j1WdfUQ78DV/hZR7o
65PzFAc78x9coXjnRb9NXjXfMy5+KyQzK3PQxndLCnZ387ELmg3RJDEEqoaaS0G9AnVZsJf1x8uX
RjE9QIR0RvWSitkTh1LsEQDyezvjGvY8w8jV7tMC+3Rq1lbAitPjSuoH799gBF9q6K9Hlie5OxbM
9GAtCV6nwpIC7be/1Scb0zJe4CcuHQaCnosYsOlErLGoPel2bft/TOF4+6KPtz1XN8LveO1zoQOk
ycUll4TeULpLybZ2fftloY/RFnkVABnX1Lr4+kilmfq+s8LKlD2dE/Ca35S7bkvKLD2b0qdxR6Qe
7xAQc9+/OmAfXB5Aydkw+IwlYAhpEt7MJq487q7vQkUG+sPDDzOKJPZ8C90SlgnBB651HK8xHE+q
FOvKKnLdvLW8bnbA5nOXKAkuxjcNhq3aDRKJRuopSC0ZKH/+p4kaMgqaXIL1VT7IKpxYeQEjVZq1
eiZXNO3hrG2aky7YixJpc7iTtmmhVEJmBPtSk4dhAjow9zr5CQOihDq18R+8z2lXWxcKg/40qv1M
9+1YwU9K01JOdrRtIp5wvSRdwtGSy2uwrkwNhDiGvm25y2idX+xcpQi1o2Nl6OROlsoKt3X3RYPr
O3u1Hq9AqCaoCtwLeLTL+GAjvV9zUg3aImToPRNsAWUbUODgFzGrczhBIuLDOqg6fQt0+yoKFrwS
hC1vi4NR+V4xFj8AKmM8HbGZ+PY7k4Hytd19gxSMMVtmLaW6ozptJpIQn9frLuVPND0WhdOivX3T
0xYZkjVdhzp7qxnGUWOGwEVoqQI7X/1ymkr8qo+MrKhXMWCNPNqnydoUM3sQi7YylRpoeTKLD7OC
/kqhZV8SOU8ByVUVRllTKONFGJdXiM1rHUT8OsFfK7r19At8ticNKOAtLkPc/eXpaRT1ZNrX3mur
ThCT8vLKaM0HACsfkI+5r3iHKJ5EulRlbWZHRQDVQ9s5fVY8vRtyJyrJkhF3qZMH8UzadYNYw3sZ
2QHMVZko5Ht3qo03XdPAaWwI8kLMQUju6BmkPWKgYJ2qeSmMu7QI/SDqyuUcayNohSGRUxAc3eHJ
FPHNYfbhUQbV9yKAuT91iBy1AMivjEgvcPEoa86gF91Wwm7elb/DSCVMsd6T/wb5L+Ctg5qXHMFz
C5WpXI2SNPjfUHHVAYnh5HxLkw8qkmDrGlKxexc5sEobmpmymiIHnvzlejRCy+S2A9nWXm52WjD/
kEsGnGOMSNXeBEFKK/R90U4MGLo3B/CPSK1XxBr9wGWCRd8PGdqjOEVmYroUf+78B4BOqBVOdEcM
Q3LlLbnc2zcaftlpIG8xjI4RMBEbvieKm2++eoWzpdvARYNelaJ5/B8ek1jibdGQucdIb415kwPt
gGKcp3uksGXZhUgyBwXqKtgs1eFuHGEibANb8tTqrgzvuz7xBaUfHvo596g6WkNXJC4BZWzRAa29
YilHa1IOdGHFguLHpiLUyo/X95FHy9k71C4MlfGE9k1AbkpcbqMjY8885aqpDtXpeQMFyCtgYkCu
2a0JuZuqLUz0XmewcjyTbKi/xf0fxd0UG9DYNdkIhn+9tb42fEURqro9+Hzjd6GFb/vopUQa9nXK
P/6aGINgSFYroR3jm+SO8gG6g1QGmCxpfMQViqPVHnrNpPOIkqpOX33sqX4aJB3X5uTNRNJUspft
1QvQC4L+fUHMie7J3U1rOXiwriZsnTflH32iicP9OquDiJ4+85oA6eI8Fkfx4Kj8JUn4Ny2pWU0e
pwI3t353Dhar+oDB+ri3PSeAXd7RGnBIAYHqO1iO6K+TUiUV1DRS26rjdOBB+tYVVtyWFTvX992+
RuO/olc7pedmvh84vC+yDxM8pOpDnI5HjgOal+rSKYt9sixKqYoznJ7hUX5Pgsz0F6/Ie6tRtbEl
1umvWw920lQJLdx8gpLGX+gvaArD/Pvh8D+mSs47UGwizNcnGUbwhEZ9g0/G1hIY2crdslJmtqY+
xoThm2BIy7Idiyuu9pL2BjPezwn7nJ5K4s4npgiuM3eiHHbOhSmbZdTsuWzJMolZtgl5bw8BOQhU
vltp/Jr57+huczwj8+xe/G952AGNl8M+nmcNnvRZDchYk3tw8dbZjT10oNeqhwnyqZdrP8pIajg5
Dy0/3O8MGedrR6jPKDGk+fDCKlfL8ZZsOkw+MtS5ltJ+WL2AspAPurdstUfz7388PFgItPlMysya
3EzgaGM3FzO7wZQSb6DhRR+rXAIqASflEl/hGxkcgyymgf7SLri6oltaj3sq5Hi57CgBdvA2VoA3
xCSJulhBdVruQV+eURkkNg/NxZX4yfI9nk2uv3UKD0RDgHngozK1KLLnBzvwq/sVsopoWA1JwIiY
wTDtwUHG0OGa9ALDAVPSlErCrI64P8kUn8542C28ESHuoPj1YNPmwcn9U01gOeX+i21VbnIOm8ll
HjW1GBHW4Fvdhvr7z6ePb1lNFXOovZEXghU/OQyzGnVFq1eTZC8kNGpA5nCdlHXP/vuR2Ph1aCcj
ciBokfo+ZVP/XBZIUuGqN1C5To5KiCzRF3MeKtxkgx6U5obWxwXVt2xBaiVvZBP6OkpJc7dyg3ZY
oJ+BTDN1tyfL24rRugXfOK7HckT73uBsdEvQ6z9lxsGVFIuLWLzjLZEqQN07jns4wj4xIF4P/NGZ
w+Vt58KcAolGNuGP9NfUxQmKhOpqOC/iu7NVwuj5M2v2WZgHQxneIVTDSh7O61k8QVGpF3aFwP9A
q99s6yNLsZSwjm88Q7Jwrcr9197WW1kZ4xanySGYey0qladiclO0/WtV95noIuucDCNFueF76zAf
zjaFtk4auWEDP2RpcqYddqL6vTc1isqo31lP+Y0x54Sv2dBZ3DfVJy2t1RzZgDyyO+6O+JcLSiDJ
lb/WotbDo4ugAv8zb77r5iyUsbVfF7KgOL+bB8G9fumyfxP4VExn+TwL5jvvoxVuQwslyf2HsRSu
SmHlpUs6JiiaGzXS3WUuuEbD+mjd6FTHxZzNJWqMaRwMWzZZt+b9k3BFf4X7LUTONwn9Dsh2yujB
e52U45FZK8pFp/p5qBKAralIclLMjZxoWXVKrojMWr4BKHAEWSg+RsqdCWS2WdTlPGtzDEUDEJUe
40gaT3FQ+ChRQRfhGyBw6AEVAfDvdWbyX4wPmMn/flNA7vfrvyqyws02V6JG9jnQ17EJWNoU0mNG
ZvEAUoza4ihrPbABz84FEDic25eVASHztgBmLuHTNfDJ2esvEDlnVIcMy22Bp4hKFUikgAoCJBT5
sxIRnO0TxMosvpVw9SYge901SaEx07hyNjc5RBPpbLODn9XWniDUnkkrvwrHlK6WSpN0bTaGNf19
UbmW44lHOuevWVlsDko5bASSMW0N61/wHJ6fuP1xOHXIm4uv4Hl7aKUkzFbsOfpvqcIeECGa/ai5
Yb1MPpfeYivaILpZmMCOsDGnh+EbzKY0+lieRG4OwklkZ3wi4yPWcG4V2fnWy1CQXp8ptyg5xu9B
Sw3vq22C/mj9lSytF6DhTaLLhzpQLjJ76MmqzH73jZ1iS9ZYaoRH72UtYprZ7rK1/HEL2gSedKyt
rCBeRGKkJJ77qPF38fuEFZHnQIUcPkclkc5zU5w7CTQ705AGy+Ss5QA3ykQ3s0ByPslOlREhs9BN
gQnQkkYzjD4dr0ZmwXDQ49rwLrlBv1+xA2WPHi6qnP4ZVSTBryhscZ4qos7Iu+1OroYNcR8ebop9
uc6JAZ2rvEOE90z3p/neG72UCpnDyxF70PPWPhYpJeLiYDCiD1OKVaYmxeX/ccKvzWqiTNcmdf7r
4BavEj1STUriuYRBPkKmMeLGnMAvcFmaSaa+wbdCiIE+PyqrWVrCMwYv+KpzkjaesE99DnpvFXKq
qYNQDzZurXfMwf/QTHb2Ioo3T/gXsAZaM0sUjtLFJWDR3OlHIvNg1mhdMMsyKb8YB6QLuW3nD+Ag
+sCaqN7MjVwmKEGPWJc5LADrfx+XMLO8gSZ+r2PGcx08UgfvBbQpM8e0xMGbKUxi4clf+Lw55bhl
Y2lWs+VNJkS9oxmE4M+rVg+O87RhQkNLn3e9G+/zrerwUAuM19+wMq285d900EJLFfolMQCd7bRj
3eEd+6uA6G4kduB9VBuKQ1rJZSNgtvo4KPpgxOHJBh6fdbkS7sfQZoS//ev/T886VeXWBuXtYysV
JphCflGsGO2Hl3v/b/EgjRDvV06zXXCZMc4M+GBGGrnyEXT06OVxE2xDbvVR9QdtC6YPby7J1ESg
m9QnaQFQS+kdwg1AA8L4Ae3lHfN4ZFnSZkw29PxpFwCuRJKRb69qzLwniC9TYMGLu8Wxp7UkNQsC
hYxRL80+KefdjHi+AH2624HJzgD6WuTwJwTYEHUsLhOfQ4Nwaw+yT19YHIiAVVsjDvFOMwSlwkz1
bR+QruYeaPVfN06E1fdL8L0/mYC7AYmDKTricL5JIsV4w2RiwxznGhLBrRqBSGoc9ytUo2qcIgmh
R0W40hxj6/dq1wtkqQDOOwJvRR46oSkzeZpM2s6BNpXhHNBxjNFBOqADSuvHsUGo1hC8CX1jzvL5
LzMep2dySQzAtmrmjpRfdPCbkgyo1mJOnrlPVW8Jl9RZH5X6b2Qyq04r8he/RvHk9DG3NqmrDXjK
S6oJoKu/cJ92+hQCPZolLOPr4DwL1KTi4wV3Du9LhZg1UVs8F1QFl2PMQO8vRDYDVMnhFs3+PhaL
s5wUhqq3F/DWqUU4i4g1lC4dTWTQncOc9rBuybadqkZZg33cadUcLzECfcB0VBBWYecG0U+CcecV
fed+/KcN6VmzMjGZd0pahkWPq8FabUxSQmjfIynLexuz4/PKRkxHdluiCqRMl8o2BEN63eBAh/KR
jNOftjDTWEUFCopioMlrV6Idq78VYb6sAUujNTVD3ArCAWuzqIjn1urc/7PoGtjhb3Ypn2cN5771
AOaqb9lRRm22iTbn543hMTxtVvwxEqz+XcbcAHZghIlUPG2iLM7WS14v60ufD7tWH56V1cP2TvWD
Uh0krT1vkXKGjVNxr4lZqCM7/t3Rcsxtz5JWXjiBxIuRrMphKuKVLBT0iQsuCJvljpve22T0nW1u
JOHr/qhAmXNESAr61CAj9RA7fS4QewP7EaLAZJ+IRJyGPDY9nVl8XWOuqIIK8ZdZCNiM/j3vQ+Ot
84T/2ozTWxucPffR1MFCPAVhvZzJAuTmI7+hHIAk6rco3yDEdi53RYD+hRkzS9BRkhc5B93ObPLZ
6+/SHLyEQntHge/mK6PbJ5ETdErtXye6msDNNAfxC9x8tYqTgJEv/L+0gctfAbkDYca6S+sIp1yD
J4qOD+T81kKyVTslMDWaXRpdilmhz41yQZxpf0hvSV6aIXuWaHaWcncE7PwARRsLFtU+qxoZqF9s
mKi/2BBygUjr8BkMP7gUxMkaQ+e+vU+vvxnWQ93MoLpXxy1dYvJuJ1F7eFzs++YV5XgNY98exQx9
fwwLjz+IzQlJLbbm0Z4626PruN560ZDOds9nbylcXLuUte7mig5XUoDJIqVRErHWpcqYEHUzUe/H
S1s9MuXc975KIYSR+3ockAi4GL11ALtRePU51yj22vXqh4pJgyKuUTNcLwyioimeF8N0a2snUOZk
vW74z3gaKxRqgPVDPuIDB0St6QGrEVBrGYXesJJ+PGuSAGWGp5sDeSBsZy2Aqp8saFkUpc8pgX5w
s4sVCz/Rwdn4LMLzw8xzAKGCelUurdQoyXemDncaNjysCauEeAlYhc8eNM5GdDmikpLUvkbyidNm
ou75b1x1L1UE2xbhs9kJ1tgu9ja2OjIyd7hSatxgiwTFdEZylrQGD0hPRY3zXXhaziiYQEaCYT+9
rFD4EjV842unVi8shwCIaVG7ePRI/xSJ4ZLexqNZAbY1Nukq0pDkGMfLpVNwzzvP+Kr26X9X1hm5
Msiko6nzcCNFi2CvEciViSi2ilk6VGh5nD29lKiZzniJcBbTr5NhMR2o9RResmoWBJTxzuagFceV
vTjRli2Ytv/9N87IEiXMdAnMT1SpmFCt2HU7J88DHZs3iXiJzb7G9GMVI75k9m8q70XWAtxhMdyI
2ro3WQPRAqLqhJiA0sV2mnVmIY+f4CRmUmflRaaoTNXW+G/V/jAD6thBo4KuAJ9vEGdz7q8qohfu
hBpgegKwszTJQ/4e9R4R4+Z3CiYE1LVpFUZQJJ5vjjZF0WcT6txGHW224nrHLm7vUIBzqz37kwMg
7cgxJEPLYl4l8tpr1MmRhJ/EoWsfS1ODILSdrNk0OAAELQXLpVg3aGLgXcT7ojarc5tkI7wkt+sm
wJkvEAe/6/inZ72EFe92Q4ekUIf2UdNsk5B1Kdp2Ro2BwvMLQz0qY3iKBKFmEQ8oFWj3/RlcH1Nu
QEXHSDgalHQHTXfkZ31hZaIotUhBTJWGToG3dNG6xdaIYZz87BPbYkoS38sFjAjv2JmhfPtfQk4P
aLJ/K8yKdo+3m/KkgaxXn/MJjSe5p23GN+7vrxYBc4My3q9eK1m1HrLuHY07vkAIlOif74hU0het
eExA2EDfz6hq5EphlkATgKfxEvI54+uOx47ndwdX78qn1WjAPmPYdihBDBn83Rbzi/PqDDXiGYTA
4lJdn/sjT1429MWe+G2kH198LU4hLLEQSziNC+SwO2VZhmjJ/EBmqTwcnUIDoO2uW5dTOd10OHTg
A74Ax8eG129XnDB4cxcZvxRROlA5SJ/dDFokjqy/vWtULCr7leSDS+72u0emT8vMyOfuVZgvbwRM
+h/4vuvCDx8NkvxNrhSEW9sP7GVlrVgyteeI7jOhH8XvR2K9YP/6+mjgBEqEWIsC1PyT7Q0GWzL/
VsHO8cqS7w1h6RfdsOGCQjswweAJZh5QUMnAsCYGPLsixnn+FH+ewjpHXvo5kM8ZJC+v3RbRwY+r
Nos9KJ11UqnYf5zyv1rJhSaWouFa54vQjSB0WYpsih8dbVkrOul6Anfe1FQEbF7Gvt3rQ5L+OjvS
CtgYmdRszeg4/il6kVCL1Vo840KINUc45yftpVhiyIkZc5r+PQse+O+1Yvr26/L/7yOD/4DUEMSv
SH3MAD25Ldn8pEapwp3bfzvfiZwTtLF6I85rDkB2/FmlN39g6Sde0Cyt5R0ePhrRMNKr2C4R+VWg
AWEgFsngKsigM5YnoEXg4EBoI7U4fa9iPmqn1YQfugxdvQR3/CHGxo9h0P+hlZdZnoH/s4AnHk2c
/htd6uDW/U0LKEHS82T2PKTccgwwzPChBRqpKHMOAXv8q0uGcyZ2wuWRZivO7algTdn4yh8J16HI
CYNPs1bB7gcwIyolhXASe91HuEynrGGQ77u39/eM7VTcu9yOTbRcNYxA55/iLCja4GhHBOy6Vqlh
VEXgNE0jZi5kYedrlu9szzbQE+WTQsiHPZjjtcz8KKaFGn760yfsP3wol4KCDS7gaFLbPMaLj/7y
956ZgavG83WUi0BUIXtF5AqSwsEUXc3EAP/l34zgr7qXxJwU/sudaWn+nVreAZI79WfEeL66V9NO
auL4coNzZ3RAkkew/kA6wrUwIGOxGuwpPFe6cTYPvoZyeAEZoESIEetRIIn+bdjivonYl/Rip/xM
OETmh3z0dhAoLXMCVqoU/j9VDlBfyCJixf5QDqx9BCpeiM+IzovDkdd1XYXSAa2aW6Z3w+EkcmRQ
QhlrkOiAIvahuCrrQZ3pdfM5ltWCzcIadZ4RKssMBYRhmxzGDi590wCA2Vdf0fUirhjIxdg+UPdK
g9phSMukWBkZeFGMoovRzg17D2CC8fMuGM0LNYMau7lJuSsGN03aMSZmhw9zLS9TQUHBOGjIyh5M
OHTsxLnZyN6exiVoOk97i4kRRi7/KpectZGLK2TxQLBTBfty1DLb01FnxzpwlpeWLqXZzA17Tinv
7HLBy26scH8+94K0V5a4qaJjShNU8j4afn27gE40MmJHz4SuZ4gFHxOoqYN7WAWSbV9XkKketgQR
Kzwbj1fOgFv401BoUIGYbHGhq2YtVzsNFl3te27s5vBIjb6q5XJYLxOjEmEVuaBmf7guYpAoeiPH
MB2058vY+CkVbqZ3IHJhWuD2hbl02U5FNMyYTg8ysH7N/5Z+Vp6oeblnhyZ84riZY/E7yGUEZMbt
EH3i9ooWOp4qGRdkZUN9GUXOXYdtsiI1afiZdXSqzSoC33XRKMdNY8I6/sAPzZijHxDgW6lAnaF0
n0Zhriq/cv0qZu+GAW/KVHu0vaRwY/+nJq7ybXbKE2Wk+xAEe+WVWa+JYRAM2yuPsm86DpWAzw9H
urT9ZqEBenFQhIcaPehmgUJQRpS93xQMquyNvb0/+EdcDq9a1cCQYXRUbmvryQR6s764f2U5jKe8
WienK8h/6F9KiBWPFiiTbbzDXhDJQgv6ZBioTA9On1jZtjB6H6bc786xVMYASJdFe6TQ2W3ENHyd
Zly2mcUvXlA86RtcE9Hh9wMf1Vhd8yQaMea+yuQdZLeM9jPdg5HOl+TClg26KLW7mfBu6VOHLnXW
EFCC9Py9KN8mHXBETwTBefYD3AyoLjEOJ6Ltv2y5uYlyWPzt1Jgi7fHOyLa1d0gpFbhGVaCdmQg5
3D4T86yeAgT2ihridrUNCsqwylb0ddBYwq8/PsmuWk/jnoJXtETl7KqQ48DQNBqjW2Kv7NT6AQRn
J4Z59nlnpCcikWYR5xaj4W8O0z5QHDjRkPv5EwcggzwHRKBJlm0Nn66EaJpyugXteuqitmj0CSr2
8TsL6oBy2sKZtudoYs9GtsGarVCtCK/r3j5xj4GzVVN15olr1r4oHe8e2nPmyEGyE2dyUT79Zkx9
TyajEvS+mzLp3Q0RPySe7v3VkNqoaYGtR1bqxs4y9lTq+83CbLo5q5aMdjg4dNaXjMJ3enYsabcJ
WZKwuz50ERLSSAiKFHwpCT4sIlzK/zo2Wmlt/8Pnnei3kraufJSKnXo8o/gbN9eApwzvuVkBtKOG
RLaghkuEf6BipyAIZkEFBdD/ZgkRQvZ8F+7UdgcGfsg6K2vjAfKWI2FD0hhsE/8n7JLXlszUWSnP
OcQrqWaG3RjPJK34/Q+o8FI6exymSmhTfrsfn/GP2SecSxA0bJkw3geJ+s+YQJ6OT5ZQ4CuRku5r
MOtHMN7I57MKKluEoDYwkK8XqT0XddGIsaIhOdtqPc52aR084/sBCZQtZ9ke+RiM3eo2EZq4aDh6
B1Lkks2KsslSqHKPemG1Y17e31Rd3RyDxfnixHSVq01qTwPqJyulcWT9lV5W4G8HcCopnkbUYeWU
1CY4U2Eiqfx8x9cBwosOsNvNeNunxTlMIGE27J4X58hu6pVDRnrDYpnlYIrlXeCqNK9+y2f6tS5F
32zMx8AcarIGNNSWu/9LSKu/f9e8sSVZ9A6eBkn1zRCAguBDdB0ezbNQgO68CDdzp6Hp9s16S2f7
agJBti7omywDIJdn/H1FP3+3zj6zfh7rnV1VQknAEnrEaIETT2gfmbRc8s8LZQftuH8L63Y2eD/9
lx+fIsTvl5GyN4G0RZw9FLFMKDheU7icvimEZmrhE+BQ9ncKwUn+G1Cm98kna8Heg/TqsvxkrpnR
My9x0AIZ3ca8jIsuLO0dFb928vkM+7k/HFEnxgkBDlXCBYQQJsuuk5hDFvGRVtj2GsStL58/WwnV
H47J6muE1HgmdhaZmm2dUmhysJDvDOEBtUMnNi/5BKOJZkPMJrpq5mcRn9UekN64aPvN65cu0++S
Ebak3ILEDOrf3pasQGdPn3J3VQmJmB4ETXtnATTXkR3w0PrPu1EKtn1smafcZAlDHs6B3GVCs4V5
rxwk5AE5mwor1twAHhYqiShnSiZ5w1i09rJ58XIXRQEiUPeIuxwX9R8N2CVchTRMF93azBET9rrm
6KyD0ulbvFGpuMq3frPT7XjzmlUcljKz1FO97GRT4zj32KF0Xw5VvCkbP9nueLXGTnafuZJsHkII
BUhppKQb1QQFzZea+FiVK6n/jlObmcPaoyPdvu67BkfQeO3NgFRLPl6+3L4W7kmGDdMdgXitk5NJ
50znzF+2kCj/8tlNS0m7QAZRQ8RKpOSZTJ4t3eXQp3dxNa6Umdz94MkYHiiWRsqGuL9wZroAapn+
znoOt1uST2g4D2DJcZ6saA6dk3O+iGdxb6bSuS6oQmVPjtGHmFtPbKZ02kdY6CxtvU55t5NUs1Bc
OkE6nA5W9D7BUs/eGfvqUjjS3KnqZ3L9+kE+uKVN2/+wGWro8hTGk7IuuCSMDyHHDqCyprrJFkHB
0AE+XSmdrsQFyrcoiFuBvyXyWsQXwZ8BYnODw4FPNBkuI0WBhgdMOcfzHVSJmcHF+AroNerhXczO
u4UTUEwxQw3+eTZPMwQMqgai4z85Yw5A87zSDtrZDSu4C6MOjYJQNYYJt+25R/FzPynM5GoIIikc
TCNz7gqS+plgd8/Dwl1TjevlrHbOeu/2dRcM1DzS8KcEUfnhsiPyqz17mysBue3KmSTKVSQcDanl
pDDr4PGOjtKWxZOh6DlXdmr+91FGjjzzpG/uBLwJLEPdOk4h+ygj2stgM+io6TUa4vO74Fv478Rg
UfOfXFjlRB5z5FgDgTfsVTl0SEeh+aQ87+U0r9bRgisV4zz2PDCDBjdpTFGvKm7ThOrUL4QzLj32
tQbDmRebKOJ6WvII+bLhSXOPVqhm2fYeasJpYols8JtxAKst1QZ1rUJDsZL6XTal7IDXuvYqHlTy
A/2WeHb5oja95TM4ij6lqaM5TNaCAKv0WuIJ3ohwBiCAM/lWPyxHQoM8Qi0t8NRIlpVA4IBt0RNg
YmRFyDp67MSRJ18ubmGxklaGZUBpZ0S5T8jfWoKK8kEwJX/109BVcrwp6DQI+trMGTe+hj4N5oAc
qaPzTvYCXoOEtuM5g/aLWpnsVeIbUqqxxJpx6sk8vqkaXbHjGYMpmlKpQyi7UHX7M6DXw73mv8ip
mewIsF2iX57KmZb2kfN1XnxvTbrbwqdB+k1v/0Wh1zlfRqFACPclnqFV5amxdTnY8cU8yxUWFlhA
Y1yRfjr35yYceWw0KVMCzTKG2ZC74JVaA03hkn0Dr+ZU+L4mK0LYhwNWGccuz0WMFUlR0LOO+IFg
UyrFQP/znuU4jVMEvm0QOgbtwzWgCCCEZWYRuremOb0/VsXaS8V3IC+bGO3YicfX3yTB7+PKzYki
VOCyJhwQyroT4Ut6R/Y3ricFDriLXKivoEWDXJ5MQKFOOmMiYltb99LU2OQCc06pAWvNN3QUTFXY
+Om9NvlvgXp29Et1FYPI8Cqz7K5K+Y6GninnRMJRom580qWHdCOqYLIe5D1STaidK3+ZmZwUlp+v
6P4wr1q+750KkGSH89VAfHnpQWSnKQWpTnAb/5+TFwtBhf5ZsXH892D18GLQRQkPA+mH6PO6h+OZ
YVkOzPF71dLY6PITiPGjpvbR5KvP0E5/vKQNm5+G/GDCpbq62aaE9Q00JUsdABUQxdb8wfYlW6tW
C6AIjhiBH0bXiyHj5LDJDN9K278kw/U7K+cpHeJRfl6ci/c87SVYyd2/ZwjD67cz1uU6Drf6Zuqu
OWiUzJYnvXjyR+E05So1drqBW6Ge0U8aglJcNjqo0LrSs3cowmrx7bvpMkzik+DdhPOCEZfzO0EY
owWmc0Rm5EH34cYY3vrg47em7WkSP/7YBMfg8oErbi/4RAWO+ciD15yXycA7bcj39iKwd8Uc3brL
ICPcWqng0eV/TVVairFVjsKV6Xxc3Xgc3vuyd0GfV5MIE6Z6A/miakaMLTHl43iabJjhhsvHoeH8
beBBktDUKa1dX1j15kIAETYKAyumFVp665+ZDmBMaOF/292/iOzwtHwuWmwuqb3tJ3R1xGSqZniX
oppj5KdHCho7ipAA5yiii4vlzRjuhfA+iPH0YFFxNHAolV2yUCHi8A5vMe5PyrSP2JLwAVSjVD2v
flfP5vPi6f0kHPZPvRKj+Wjyl1jcwDDcrC1M9rdYivEaDSA782XGpYe8eueOgYDnmqFnwNCw/A0L
Ic/98UTQanrErCHTp6dSPWEE50QQoE3iJdS1G85oeu3YCAPBRlJW7kE9j5P8d4P9aFW5FbLU+4TO
UCSLHYxbT5/Bx6AikvAj2eP8CkHXYth0e6xSM8e+NiB2ByExyhjZ/GuRYjJNzCOTTCB1GUN7XsiA
eTDeYTMXSx1HljAcsy8ncJo8H+zvJn5jdmLUlUPzC7ZHK09owqfnkfF/qhXhw0jP1VBZe6sGgesg
ViTRISRf1iMRCAjG5znCOUdL5SNp6V1VpzEEiJj5/D7b/0WxOtL9wWtpPQRX/wwl4HEMQjdSLjHy
J/B1aAmG0fkh487Rawy2m6nyWZxSfpApUr7R9o2T9bHM56Jle+OYCQkdsn9xW9d6J/1Q1vxOHUaU
WEjuR8+kXJTgacWyAfIaO0bYB0pZmm3PmDITQLRDh+gj9LNa26L0xu5ASflNjlNb403QrCB9hMhU
wLEDQuWKPVUF610QfshqiYvj7kmVU8h6dBbEfPFrspXVjh1JUmlBPt7t85v77l8VjVdveJTTdhHh
jCUQkC7F+ty+U0bq+roIKeMyuWzZowM96BS/Jm7GmQTzeMpeQM4MVZ9wIOF+Vy/pIGJnm9lW/uLz
mwEu93dwpQDhS3YrS46jZHPw8JqPblq0INaV66PdDFfxpWyRL+hFLghYTMH5EFo2CtYZAlU4VbuE
JrWbIYVwthYA6xhcJmlBhjjnRLjPIcYey9QLTFpSyjMblhlc7CrCoagsmwCoo74190ZOgPmA96Uq
6+lDm1iJJPraEmHNSg5VCDn76QFDTwV9+X7f/27NN1U8KKeIXsmWbNFd/DYTFdwM1I6T6IM+WcQJ
+LjRJIjmUGzYpgMzqAz9w0pLd+qj2VhzGp5Z1UYgTGGVPToZTMku2XGnBKgdDQlz0M2piMV5CqrU
0cg27uqFE56bI+BHjZpko05BW5wEskgsAIQObX9Cu/AW11242Dy8Ekn9Z1bvNYNYy1gvnOhg47c/
0d/m+3pG1Sh34ND1TJhDdbd5my1Cwbpl8/jVgbqmffKJVoTYQRh2q5J1E77jK/mO9eDVBOuuVcqy
23is4RhmEUj8xEl4hW7A4UntleffV5iNxY/OR2hnPsNo0JiEePnea2yJQC1AuF/+Fz1NbO9tvjt5
jIK4oH/W3wVL0ABsJy75I1GskSUjJID52Marh7OXynpzKuGALiFQqrTdLj6jiXZyslVyquRcApyB
azYWBPus+4m/FQ9Jjyg2SNvgARR3XM8YNKcxlgBuOuTxi7ilJdWxys6Vw3oWlgg8exinHX247XwX
GiPJgKgty+/IqpM6T3cj8hSDKXI/8Y3Wyc5FG7zwnnhaQEUX/NtpkjT6L9D2kPH+18tY2U/JFWNA
Y3CHkBOty5horQQ1QxoQ7Ing1ekWPe0YdC9OcKDrovKpswA1FtglJ+OhpY1n4GDAamuIKdVDsabl
RM3xz+CCSOJ/j2qIVcR9Z277PDc7YSZDV3ImtjHL5jZ/Y7spLyjAZPyAD2vzpYYDQAiIu4a3X3lM
ZgzO5kipiqb6wkFbPu+gYHyEQDVWHL0YD8nNaKld6bxHaRtC/dIjqSrIdgdmBlIyNMxPMJhVsnNy
UaqqIZw/+gVCsSSwEEMIdVu4u8NGacZc58lLvquUCpnUz8l3+NYz7cPG3Z4yisAbQCtCPgIgdXa1
7tQg8BskrwsAguGVuJHXitVaPFSfNGpvuNjITHjIMzab3x5Yq5T1BMC1KV49s2OER88LyZy/hjwb
0v37I1pbcM0mpJ14loBRyze46AxLUFaq4aJa3R05Fpn1lrWu6QYG3TqhrV65n1E/Rbg6S4ZgcL8F
85x40+SVWBqw5CNx8FDs0zJq3cw5LvFUzWzimiJOr8OCOIfSlFS3QlWnOPsxwsjWVObw1yO3gY76
hQWgaA/caa31htGAK44BgW7ngABk1gVfvIcGzLPBieVMjtxpcD49WudL6pxa1EdqIFEulOWO1yCn
JDGCKlA3OsQmpl22gE9fFC3JYiu2O6Ds9fWcW/U+ok2uT+1DEVj9/sD+X+9n8hguSU3wONEWrYnm
/TzD548SxUqrgHkuLKASKJicx3E8ctaGzKsisolq83s4LAj8ianJhwXgAnWyUPhK7KmyVT9VOsj1
cz+FzzOwbf1JtNrQIShw2CV/9IaP3QSz0wojmQXKLxk8V6aahpw+RVLipW3SJb+5Tqh4L5J+37xB
/wQ32aRS2/Ji0g6Gmzu9p/0j9VVWonOJN3Nkmwx0lE5r/PkBPMcKaC4yh+2jvm4d6ZY97WQJQajm
sxDvoj5d9bcovBAbAkvQ0/1pAKGMn9muGueEU6QQwZea8rCMwZLsNnOcbvDbX06ljcLaLIdu1qHR
QYZYKX0EKwpNsfwVAfG7Mefe2s5o8aeeS6TOe4zQzjQqWdfyOeL+4LQC6PrfQEhLitkH2a0JjfhT
wZfGXH7dU6B77WZy5eVRpebX3Lt/ll4vnUVXy564uSmSiSIIewAOCJt5RIz25vOl1IGiPSbGISAe
pYn6p2AvwFtHDWUy0OPfE6ZFNOUwHSbQJwFeAg8LWGUnHV9KsiDDiwu/F4Vf65FChgpTaMWMkVjF
3nzoNrs0PuXqxS5xtpPOQXFZSnn2hrNehiuVtXI2FKc++JcJRwcSSB2/5QEk9+wYwMEEb0m4ECUU
ZLr9shw2j3XZkx5PVx0joPfxyhkBw+TpPdqI9y1mSnkQd6HcUrXUuHywkBzq1EXG/g45NVEVVwgL
58g3IjX6F+Z3Hlgj8B+5tuYvPoNZ9NkyCfjw03j6KiXc6B6Xxmku+hKEnMpIOrPygvpkHRM+9vfp
tddq3h8pxg0idR8eQPKGbwxDj7vnPxub12votDs9OHOTXTTNKWkiqHFK2tlyb4X1/6OvnBc9vPJc
31F2UCvdcr9FS8LZ8HTVaDUlqh0oUr1GxCP5VPzh8JybG3nf/9tV/277DgQB5HH/XimB2dGuPqud
cK3BQj/vFQCm4X9a2U43Gl9EXsHOUgJ8AP01QBb+fCaal1sy8uhWqCyrQYCz7T60dmEbe9gA/+/s
ntV+Z3xiShgl7NPeaDGmb9PUvaS7YUdrYGX7Xu9n73/uZYAt3GwZCPCXoY+O4ipAxI0wkPHQ404I
piOL51S8F1YqiWiIZBSq1s+cauZpeGJWE6oknU0BA9dSd98hmAB5NW+zSTQ9M3vo68kktw4WP1he
sovs8m+sw0172B1ADd5vRP5WzJDgHlVih5oCiiTXBYQuVoHrY0vljR/GjvPhCb9NVIanoxNWcmuk
ulu78X2FLJKh3QlHjeo1uPRG6lu/usgn19T1ISpkilcEKFgypPqDWCCGG6MPADMRl1ekEWYRrOAW
05QT3MTGwvk+VSZTjHHlWkhhP61ZCtN2QfFzSOh2Qgsl2Jp2luayopJbr4JdT6bmVgVdksJAMPd9
P6WbfneFymjifsWLCL/6Qsafe9WvqyRapUN3KaKZfyDZrBp3MsU1ghzgPvE+xSQT/CbMwIBiXzJO
jOx5nZdkhkzkWUsXWz0CuVFRybtkaq+n0O+O6n2GlycF/3I9UXYT0TujS8tgqpWB4FE3u3Gczm68
evOqyCclqayfxyujAx7HO7HTro1PDrKyImWNpDXEgzZ1u60SlL9JHh2eLCAeTHHnnDCO+DQOwUpi
soaQY3rSUmBRGM6ihDt7hpmbLxJCzge8386fpxTLC1UNTbtR0fRW4/GFNH9VNLakek2SF5rtVwiO
KOokviz+hzL65bVxjKCliUQImchbbz1wrgsRnqx80ALVeVahCHYTbReirWklgXWTj1xIojFTIvX9
gaIFBCVIlYL1hzbKitIwK568l25Fe1ZrkHF5vNbWrSrakFD3M+Gvl6hqzwRg6PgoiXlqVm5YbQmn
aNnto+hpvI/DFgdYZIBLDmYvd9lbzqwWjGXNdRFOPsZONpVl2PMR/nTZ9Nnuj6I8UJjXtjZpWvRa
PLVNrr27Qs8NWJdpIfVUqTEdLtOum7zzL1k4izD67AeyD0XzeyVJdcMbtqVLml/23nSIjh1ngZ08
7aYHbcLvrTJI8ExkGhPgSCvdDVr1Kdgq+HCAVLjez8tRWIwCfDy6TuCru2Orap+XLUucmnZDXBdY
Dwpg65GkFszBJBLFlkzPWSYsTMcvQloS5lVr0ipF8L6Kysfes6/6EEJdnvMmBS328BPki+xR15+w
EKzgBqx4NVj/jKRXeixXQ9te2st6dh0P+DCM8n2H4+gC+vx4NzQ5ByH2o3bmV9m17OlTseq+LGdD
KBOK8rjzyqY52qZ7KhZ0W16sRH3hDk3SqYwkKZ6jShy3QHrLWZMKOY3Vbgk3Yqld3K7mAE+KfRgQ
F4M5kVLOwwz5lTj0Eg8+3xS5cQMBakfAsObEMq5fp4i71FS9A1rTTwqGT1JCSFfmo3/jp0dnHYLc
hOmBlP5Kg/Qhh0omSMGdPbUju5L/j33abRhQqrgRfJN8azXWt/0/viUb7KXQtt66bY3iT1EMouLy
E1C8P8iO15jpC8+mK0VklRpN2qwopHXP1Y0EV7oykRNErz2Bb7gVjM4UfwWrulTzSvVsxxPa6DA3
wgTpibtneLiAGOsUDxGRCNOc2un8EmXbOa8RhqiF4aTgDqZBGWqYCOBIzj+xP6BQ7UOINgXbD6Kn
BQMApZsCNWDzNLKguXKKhOoKtG6kNwURz693qwiuOed8Zv+vZyHeKdK+uJeNAplHj/zh8Bgyshw3
ywuYv5CmfqeZ0KCYmPDKYG7xqYKZ+sKJ3BS69g0SICfnAngM8V6vdagh1M9jm25yGataabsaPkWT
PIah+bSGcGyk9QhkiKZBs4NED8nzSr4IPi4mfTvtfPGVphBuGM2bYVtQmkb3Fpd4JGDxGSo7jYaF
WukFhodFkkfH7KpPbNYsC/xPApGEjECDyttrO5vx2ZOaYg+rDEcyD4nP1k0G1e67depu6dbEXIHf
qQDg70ckKDzU6K5nBOd2Aw5Wp4n1RdaD1AHkYItLur5zceLlwuQr6OLffLE/vsalXXd2QYic9blX
aySFEWqgTOZOrDqNczXRXhPKFrfOwujN0AWHxSBHfhtDrSU7TRuJjBKBI5GUdo6wxGXFsrjdLVsL
As7wev6i+bfu21Ne7hFI+v34d1cl/QlnPGtrZqjcm0sr9WIFEL/Ttq3LfWlxhgOB+/TgbwVYnUjA
J7LVQnPJYClY7G023aB5VSbt0VPW+YNQYjzMmrfWleK9MpkRNY5wKCBRifuyrFGgnSK95CpvnWaR
S3B+0047Gl2o1ckHt8zAvmjthys0h8apVI1nh3erAeqPe4tI54Kp/2N0Ji/ZdnYRTX/jMyeUKdri
MkeC5i+/AQY4I8/ekUiWhxL2bl5mTL3VctE+PSZ8Xk6kCdA0HthLPvIBEQNy2klI6Mth4P8tO1n9
UqP+fb0OIMhDKkO4d1BHLcGcea7Z7yuYrMcz36MHANYBzZVecmxa9ffpRDp4kpqKgVeMyjJaUEq8
26pC7VYaAx8VSjJSb3qWpjCqBjJ52aRiztrpJVvLc2sSQ4coS43Be52SRNR6+6UtBm23F59xIQKe
h6TgLhSoii1XLbjoNj1mMWKjV1DHzhtLX5wjnR1kqKMYK/iSVJn7No4zcaZlkwkJi7lINyYHgCLa
lcf1VYrMZ2+6aBTWffHTZIEwuxQN0uQB7Pj92Os2Baa2hSWhbu7kbU034K2r0knwM+P7xcKl3tSq
sTKfIKaAigfv5jeDAmCYaI0arV3mfRfOklEGPtoZTZ49C3eldMMafArhgQCPL0q9nuRTiAU4hyTm
3wIhPoE01hN5uWtfJH6fCgv54w6ffP06KpUG4NmAQxUB3HKGXuctMdgSrVJx94mdkXqxJyRHmjXa
7jGPzK7dFyg5+hDbP76uyl4IbMMmztW9wqtub/yckXFv4MTS3v+Kx7CpS8qUNO6W0hLo4cY1lpRJ
s6sqc4702Mf2Cj8UTUQ6ryerRvmZjpTtDNsFqGj032tA1DvlZ/Y7g6F9Q5sfrRJ7PQWTfp9evNP/
YlDpVxU/U55/Zix0aNjLXrxbj5es2dGQNU9uHlqNy4kH+QuQ/oF/QAxgj1GsAk1LDgJ6YJBtRrPO
+7H0xVlSfcNVYUNrNynrcaSXXghalwpMXnCJO6iUk/Y/08WTy5c5NgIjfXW0FkSklCw69RVqYVZt
/ukqZA/pDIamQ6q8nMDLfWmepe9oJPDRqV1lGIChY+CkXCQHSjVHzKbHdUcN6d/6WtG0ElCF9Hp4
3DCIwqe6xbdK53LeM26G3HLlEBa8LvWO4PL8X+N9R0qivDQhQ8ElJoNj33nYFsTiAXWIMdOr/Wkr
K3/MmXZNHkzTo8RpvglOMOa5BXY86chOMoXgT5nbIPeNmP6Zn5MstGM/796Fw0YPPdkuFij6ynNu
J/mK5o/i5ApFdZK7TzerEW9Qe6fhPvijgYvWPkXOdc/U1WzfIE7q5WJv1rMYUO6E02fvK45KzpsF
h4ZW13sW7FsIOU4kqHxAZ9OB8ni694hVGE64olh1335UMjWyrovEFSM3nr76cAzhbEaMbo9kdWq4
XMwfsM+1XXXF5oBaoKHN2M0z/7rflu5UCLr/GEkwkE5NvgBeY3FoeIODV3+bYvvf71RwxLSgdToH
bb5yl3rlXuUDiAQ1eVj5K5hHECfczxtiCIYbaA5lJmlSffS2/vI7QhqBJAJze7a5dURbr3J6MLaN
9Ad3BFLP6+1PcYzDVc1ffk/WQeEcL5XwKZNuCa3z0W0BeODOzMN86/bTVXH7DPlrIF2sEmSJgs4a
kZVYtAQMs57jn9k6lCR/WmchUwq5+FT7opZ1FT5C4c4bV8wcXTYYLTX1FnlJ2mRwOlI7hk9clV/Q
tCVHcd9zevUwLYT2WQdZUBqo2x4Fbk9w8nLA1auyVFlRycVWuSyZP+zxNJI90VurtO9b5/Ieo/4l
scQWuUY28jOJ8O8yyAaQ2g00Mpmrdunbaf+zVFv+N7ZG1boOm94aMKHAT3QI4t5byO0IXNPkj92v
kINvovoB8VRebSI5wVRras2XHOy2hdVI6MehvebZnzwqZEImS6RTaDaJFdEfU3KGrVJQgsc7/N4k
ECk4RoRpSL2LkHLnvSNeVd0K+dQ7DHzvrCMibr5mSDjqXF3lwej3+57cHGjbS0IyFXa7QFBT33eb
Oiy3DG87im26o5IGxYDqt7ElOAJdbzy6/dN3JmJW8ODeaVBCD8XHOP9X1wo55OmjHkb2zmV+rBJM
ylf9iGKDv6u4vqFlBARUiAhkeG2X7EBxo0POafoD/315WAV89hJ5HjFLE2cdpNqU4D3+n9iLaGeb
nDFTBUXH6cyPOhMAD2DwD9lR1mcOtX3rG6BBVcVWriIsevS3SOJzpldhYOd/Bc1DKhllkAOAIHnI
88qDhfYgOlGvj7CqMld9wpPg0+OzuNdaAzKkjltCHVnOKDrAjQQY9SLJGYO4XKUFvi0UMZHqJmkF
hDSIir/YQ4+qoqlyc5Rx4sb82vZREKhZlN4xzye84bS94q5olZyAPw7I2mv5ScsSEiB9hZ8GN8c+
Xncu9aYq+AZAGdtynyOnustw3LJVrVp6DVYu9uOWpUIDJOWrODSVCQ1/SI3395W0507PuVo9EWLT
pRsa3KhgYHFySReQK2TNbZODCsOgde32xTNJ/XVmJlTLdusA9xss6LqhDRNrH+6p6OaoKd8TfOK2
FTx7pg57P/5OK0hO+u9/umQNbiIMh+QoVya9JAZ+EN3FmeXzFfz+IUXeRLKty7gSajtXuGUd1u80
xJvjr9rvxNmyCDTDD8UtWl5TxMQAFcFziyI1qizqWAyyD6imn6aLyXwEwds6XH6eJw+R3RuaK7+/
VmmG0Wx38ppWseLMc8+6WLLpCN+DFQFjDpTgcN/LDP88lioLGX21IWxMmEBIx7kC2pfP7KaPuLMi
qS365SyO160Zgivh66Ecf6472bUX6PetPqRTGcbY9HFyIGZ9n+h2OHyXYZjD3GxVhdpRWY9SKqIu
yvant5KWTIgaVeK+Ojvmro00FuElD7SMI2zz/cOr6l7FpjinK5bJAd274PS3wrA+SEfLvRR9NhEX
00iuLKBr2g+QFA7yCTf0qlHsJqYaVupw4pWo7PVhZV4m3IZB3gpkMoR4bWDSQhNG6nDndQl9Zkd/
qIlVPfcrem1syyHivbYnIVwQFwFk3aF4KHYy8WjfBBWOuv3bu72d/csHoXjPTYHKSGpp7zd5MPON
XQkti+DdWBYOiWDokZalGZSHlDNx94z18cVEGLJZk4m6FnXmFwAFLp3qy9MEIZic0DvJeQG3T9y9
kfTMPpSLZkpzVbiKmnKg3quPrJX0YgYnR9/UwSz4p1XF/FOxwWbbkGkLH7sCSw8zv2XRm4M66v0W
hfAvhntFa6JPx8oD20SxBBUjFtiYnUvUZMNyXYi+PdO/VBjdx0Zy1uCAiDorBi2DMHiRkEnyTtxe
05A6m/AqhNzTWr59nDtOcA9lWtYj9DawyTq0lCs8WVMa3k0pRpgm7kH5lQbU7aPfI9ynlUgOqjjc
bw056pU9+hzDOm5EO23eWkiwtHTGlla92gDXYeRrUJNZ3k3owRqTCnRsdXRPml3TJTQO0iHsmGR7
Icx5UMJ85KUScMZ+KZTv67TDELU2NxsWYaNOeLELpqOASHAKM4Buv7q5xv7YRxHNYMky5NRRBDFN
l/m2ttKRMb57h917ChXDPNGHJG3REcU+SRUnlA29EdvkENmQ0mbFRFFQS66CRm3DgZsSl5k63wvJ
hRYPSVGfRbUW7ra1SwxCs3BW7fMp6++oEb4yTG6iDtna2Q3J6rypWaD51GHhSEpUDOTDfUOOusDc
eFNEn+BnZBLLuKJr4A26NG0T5wyT3kbJvtiCeW9iwy4eUnTloZbz5Nxs8k5hbotIGiSVtKA14+U2
SYlVx9sQ4voTTeWTX91OXq6DRdOHGynR1vSyYR7h1r9MP5OCPkTepbVTbR4ho4hoyHkWEgmWhKw+
bwqnEyLfQeAaV6AgG1Fe/OmfSXmRYRpaXTVOi9uVS6VbHN8S/BTdb8+2MBtNZ5yfDNNqF3LQep/x
QHSAIlT+fDTtTcTCPpoacPvXhK92P0aO3lf73JNFGhiQ+3QCtMZRYg8H9JbzLfd/p0/Jv1HE4LwJ
5DcsWPOZtRwOlUNgERMNX88rQ9Su90hhuAI0zAEwJbiXPbfhrbxWEwHBsQ4rFAQAcsZJwl3Er1Zl
Qfjz4dIoOmgi/+gQ9xtqZrKR+8KRKL/8MQlOpYkf6ilpN9luu5sLrV7lQU51YqG4DdqOhefSttpk
Pm1NJjEH+FaUJ+yToTg1zV4CUJoqO1eF75Ts3ZpHcX/hNRUrPOKiSdZ5E+5xL0SyiOZojOQA4bPF
eZbvw2+OMHlcQ1UAAUmYPxQ/sFtsl0wEciAJyWTgxYVEr7o9sUrXRGn+dcH4WwKYjyrOobrDIcv+
9Gps+2Xu4XQTcXbnsh3rie+yiKfqvjxJ6Gp/1sEpuNnCNUq0qutDx+DaKwjgWZNSuHrEJ62MQ5Hz
ZXisrxLLz8qChOkKdAUQguYuWG6Zivzx/iccdoP9Df4v9Lr+ohF4+iCbxxnpeOSl+WJo3Ujz44vR
lujs43uySqp9UGNyZVhiHf47uOHT5KIX9x0eXxc6pwPEF7ovkKFtXHVphgUZkw51yBedqLZM8mFy
tofr6r26EL63rgPkcM4Y3CtzUth95MkvuqLurQpVrMH7KSNaEroRxLI4t9UpdUvrAbkuDNelp7BK
Gtj57Nq3kwObS9i9eAZSoFxgnNvQny/TN9HXZonb6MSSb7IkUN2yBn1WNUYfIo2+/TfrLC3nuzkt
IZXhiuRmilKbgZV9eT2YgB1dKGjFeIjPRYbFGmrqpdsQLhC8IgkKBtCAu3p41Ufs4rYarw/M2CcW
tL56NNkxpo++Xkj4d7owX2wQMW5g+V1zqMe2ohh7Q9Kpycah/bAhfpIdgOuFtM0eDvNltItYPA2F
LbAITMbcGi4UsBS1ARKz8b0huXIfVzcG3jwEcIOsTH64TZie85Kd2KmE2DnlmgP9GZ2qPaPinbFx
NZswlzzfEcLMJaIXyXYnIoA+NLJXvpLZFM3WOUkj8NWl9f8oL1I1rd+IvROEZKFMcKuDUQoIxfXV
7CTAMlo9VRU3wgf226hrMJhTY+5lt8x4NAW7NBhpnnZluKP360tr79w8ATZW0M3n9Y6lxZ5QBLIX
XfLvEiHAU1yDP1H22VApGV+uxOiaa9BpXFUu7kjT03ujUlFgW6BtiHUV5RDrPvrQUaZHaAvCF0KY
iOdXiuR4xcJP4rOfqBqsZthCHzxxJpw44YPoSeYwM06ZC6JwazhgYNPKWSn2iQ91IkpP8e7twSDt
OwxPLEnrAv1IIoQuTqmUpOIbqANN9K+A2aMo8gdlNi2UcnoTlnOJwexm8G/ZAvay2j5ArlSSShHo
F/s69Kq4nEvgQ9SAA2MipIJDOrZlOBsAtanwKgSHzwkQHXTFEgeevA5fsY9pVI5JwgMrGDoCLsUQ
ba3xBO2auWhEXopOo3JlgzRrxf8V25iR1rWMJcFkf9Ur+VMVzOD4HlDgmNwK0v08QbXsRKrSW8nJ
HM3gTnYKRl1ZLty1T9DNtQrC/MJCNQyptExz3UnM7AH6wpdQBFk2uPKUjm+atrK2Y9ktSTS5Ked5
iuBxnNP1oPuCE2b1BHAVQLqUxaiViZb3Geod8qpLmShnS+Li6U7asYIcGfDBgmYAHlrjFebb75ul
kbj0+csCErQtiFobsm+r/jrEFeBEtxfvbBHO6TTrUKpDuD3dSG9aiovVPLrU+Y39tAprTPt0ye+K
VzIpJcPiRd3pYbmbzte7rf1P2jEBRLQOGvUCnYVRrzqXyf9HV+F5nnIRyFYVEYiWk4bWiaZuG4oV
LWerMsYiwCxCOLqN6FZNjcFXAun/eRu+USsZiRK9ULplFtAEVb67QR4wcrNHNI/gf/++G3frsTLq
ApIc5z+GttOvJ/IlGCvKS7Wun3d4tq1mVjyqqWfnfUvohBquwBFru9Nq5zqmpQ648i2bJIWjPN8c
ql5IpVAn7utUqGsnbE7qL8f7A3oH4OUFV9vB0hwNMKxWp1Z0kKdBOXUXzXbgbOjwg4/P0a75ax5P
dq0CMILpAsiPh58kfPPThGeIUPTfCF9ox88K2fm+yAfLuP6EJ4OyB581gtB5raArnVsFMgbxrxh3
AF++5NR3Oc4y+/OttxY+4icFMxz0ZMQTYnS1JnE9Mg/pArpSVUFLDNoEnQkhtxaLORGD5ce0PivI
ToLL+jZdpkOvWdJyKXe1SqHaGxYvYrx6A7MQlHtzU2KqXnpeAw8xqvbUgXCz/CbuzZKBzwEjBunB
f67ZOe+h9wENivwYj3bsV7cuuP8FLpmJoMZapeOxOdc6RqR0IpswYFSIcUODn1jRBthbQ0tF3PxL
PFVDN4mP8nI95L52mZBDFXWVEvXMp4NdqRi4fgSUuEyS4Ksdxz9NkMObAOQfLVP1vhn/6TOy+9yG
PawhX/RcDy7EaeXyytNHjMGIx8P+XFvHVjlgs0q+gv1VFalaHG0kArfgMsYurCe90m5yYQq9iIfo
O4r2NnwZFI7TtY4H9WOl2f18dhCvVF7Garix9uLDytVLbDr4Fa9L4ylwWMltEkvwonZERV+0e8wR
qyuGLPNwoT8QAqH38ZOETau3QA88nPLyGGBtR32Y+U6V1jHCYOp2NYlDUFNg5CRCiC6RL5PAO61G
eZX9JvKk60iJONfrzw6ppReY6R1vDdBHDZXV2w3ENkU28uvViiIe82mELTFhG9oTN6jS8pOu2rAa
dh8kyL7i//avtK+8ndRvKShGX5n3mtuWoM9vpZml0jCsbL8uwJBDvEthyWekbPXTSn3F+8jtwPGs
Q3ltMEKjO9IB0ajb9l380GlCcaFHJ2ov9EPCCpulBzxsd7KQxlHNtroyg/SWwJNIeiHfJq9tys5l
liPVLQpPfzN2kGxFzBxYj2p4RJmQ1A9NgBo4ZRJubZ8posjf8xzzGCaPyRzB040YNeTmBT0N22LV
f6rDZY2/uJvt8qOpmNNp8kbQXe0OdMcsju0WYrdX+v+gTHs+35isMA7oYdveXvbx7ZNK/AQGG18S
Sk0faI1LNWUM2hKLU6qOanyYxVmo9a6uY0NA2K0qhtJM2fPq1g2KWeiu1QWR9Ep/e1Xi8cezogJm
ULBSjtoQNmQ0lgZ9HNoDEIeINwltinjKrzN6aq+WOMK6150Oslg6dJ5zrzPHFcxssB5DeORqkBL9
/zwLvpzC3TU/1I5Db8+QP4icztfYOqbJBv6AXDk8VJp/1Eeh/PI/nbfXZvU3jwXV1hXLm1BaGcWt
p2uVucSTKn0+17+SoEAlgXFgSKLW+z9UjBNM97c4ifXG6OglwE5RIZ08/xdEEAlmcO/Dfamv7h2p
VYI3kahqj6xc3yGSyeOuEDNCuE4FOAtK+emONhmU+L7wL2aKSwSew54jRXYdHO0WNDJZ+wEfK0Tm
/JWM6+kYw40pCOND9bcOZlhvOhIgxGQd+rAAU4e6lb6X1hpm6fnn6TeZRs2V8C2CPlCdu391IFf5
4A3OjXFjHLgF3VqeDIq+uAU2NOfRHlscwuhHofdP7nid/RgpA/+UTiIaahnnOkCPTAGTRi0I7lg/
ooHuh8tS8dA9R4Ws162OrArShCMiwPmVvL1gaaiuj1zq812PGryvR5tE65nwyxS7qWVFVTw0eiJ+
Mp5f5sH5tgnZ20ahBjcLMPDn3B1JwV1B4p7dtg70WnYzp4eOH/AN/uuq/yxXctxxCgtLrrBP9RzV
HyhCODBVNHYPsgF4nDmSFmpKEzy00XIm9E4av75CM34A6SISd6Wd3pq9S51LTFsD3h93wRhMUGlB
EpraMSnowDJN0/+tSfOrK5YAOkdqPthPqqspQOu8pdQ0z8oudNYWI6uO/c5dXibfeOgPncJEfreY
jzo1tUauW0TpOumr+91ucma4XVsdheVtV5U90EdjUPHZbSp2iBri4abo0bmcgRH1pAOk4WeeGHEF
BSJ1BSqduQaJUntsUTj1g7Z2h90+GWzGD8EvMarKrvd7pc3w0ZmLUhMTishJ7HSTtqc4P2Rjj0pX
B1fksmqdPYqiWqLm0DFTjFWR7t9967f+DPsPUfaaHh/QWnlZTYfzhF9TnaFGsW/nAO4/0W+MYADn
I2VIdak89vK1Kw0pJRc6WNyVjQHoeRuw90wniv72pXo0HXRO8eBB5aqUSeSbPj8pevW1NOpFQnVl
O+KJceUxDXz6Y732U4ro11MADE0wppR1K8hAx43FRMwPfyzYQJ8jL25t/B3EM3LbRqIwmBLyMlSj
d2CxoIuCzDCyJ4esObug+GaQ1Hw6ZSGt4wU+gMtD2nU02n4r+oJ0215GrZSdvWXNI03TD97ojVVA
/jbScbwr3TbSE9L9WanczA9b7tT9fVYAnMB3xq9rertSd8Y8sEeWA84p/qNgFhFq55LBZJSefLH6
37uOpzV6UCBCfBZoh3Bfho8R/Mk6zAKHT9h+xZp9HslEhHdtXBY7HNY8fS0XDjOaY6zOF7N5qFK4
6+H/SJq8TqVG0aPfm5A9gTtL0m+jRKnV/eJnwiTG8fL165DT/0QfxwugFeliZ2MMyPIEwswYve7T
UzuepEQzcJ0mVV4QkV8/5EPPMBEtlLyaH9f7z45gWTUI47CC6NqpRfLKpiUgWE6coz49DPpXR/FT
KYUOAHd+NlC2h8kf23HgrZl0rNEuHYP/NH28/BztoG969gX7RQeqWhH167TbVg2M3HfpHeCtc3UA
DrMpMPBU9NUiUN4BpmjvC2iAByUlLWgRDFKR42ei9pP1xdiEiOHf59tTl1wJjumjiM5mcKYexP3P
rlQooqqfGkCjk/ofTjTup33APFwufDrPBqZ+Qr2emkdnNP82vuPSMh3Uap1hR8jaJEPJjBdlC3Ba
iEPgRvStxAa/7uVNlRyPqm4mfIkO49fSKz2PGgFve2hYVBFui1eaGKRAnwgulfbM0rmOhIR2fpZV
QImntTaJWc7Sg67Umg1uLaU8CXQmTbdm87naccOvW28FCBKXWX5q9pirmKHKDcOLjn3As893eaIV
AW3KQNn0FYk3EnGznqE9UUvAHb+XWBGbnV8ey6/7D8CRMBGQ+yTNKXnvOPvmdx6wEjH9SH6EBDxU
kl2LGKWLV9XydT0pgdQDQhufPsGCpqN5HhlKBllO2RX2OfqpW3LsUbXLUPoRUOjx1qRriq57FMnn
GyycJpHdsutpG5Y3IC8ZBNl1FjodrVeYcKq4pgjPNRcQ9OJVoBPNCv0mNj4/sW1r/mHu2KybEVEE
P80zrmDZEG0dhVjROKCfDgkCwzTUkSTguCMoU9SICW87/CBcFLdL8Hsvv2ftWoQHo5lYMc4/inG2
Pj8wWM7kQlIrMNcWZUx1AcWWlasvhhOMWAExERAyHG50tIJ8LOheanigkFAL62pDAjyc0HI7Sxi8
dmhf75LMLbMz0eygeoj7TRIRE4BTLHhXIe54Ht2jjQDfmKhjXHpCkjJh8UiSuXWHfDW764k9YN3n
jdq4FfSHn++XKzyHh6B4bADFBlG0Dz9+JeC/3S7X9BRXQh8uW0zUIXAoSGEsCCJM9eB8e3TMNk9H
j72hPEJRHfjZqv6iAm37sfZsW/D4KQAOShxtbMloPy6fXxJfCxsU/71Vt08FLZMhquPXRltjHJ05
laNHA461RYKXSMVDbSGWptpMUTr8GgrNDAQzrU153qZ4T2yW6yCSqvQOYjDMb4rBiq0/3tqU2Q14
ipeXymawZov8weuO7gWV5kOs8kn+JsSQARBD1BUMBEhBOOycD0+LmA7xzRrNBlBv/1n1bpLu9qs8
QA7Hsu+fdBNyY5n4gzIJd++FTFZ31+DxeDMq2ntoZfVRgU/IA8wCgPkBvlUIK+kl+qtFJBjBqnVZ
1lXdl0r2nyE+0weOpmOfsowJDGpOTrr9TyJP+16e8X203pAtblugwGhEwgAimiy1qaIqg4Tp876L
IQWfuXcs13eOCCoFeB0xJinnjefmAByGC2Bvqycwavu35m/KTJcldNl6vR7GIvMKsV/xLxvoBf9Y
y0yiFyM59CqhZM+Z8id/fw6PySdVqyFddS9s5A8gV0qQZg99DE5O072YqfNuyPiG31/dc/6IgMO3
iEDD69swyiQmHdDHdweKbL3G7/JnSXgIk3N5f17Zz1ywSVUQii2w+HX2nsbPQuV4HnxV+wDFVLkY
zhcyCYZfwIJbk+FzEhCDmjcRF7jcEWJ8f1uj0BV72Lg6yYnyhyUdgn7ighoRA1J/K8LSjPQ/p2F2
HQy9/K+eer36bio3ooH96PZkDISHRA+GX3/+5H4frSmYRzKbgdzFGjlYQiUBZa1xTRXcp8QZMZNm
DSvpDf6b3jyOi3RNK7HMZxlVZVW8i3U4YKdZ/vH44yUtCGfFtYSYlYLWXQhI1NbRnRcUY4KWzGiI
jvo60hRXcEpxH2c+3qiB2cGStD2sBGq1k+NvVfCGotGn8YU0ZIF/5RfpUXNSxrYicfqBxtrdoIrb
7k6uvDjhz54dNjv0Cg8ugYHQYm+auByBlzDaRpMBiV7G6paJo0jJIwagjh7Orx/2KaElMYRCn+Tz
rQ7g0ZEy6tI+jCx85PhgCHgeqLXoEXklC0XOCEUFuxQP4QqdLQ4Lc/oMGcJozRTD2zF8E1gtu/p1
X283SCI0GOLcnWQRVY2FEYPjsaxWBQrgLqK9qvkemKcjnkSZ6uncWT+rPywXOxXKrCBfEA5BjSsy
6FkOsopmxu9u2sZ1PYLchZSEWK6WIdxGNAkZ3cDEWunMpzt23UMhtkgvORWI1it0a2uQkC1azRkD
8JWlWWZI5tIHbX4FUhSRFNL4Y/gAOBxb1o2t48s/iCYRo8M+biDs5atcAvNQ/lO8F16knB2pN+Xe
ukqz6SSBXBR/VcsAVvRSDKQrr8iQjyf4DgN7hkflX0VgoUyXVKD8irgW0XOJwNNu0+GNQ89fly7a
BII41003x9UI4SSrCX/nUTwMzFWkF1QFR/WYQfMm13xHoLtB6TW9zv/8t02sd1isjaAn47uBuSZR
5vSBvu5YsCOPhtzsfVYGd13k5XOAPbfhKwDv+YCQycQWyJodma6DCXuQIy4NXfymKQxMJWVbZrZh
+2//zN9ErXUpt8czj8dVHotUvMd7dZrSeeVz9/Foi6WyI6X9dqPiKqBqe8Gm+tcZgkQ6cu5ef5Sf
bpGseAzcUtTC9roZSvt1Va4SK7b+apLhL1rtCwDc9fbCaV/TEUhLDml3P6EiMuUBtDS4nRO2Vxjb
HhCURDC2UdUdA96Kv17z5/JIodSnN1Xaa+SXqw3mIMYb++zuxK2jfhGRINy2JcBH0Jb4Vm1fk0qg
ICCGOHWfbogBe2AqaRygYVRASt8ghiqzeCnYiiHfVGxz9vF6mWLnvTT2SMMrHPlCopKsx5fs2QGV
4j1S/9hr6jt3nLcbhtAcsYdE+FFd9wuN4HNiHqJNwTOLQklWVvP/dGKGD0x6jWojbiWNLe8e/bCz
wq9NKyGYGVPuRcAb1fSNfSq7yaSIdqYn+5v5SMxziehpaECLyKfW0QAT9yyHeT0kR6fN1KpEklKN
eY1kERB6Ns+sbtNUGdZv0R8uG1Iyf23GDKyG/wUchVvDZgXQAN+a2HAvEMLmz05+PDSJ+HVa16Of
WEgIOSxw6fqokHsezpH2VvxBogATrIo25xe7Pv/a/e5w+6cVA4mmeJvcnMzkfJ0uLV6mALE6f1ne
0Z9ClvFcInrGKNGnq/hxIJPZUHmlPFz1FxrF0Ufsk2FJ5pyW3+042vWGYGFUM1JaPG24ZZ2rAEhJ
0mXxXUO3GM1vAgdUEidOBBOUOxTT8BrBYzZP3nSiMGtLMnfVDxrIkpD/iP0aGcEL/l9Dq4ab8I1B
A8OOUi8CGDOBmUoCwB+6oE0HG9YkKT3ZMeiL4vVz4igN/JcYwKE7iw0Pstw9lLqZKoPu23/gMKRc
2OdKOyyUnNs8RAqv7tcZTnbfvOGN5k0ZO3cYxDgM1NF82F/ar/bxX0siuqcIoz5qjNjuZuuUUH8z
lhgE0Um1F+sRAPMx8OmfG/8H+pJHTyjHKwfUeu/eoR3BarpS9p8t/WbmPgL4JZaa6tCakiN1d83x
G9hOqSUC7hvyrh6jJ0XJy706IuMABpUC8li0QyH9bM6fXpohIMJb0j3NjKJ+yHNCRWU08mK1Bl1s
6GHm8QXvkarWyLySLPm01lI1nGwB9M6hNq3Q1MtuAr/qxJVqWVH2iyBFZ6TJK3FgyhSsCHfjq2lP
0KatFl+SSG8fLOc04uVjtQ0iG3ChKsHwqs0O3gZJqhGkdJ2/QjSnpGpCKqeQ557Q4hEGBbNs3b5g
S/lNPrlDsNEgZiPZYgR0mE5/XGwvEzKAea7l7tsn7/fcU7mL9V1yqz2PSYqnaTM6UZPD7CBVkMjN
Y7319SAn8CY35aP6iNLz7PR6wYCDdiak3DSLBFPNh87Wlwv7Lbi2Oj42O+epMO2VBaBWKOYwAvII
/emwnmvOWE+tFbEz4RgqZ33hppy7EUMi+MdNrusXVnRSj2gnlLAvkSCTkdaSFNgAS7sSBvWpAF1O
hXeqm+yqvfKhl0UUmSu20Ajnt1E2ESE95+2JNK81xauLMyEHNvR+g0fbc0yh1sCOehEKAnH917D/
yDuYNoMpCYJucm/7acA8LixlvyDmS2Lc8vwO+pn9ePWcKK5+KjfAxNGasJUUmAltf3UsIBHvPaZD
wm1iO0sjDf+WkE7bhCJtZrj1KzTRqIFG47YGUalj5cuHk2UdxOvRz6Xcc744gYn13U6t25GVUn+N
pfJJKmJDpTmDSqe7cEkBQNC+R0pSUZTuD8wAi8C1ygXpqZ2cb0Ke9Nf+6Djz23sGaMRStKfLtbEf
2wAhjrLt0/5FMwE5pjkjcUGFkyL45/Ol+/o1Z9sFscKdQyDEjEylm+CeUTpDQo7sT3HzcZbcLyvy
vP8FMiu26OPxc68SNgavwyre6u43BhMNRu0fs21fpA7qVy85RG15vppcKF923FWcbVNTO4CILTkj
AJUiSPY4ptR41GYIhlX/8I+rN+z24dRI+oWxMLmZcQtZ/jLkliOLmrOYVvi+GVUHf8OFXoimdKpe
OCvIhlrEv6/pdVvq837qXCSHYTxw/RPlWe/ZCCVhpyEQPrVca4MQxlGE/IXEznAHjqz4kOcza9Pw
15UQWFXnd1XT3mDzZ4cDhg7PWnJ/95oiNV/yVpvDepfXm36RFYpsmAxvJ/y9cZFNn+fGL+h5VBUo
b5PhhSK6PnWRnhoxtqwJUc4pHiqltR+Okh/wMqTT10ueiONEDduoJYtDEbySzUH60TiDDyW42uWy
ksnq4WKnTYMtla5VacyzAnW0NF0+VD6oL1AdjnX+bnS5g2iGGG+FuHDy80E5CuvuSzQhWItfMl9X
J5JHmlaN9Zj4ILNOOVyDkSmyS4STHDoCnLy1Nyr9D5TQlRHmqY8QE5Gk8d7qB6saAu/8GFHot0qc
AljuLWt1qBZMAElDrPQW5oYqPNkjfRaUm+xrems0iDZmHt2YAh+gR13FyR7kEv3y8T8sAqjzWZw8
OPeWGNiRUg92p0lb5FCPFs7UpjTlx0nCGbmf42my4Xbux/z/Ixbm1DvzwZ8n479tc2whZgYfUQso
q5rHI2EFD1ePlErurjP/N7cFVTeHIklzOxvNXn4v31ZRm611DdeuhcsoLNVAl6qR3PiQT9239eof
i05JnX9fZjGAx/xmk2g2jFcupwaAWdHwd+Rm8BuJxNrrAyCRE54h5vgUu6PlS9i8WwFk1+p20jeB
X9pHKuFvTti6CFw5GJihmezh0uXtCJ5lUhGcGJli3pQmyLU8QvL+I3vxPgvkKn1VAFSbXrc/bRTv
gr+SfkaQpDehm17kuolgKK+ckYrIJceH03Cc700cMR1gPJnCihvEEwLRnGhkMjhnwGURUrNhuuhp
17Sk0Gm0MyJ/6paftROogyFlTpA2BvW0DNcAgZqopfL5Ua4hzNPFp/jLP3CBz7SU5WLYGp81s0VT
jyWuf0O+gXsBcd589umZurDgO8iPWNbNRKGs2mBOQ2nDoqPsYQOp2zBd8eAP/vxuTK2QIrF9nSOb
hdVMFAnScUaStzyYdyZtzEGSYRvXqYCzQ6XnXxQS30sGrmeQ9rwMs/FJrZMj+99+ve3/C+zOJ3em
mRJ2cwwM81MY3yF3pyt3ccMVECC2yrshkZrpkwAqRHWxuBvgNjVr761vetpz6QGKFEfIqvrOFIDH
OOl+fgtpI23wNDL4qGk+a//ii4fZ4Zcf4NrIdUQpD9RDVRzanqFihpfdRpzlEt0cSehDlHJ5o4K3
dOhRNWkbl0Hi1IrNjhBo0dfRmDjwVuFmdOj8cTHLzAS0lMoU5ArceVfm/uNa7be5tH03RTJHRbtZ
P3NcpYj+aX42OarWMhVBLCNeqiqgnG7UoMrsH9FKhhD1sX5NGOKh6S3hoxAOx2VyrkbxFT9cG3D2
oxcgvgpHQez+KK/qui2MIzXJaSYxniT5BrjVuI04RifV0XnWoJK6y5AoFMY6seqKieNGEKQgG+py
K0hwjA/y7neTgGqpetlibjk5l9GYac16fqozVo9M05XDuNKY41FRG3Q9Vq11rZglm4oezLnDMyg6
32YOoL0to1+14jrIKi7zBp0izPAhsZq54plgTlVIOGOHv/lmGnJeEu+DZBV3TJ+uBC3lrJJTBWRw
Bh76ytNNW4t+KH8DkKimF2joSuoXIsa195Oj3HkFTqDMymICGQlkQ3ojcpn5qjkGYwW/cynvTC7d
yBlwJ9GyOqobSeaSUrVIk0Jouu+07NkqXHNwoz9RVqhRUxQ9i4WVKgjfgQzDwyFTdhUdaZCn6oet
UPfXsXBsZ9pEfx4FzN7RQFAxcJjZf6pmo4Zp7n7/yPqV04zsht8T8xBq61xqAIOx5J6UqHw3EFsL
n2C9yyOe1Gu91k8dU+wiTavFxwJG+9MwvpT/827EJ5Mus7ofMEex1+/ICpKmwxCe+RSX1vjH9p8g
S1GGJBGmK3larYpbTkeeBInMb6XwBOewL6dKtsrWOZHpNR/wuYtkJtdevnvtQpxHeUfdMEe9uwFd
SQPNue8/H4CVWVhGxnAdw+oobZsB/hYeh+dfCIQuL3SygS9YkSkZLcoku0wDBK5e1GSIXDM2U/s0
rswh/dO9Q+w6dMemNveTY5YV3cknzN6J2HeSNLI+yozDs9mK65oUrqdp/uTA5f2KTs4QutOvmHqI
WJMFLNzh2y0VQ/c/1V2RyPI+5XHfp9waA4ek10+7eQjFtQ5Cpzc4hPVAeDLsiuGrKFb8nIDkTouy
OBTpH0YKdEBHFvx3GBWG3d4EbedJ9kDmsdwCiqZuLsPbX4xDV16ogtcka3Hnd/X3mjaunnz+YGBU
VNE0FOP0T0tSpNV4ohnJ4oMzy2zsTl6uBJlSCRLqOYooHE030ReZDQpArdFvTjpIcYP3IGT0daQP
8piuKoHFXyV2c3eNtkDIpOnVnM1pL6vBSkYQLMlxh21cEB5T928Cxm7hWbgm2w7GygLEsRyIPpe3
U3jdu0rHIGGMT4i+VyRm30zzbzAp5JO3+9C35rNoKzASZgsEdsSsHHtyLplf76Bvexv6oUIxzFuO
yWZ08coGfTCinSuu0RO3rI/9EybR+byXUEPc2B8a4+n+8myufoPtWBV9oEg76RdSuEjfjXon6p9B
VNvhqt7mij/EBxnqQ4KfbdRJ8DKH7hzj0Zv+KV6ED2qWabvBomqyQiV175Zw6kedeYGUkq7xWC/E
/OAXMLgvOvaiuhgzCnDC2/onhBTIDoM5OxIpjznvta+Hdtr4Fky+T0ZetDILwLa7gOd0ZxFs/Niv
ovkati3KfPzMm8ZXRNeu8ooevWI0w+pa3JuyK0JSZ4ymi+UutEXtKmOityOdNysC0t6Wa8k9PXpF
UKN8uBOuglZOp6a6CEBbCyMOU9b2bkKcIFy75KqZps87D1L94IN38QAwlcB+0JuThV1UcLMMvcxO
KrsXqN30qn6yvF4yY2xyFHIpS09G1sLL/T0HKLdoMc2H+nDazbhYXnoYZAXSV09AT8bYfWWk8BM8
Pw0kGzEARRCXbpVkkXO9SRN2mVL733DzhQV89S9U1FLUZQ9WGe6WDPKCIPzaDSd2/qS38cMLFGFj
q4F/LAq8pnoIqEUlXmIW916gf1ju+IU8C6lv0AYWYcYL94KajJMAyrZgMLIRvm2AM5bJv00uaBwm
qMDEFOLXl+uEt9drACNaTSUfUs5C+MtfskqRGkz9PKkGyhbwuRlZbZCkB8hxDM8EaSuI7EbM56Dh
d4m0cEmMZDVx2l0uX8okuXLsFX6x30VCNFclLZmgGPL4tTSjSOsh7sX0nR1i4fh8dJNjGjVWXYvu
otZKyymXRAcj1KBzcviuwKTENjgCH3ujM3RtQyt0V9iEvHMGi2rOU8W4PlO0qrphmT05fGmlPn9o
LeAqTU80SPfgEy3tz752FsgKkln2QmXU62uxYUo2c4uD52RBkoX+NC8Ch4ooy+s/8GBMZdL+ayw/
BIr2asZd+k1QAOs8HSyRiiVkrzr/Bs+8/wHlCeghfvyC8Nczop4OzYqIb7Op84mZhmmb3uzkHeh/
cgpBs1PPMgtGNZyVqImJAi53B9JeRx16BJn8w/tCHJ0Q1RAJChtoI8bv/ZWgIYiojeAHnfZzIl7J
2dKW940xmLfPQ3X20wQKzrmrShk2t+I1ASnXyL0JNYlsfuT7siI7aiMSnXKeB/5h72wMj/qsOpIc
v0oJfB8UIwpCIWm4RwkByRZ2sgynw7Pb0Jy0nzyYh2bHicQ+QXNdmDyr3HW4Zm4WZqKJzi9M4rEO
85r/D0YyxECYfuUNYGExUdADV5rBYNjwdAr0t7CWqBpOTbXmtq5ZI4c19aeCaM80rDGwZthmFv2I
+8Y/Xu9XZEz5dNU2KSAm2SKqcFM+r33GevXfmYkJULRjOHJXDPoajmFbNcZuCvmKHGtlQ5h+v4dP
TmFjxKgdg6yBEMYpM1lEGGZ5Sx6LOlM1hCvX/Xw8EDXXBYRmbgJOXQxDvNAzJ4nqQNbrut0w5bR+
OhSNw6BH1E1gJkChmItmhp6kp2Cns1dxjk488moE2bubE3dEaxkRz8rQviqTcuqseN11FQLY5gle
ts4LE/+cU0Ca8XBitiZt2JDVuszdOwb8BQrofgoit2dp87qcuDMGF6XDMdTE+yCw2bRERLAcTyhp
WaytrXZM6/1qtiCJmvxDPpDDBdNCwfdk2EMVItnBHzEWxJCRJ4sBgOMdg23utzLbHSv5plZzkLFV
Iwha+KS9E1+r/0uM/m7k5NpF5ARfIi9RTHPctLVVmEWgmaERtutFiX4qM7kszBWk31/leOAUaBhV
zUVsbmP0hUfHO/sY23UmRTGy7PwR11TIcHrnWm9M/8tO0nVINr2iG5n9L++xEcDHX+En1Fv2kJ18
J45rqDzie2NQXL+lHXi2Kv1aEneyhxez10FstIwSZTvhQpHsgTiGA1h99PJqER8ai2JkWhDxW6UE
KER0E4Cmf5aGEqTNrNWEGgDqPnStNt6VVshdiwZKV0AJHheZQnbxr7EbPJY145gvGAJHbhc3SQIS
FXRDK3mgLfZdlxNPfW9bPTXplka2SM8250sVHrD5Q4ZYT9AJRYZTP40hm+0YbfcFX2AYeWQw54Si
r81Gmv/PyRqF8jpXxg9FOZApOoDZ3GiQctfdCyX6lH+ftSK3JKJzLkeVFo4N86HLaiHSIJC7TdFu
GtEjUW5OZOYGoiX37yn3RDxKEoK1Zwq4O+fROWQj7mqyhEVtaIjZBX+DkPaelnXS1F7HJsIxaG7b
QDxu1Lpbpl6B4X3XoB+t9L1peUHwYCgThg8o2LurXr2wvLiW4PLuOkT0hoFxoCaYbw/YauBHnfdm
1VgY2swWXwSoBOADEV0hot/0w3lNQFfSSfBVXiN1UD+cPhknaa28M00Hlm6ksETNxK5ebCrwnXHb
WiSMpuBXXgy1/3iKbPFXWQEv2Qp22h/8FktZdRYBI4nbdpJk3+Brkn/DeMsIei0bmiRh4OgPvala
lhYZLrU/EDKQVGn6vVoNDfBjdvfjjr34BCtdaH2Pz73zPyzM12N2WDg7Ait3c/YBHJA7YY73SJVB
AMhQgJah822iSF8PssjAsmNI25W8ti0MmupM0fVJVbkuCjBbHZ62UlNvevSqfIHmXOs79F7K0ahd
9d4aksZxr+CdpEgVshMkHwwTyFmemB2QYgYLor8Rs2rQj16FpJXzXH5U4s8S/k/kEinNVvoGIygq
sMJafMkhUsBws3/zCkCCu+FdEpqAWu3sXs3htm4qvkiAbcgd45zYjhcME3ybehoP5MnAlep8IfNU
5oH7jS+PYU1UxL6P2OYUrwfsKc1MpwLpekrg3kHqt+6hpaZDiRQRvUPrxs6XfTDymqGM+VhOYpar
5EoC2ya8707+g7Q2yA00+V7ezCYBbxd/QtwPLr8e+CVgmZkQawhHvbkYLERp/T+VCPZNTVBQRhBP
svPQqy4ef0QhkLeASgNmqVr2UaNC0wp6iSnQhd0vU9iFM0S7kNd11yuPMJaWylrUXAs6d5//aSiC
PgNzC+/UR5ZUbnmrP+2LnRCrbD+zc0gN7XWs+OOLMFHMOisfiR9xn0cnUPWMzEGBEdOFWaKmy2F6
8W+6hONkIgmVjxs2qJGfEGp2OFSR+GWZ7XTNwA8LIpXdQjSXVn3ddle8yS/3SdnHn1XN+PJIZi6J
ncfQtyTzOglDMpXCzTGzgQVkYTFGKx3+L1e1T7AW71O4bml7OGA+SrxHbgugaEdkvZ/tHKuUemkn
un0waGxN1dVl6bgKcYvRy4cNY4y2kzZ2Z31IH1VcqtAbIFx+Ycay6FqvFKaLDo808UjseboIWl6+
2oaYITdwS7qWai+Wh/jwMKldF6bFHFt4CAOK1Jmk7a70ML9GnyxIXLtL4CVBSrn+sOBxZyEKjr6l
tRvxUi+mwXT398HB2BiHxlCAgN3XWWzxfw0ulLmSIQkcBOAeb2nNgr9HzzhZeBVB3Ebbi8cRlpd8
BEsS76lAMNNhkIIK4xp+FcxCTLtvk1ouKvvXkEOhi8WQDSSedcntTVtGzpckJVOmxRUixutPDHwG
0YB/phc9rsLRYmcP67mJ9+8L9z58PUreyepp5ZW7GNXsopU7DU9apkWHOIUgioNJdTUoOech0RhJ
c8Ns2H5gxPOlTZjcOQKxUoNwxZZiM+KCo7p9zJgg4fGM1YAvHmohICM5WJPhIJdeMC6RaPlQphAb
PYANWw0FKVrSws8GOeknisZkhliZxyrIwp9P+1MZmACxJ+R2zHakMsIErebZm/vOiEEFumBUGdEb
8quXqb20QHGZ8WRcBpPRNqB7rTY+elel51k30C6FdO66xlx92MX0KZ2IQxh19jZVofCzOcKy2CXO
xislE/pinUHxL7a13HP7fVHNN8tdCCy4GFz3d4Q+DCgarOQ2ofr70bMGu9lbk20Gp6qwPaPiugLc
fa22gfwynJ56atX4BXaDsuHl672Dan90jxDALLfnxR4wdV7A05Py7/Lwfn4ot+1Aw6+DUqF6PP2o
Jf8dkSYqphMYiRAdLTqVlkChX+wOnrJWG65kG/bXGoOIqDtECFHOQVz8VkaEB+JTnaa1PNyDPRIL
MbYXwtMUJJfrdXak+klXBCObKDlV5Zrz+kpXOuWSXJdmMqQyp5DQeM41kTfWNuSfArVjcw/H24jS
803Shn5QKIGtViX3MvosFF+V6FoF4940U9paed4kUv+8RlMor5o7BDDsie9q1g7ZMwgBCCkSg01T
r7oN08u4KTT+vPmtom24oUzNVm9fsl0qGeNjnZ8R3Nw4b02ikxBVH4ErD00Dphwe/isC+ccj52Mf
EpeSV6t8UdTuuMVe8n0+tDHITGKx2iv40/OnHqvmu7Fdkhiy1VidAvuJpDc9M7u4gRsM76BELEtv
U0tvDszCzH4/W3nBGltsz9nKMUknrLb2MrY27e6fLFsjzvoyxBUq8tMJSFK7qoeCobitLJ62smP2
OslGSjOGpYbwEKLWrHRSTIuz1/8BrBPYmFzNxNWzsfbuDOI4hnfNPzKBQ6GBLlidPjexuOrMl138
4hASJyKFNnQ2N5beH3MRPnCQhzNA6OjoziBqwSN+h4MXMq7Zjrn8zX0/MgwNnyyFLT4n40AlR9U6
tmanecjeZSkFENwMDdlJWCEKXHPEaORl+K58nkQ/5I9/yjsDedS6k1YqgYRSQHUM00sqOYdGuThw
b8zmeM34IyaiMCS7EcAMpYHsTZrry2crqbGMQDdabDj6H5j8o2aEzULWjitGkJokN8OMA9gCOGZ4
JXeBzvF4Y4GqFd/D0nVO0cnTLRwWKZE9TlvO2S9o0g/oS2jEx3qrMDtHBIi5wZO7rS8zhUcc46r/
aCVTIp+CesAKn4yv7uqitg5ywl7D1baooPXQZE9i0Xdw+Feq9Pe3GEa2+V4oVJG7AjIWxGihNM0n
FI4JWrjf2L6OQM/atHwtIMksoz1WDnHgNwZfsXGVXxtqGPBykKgKPEzTRrOibUG7yMxrHf61pXH3
9rqR4sjHK1VGIoJzVHEXoEdG9+fs7KZO7NF+caHid9Hb/T74YrsFTo5hqSYzwmYlMTjREgAWQKBt
0NYHLIH73twCxqNypJJWG7woPZqBYQfmaEIN4A9mE8o8yHma4S4Tt9B+w87q4Pij3HG8p1/eXUGl
rLQTAFByX0hQxkOJIVsCPzkOljiolot7pDN1703CV+e/oIHr5QOSJrb4JV1wtDtIIMt0xcYmstDS
AYrdAlMOHYL3Cyu+zncemXzNAHaAev6RlZJ9h9s/9JC4dbAqo+DyceghyLm42kTXiOZVHLIBUqpt
HCdLzQoMo/5ndKQVfN9MshdHn3/sXV8ht6SKli5z1RpIq6o9gV3OXCC6iYDvV5opkWaVh3r0wfRM
cNWmsmWKh6pXlzZFx6PkoSooj9ZjDrCZpFPjwrMfyvSP0+VMxQz10xyo9AdxkyZLlEA7j45Dti/z
X/WJopim7ANJKHqAmCuU5YJckJ4Y7hqwdbnVk4cUTf36IDUizhJ+/F3k81aVYzSgXL1aI6kFHd2z
LE+pfTZia/x05xCy2UCXobM73ZmFUCLJ5rjosvq3tH/kZQsyaQTw28elvMesDlSbRHT+mmERLZov
kCalkr2fHT7d+EzdLLBKLwB1aDRtNvPbiBFjGSp4KOeuAh9MKpkf+WoNjdLa99cCk1vvQmgYRjg4
A3XuWJ5Exk7bPzFKKP+NUtpVB7zDO/kY2np4afoir32JAH8nTJUePlcuChVQHL33+XPPuVybk+TW
0mxV8Hpc5/9s2i/wNPlfFyoHIRvTlR7HmIIwLT9KOrITJ15L1f+jlJYGKqk1uJ2h7IXW4v4IClHO
0zAMCKMMgPM+I+GTq+Nwq+QszltyGsH1P1kxqowUdVVVaBEvfbuNVhBNDPt81pmwXruYfr5cz1EP
G9iOwe4eyK24DLdqgOV48nowjFWvkI6ctWk14EmMhPAfz4zG+19xVImEOnzjOgw/8lOpXmp7YwvD
EJhViLEgL5s5IfpJuOvZp17NnjmcwyNno8uSeYgW+w1gmSYJBlGRf6A8BtBej993+M4cUGSL+9K8
+3tfMzSpE4sQprgPkAxGaeACh8ySIqqBbGAReVINGOEoczIRHzq+dQqrBw6evNQDoKSjiFtpbPOj
QNfvikagLoarV+bwU+GF2+NGPO2sHkT1I2z1tT2CMxDQ07bXDKcgrSzcP44ACEhM+yhZ2/zIYEWT
Muhyq6JEQuanHpjuKHeB4c3to8L4ebecsLudtIs9A1+KkafrKDCoWK/cE1BsMbCCfnOzEzq1Z8Yk
Bzwi4oD8YGqoy2yX9reJFwcX5BmuUlEFhDHTIL+A7oi3PNKw0j3Fna51PwvJHSpnReLrUsNM09t4
sGo7wtFuOKGna3smeg3/v7wMnaf5AJiNTqoRGI2RNLmHh/qu0gt8PcxxQlvhaYo15X00qbwCMeqx
jiokq5h2JS/jsEOF/yb2hPCFvFXoswXgmILxU700wn0KinUBINiAcy5xiZ2BgHXB4bKo0cyjwn6R
dRw0haotI2JGugjOXMUoGgiGY9XFPhATUuiRUNmEHqVWMU1CVOdmCjB0v/dFihL3ZBA2WpVHihJn
q0fji95g6Ywtt/z4s85iD+LnJGHDX63NQP0gOhn8pv0UFQYmQSiS+13CBy11O9o9a0fEIkiZef2Q
zVsejjEiYEw3bfhnlqtzqDkl0NhIdpJdWNvnpMxN5PO6DMHfzmYBi9hEgXDbsMWvKiDY1WNRaelm
yh2ZheNSMPXRkZi/tE1KbRHOM5uYxbZy4Ulg/U522ieYuetOBbMty0GgMDLoArive2VG0qHSqRgW
C+nq62j//OmKwlWnzPx+UcEcVyz5dfVUcGHp/Yc3Tt4Rae8fSExffd6kptRYC2fu47LtUFhpepqU
2xhDyUzq84uYcj4vzMpFW9/V0bFp4Jtq+U27aVXc5FOVqulGK3QvnpQLA0hgNN37UdsZhxhaH8H9
2yjyCwqYOJ+tAt2qiOspiZphWBadtEF6RYxQCtGxEPnhroBUgeZ0P83Y1gQmGAoyKn32n9Z3kvcY
Bh7EMpQmZwuCP8ocNKNrHOMOcZkxGHzlzIVhJhhhYyhS9LGOrheFhoEL6AxiTjgEoVrYvXjrp8YV
QOMrKqiIF+3bI+sH8/fckniROk/OP2c8+nm7QyvLBxUvzr8mrrygQQ5YBgZ/X7x1oy8euL2nSS1w
fTAn7z5otD/bV5ElygsVmErUsvFyTX0+nueHQgVZoRNtM7dHXS4+A42yHM3YmH0ALfjgHvbMn5z/
cRwWw2KbzvI0un4HPz2O8JR3q/NvltSCX1rGbRoQVxaiTo6rbsrYbVRJtlykjpzEr3uuO2X0H8q5
BxHTxpBeTrkh0eIwH8D3TqGuQUzTsq6kwSaQUucTr1bnNuoXdrs3p8vtPBFJXVcqqXWYT8NMJYCa
rRZd6XusLwi2yP85BEJA7pyY2v5wT8wD660XEigHmMA0+GafTivrdlqc1mUlIVG/n5zLIuCL4iWu
qqz8jct613k79DL79x8mR0Luo0JnDTQyrEIEw7QUxUFul13L2BGA1Nwjyzs4ItLH1FS4uZzkk5eE
J/f8OK9pdojBrJ/vQDQhEZl1LFmJaryowkOMGMYNuTJ3H5y4KDp38CpT2vNJV+/ufNr/Mi5v/82+
H5byuEo/5fH4pHqb6/YXnOo8hHoa4ZwtkO7vRVjO9FQiZ9ilzVc0cm9ZKSIfBuPfsOH2pg1Dq6mQ
ShXCOc1n7G2RcdyC24dkNacCRsNaIQ+lurfOQEiQUjjuSWsIDeWLbPQYO4uynxJVGq5FwgT1bAh+
lZcSStygA5J3mXINENEHJhB+Y2HPfSwDAlOM3x/MXuHXZYHoCM+i4Tq7z8lv4wY/99y01vpBfaXu
TvPiAmcmJ9e//JPTgGIe8jZOvulYHFrxt+pVR0xd7dh1/evb+4axfHqIAgzFkPtF/r/TaXIM9fkg
niBlQd4P0NOLMJsU/3T9JX6jiAb8kh225U3yKYhriYNPxJXZdmpcxq6PFpure0GhKxZgv4cHW+Sw
1UpvhY8/BrNWtAXZbDOXZcwOA7+lm0YwXemz0Xs7PucB7Kdv6FhaJkqcUZIdlwkPR1j8dr89MSzb
0rw9st3g4wrtfZHoR3NctrKiYhMeiSI5ifMprG9fFG1wwzFpTIQ3FicnMYv/dLWmDAGCu5pFfmJ8
Oy9tfTW5cwsn1d6zt12FtZwYHJ0P1fxG6wxEAg4a6dUiUO2/TtlFSUOTxJcZ05itvzfdlq3Xg+M+
Ib+VVa3leF7KQmjq4yiwOo69OVQ6aQgSGNT9C5bvqr+KMFCU1NlwhhZ+J7HXJKByNxBihopa8TlM
LGmHxleYVHsgwvO/HTGWsemd/bfXH3seybxEjNuqdQhBPRIB+jMSyToWOPgSJcXZLpEe0DWBz7hK
xCk6FYdgDyP2/5MzaRMw4ICodp7YY21an5CY9kbW+fmNdYRE0jk5GicVOmDwr5aiXeYpGhKOTT6k
CTyoopDeNFcf7zdMvmU6gaX+HmUyo/TIDMe0g+c8u8dNRitguc7C41quuo1VvIPIE9+cMVZPfWY0
+X1YdQ5MS/JGxzrtsGX44PckXMfl7yzCvGrU2yEAFQHKXl2yNYkMXyeetNRV8kP2q3r7zpuKuYYz
0dVIerfoHzMqcf2qHuoMH54L4uI2A9wSFHu4f9bhHqkOworLzIKKZLROcH8z3oBO0xKHNLF8tKL1
pAlqwgimYJcz1gRPrruTNoH1LI7D+j5Lzfi/wZAbtdC31eNP1HTEC/2zgYfwt1Bz1Vty7XD3MeA0
behkT4kAN54euozMqrdsjfQM2FZh5kkeT4cQoqVGyBxk6fFqQ8siQkke7i6KRDGAjRVzpLl32RJl
GdhsGrkgDobBd8Iw8KI+hYkX20HoM2+/L2wpYz4iaeoFqdtUfQrsA4jHwscWGZiP0xabHD6V0TLK
mh6W1JH6PGAZrNTbsTA6QYqgb8yVUpIQISTSFqYKZ/QsLrvwZ1QcXG56OK6Mi44igjUH7jlV4CFq
BE9JRg4JQZav5OuHxxu5/JxouWbpdNJm4Z4pxWbBZ9J+bXCvcwZb1X0tdapGCNxLgwvSjxhiRPW8
p1AOGUpejnFvqn1UaqW0Iw1a5ATwGFKjY4QvRUj8d4y9KCO9TQwD8mKrl2t743adBjs5bwCRv8X2
+mai6OUQHV3seN2v8WI1rXXxBPlgsaI/+J8OGu4zH6RFzvZN/CJzFFajuTfag3b61h3tMtqr36q6
dRsk7lqtG9pzoeOMWq6L1EmmP1tmD2ullGW8DRVKtpFTRtbNQmxuzZiQOWOMW1O80HK/EE3hBBr0
GvH/cJhlEa+OYMz6BC5MTQkOWEUvXVRC4e0uBtxk2g/7abjSH0hLb8QWxAftCoon1V0oB4nNgBua
YYx/U+87vJH/a8XW956+bJdLzimNiz2ADaceGaJaXBVraWa8HdJ32xrkMtCLL3slr5wQj1mPgQm2
P9ZE7Mo+qvyjGD5j0GI3nZslDETCqUCJCuIU+i8wJ8+R9zkRB8ZJMx0JKtuuenM2VxnQgZCpqXf3
0zRzcdAzq5COAsfced62OJPqJ2XEwujol2/mvJZ8z+PPY50LaBNe8vSw54Ny8OEmYxGAVSsEga8n
rao6MxTzD77//JH8d1WVFRN2YHFwRnldLGayVXopIp4c0gK0eApiVRYDpIjQ4y//I99FhzkHiE2H
QWuTM3GTAvUZ992Pq8VCzGCkRa/dNQ2DKa/tYx2XKUnWxarKgtYgWODKsvh0tFj8uz10W0p83rv5
jGpz9yCA9BcpGYmiW7MuxVXMF49uSJEx/egPLytSp17ks7KlBqrfOq91puUCsvCqd6ypYYlsdbTL
0SPEcDnkqydXBl/1fX+hMt3FUCNXi84hsZEf2vVOK2T8zs8Aya49gCsItOLGoKT1eUZQ0HSbtQt+
+hmxHpFTK2br755HOUCwM0a95ZnAjW51+WtQAOjkLHimny84HtnnTO/LozZdXxWirWMpwOsWyBLH
I6RROqLkkZ2LUBhFAd4z8/2f1tqe8NVcvdYgeJdJp6iczSVVBqldcn+9CxG8RdRs6FcleqA3u/oO
W2z5/2C8RTJLWBsGNyrP+GAHrnpL4iKMbrlhX/iWTzRvmEs596Yis4gIdjqmypH7umOtnnmA3Tqh
1BeWN6QzIk0Gqe2j1MWdU+MFzY1yGFeNC/1HosS/eMpRFNgGgVMFvEaXTesstvx5BSSkzluCC9kN
cFcXomi5e1S3w/db8VMCvRztpaHdDzYiymqIvboPvx56xv0+LPcTqXShYVXU130hjXV+wxpm1aM2
wA0cTrj3iFVlXTp9CBl8Tn0nZihEd3U1BiK/0DUFx2ZMNiZp5skjV++BmxC138pQmb2zGWaY2Sel
4/HGe+jT9TzZGAvvSZp12natYgeMnB7oESmCamrrb4+EgpfNSHaDkGgRHTqn4lViBWWZ/QyF3/er
PiCMiV5248mzgvuHK/Dw8ZWNxePv9uOm0cfXdKdtPGaEhDlgq5OxVtgU+BAdi9Eftyu7j9hI0h6F
vRV0K8qXxkUcSnBhOZabg9G/QxGBFlhyzUyWrFcyyFs9ElGsb1iTLnqi3HOeM7X5MEXOV3/XAuqN
SEJXV1eMYLXzH8xJ6XyLyHc2DcPR7Rx8R+UsAPwq2XmtuUqgFTkFEQRdJh3alhfX3IVQQy3sf5Ys
oPyWdf2a48eSeM81aGar2773crnBog4b+CtvonTK4NVCclAUpMbXQ2vCYhnGFXBwVulfm3793JM6
mnwa555GxaTzcVa0pFlKrAPriLSEZxA9q0Wfvhoa6im1O8E+ng9N6KBBVCIW04giFWZZ/S2oFT3M
mRzCgApsJLXl6dkJ/Or0y+E/rnqi9cC/WqwHF/TnpqwsYkbldoIuqyiPedv4+7RogUwTlHuh8vjl
+nAz5TVoUiapglVPb8ZCDLuzrjXc3Zheh7RYgSq1ofLmH9KmKg0/c5xdpIZeOvk0KEIKODD5R47r
WRqp26qHsq544s27hsJV03b3ETMo2h8UwvxLQHvIP/iFJ20oMfDcygX+0qPyH5S05+RD1fBxqk+G
D7U/ExFGSzthROjBGmBCacgd1MnD3zSSu2h4JsgNBHx1e2twYwf/WbOT97wfBqhHx6RiKQhXmmv9
EbaK89F6KNs7trqD0t639+ZyNKkmmhSMW/pMy8aGnTj5dvjAqstMFWhA1GvzhlUQMC1qhXUakv8g
gthotDPRt2gcGogVvrmGWQvzmBf8T4tUgqCFHZZOIkiffL8j3vg2dQ7gBwkMnM/oK3E/QaLT3J4/
KUcLHQ2RW6Qx6Hvgm2c+6ZXskaPHBtCGKxKfVLZhCIjOAWbmxTK7Yn6i/bLwf6A6CFylp0B87zHn
8BhcrN/03JCN5Q2k7r49IQ41mp1RAHCppNrjujEdGNR92r7YA7oVoc2bU89x/6aiT8aKbQRVgNtI
QWI5LesUHQs8va/S73Zf2tlL1I7snZgChP1yQjGvxKEJfnn8kUHAhzekgYLuSr8y+uVbQ1jwKiRB
FYLQzp+lU5qOwVAwtdd1kx76iRqZC/4EUizrjuAi/RR8U3YF6XXGwf0dszusFDWPo4Wi7cugdWVU
oh5MFGzR+yH3aC8Cik8X2U1vgoxxi8v8W1lOrpmn3B0+7LI5mhQt6ovruTrZXFz+P+6G5d7H0Bg0
e6njiC7IjPU7/E8gUufuC9XLWDbD9ovoCi0VlzmV5VaJFXB6+3S7e9Uy99L7EbaWgN2+xr7iBb14
5SQ5NbQLxSJU55OeHpu7bPkZP5RIzVZGa30YkGRYU6bXgUMUCA0X0lkIeYxmKyZLVbQtEsA0AcgZ
V4gNo7f5acyOxJKrMBVVFS19svTRXs2v49FSDSKbIXCZ33yTXAKyGrqshgsoDcQAGmf9dfSHffJ6
ZRo/+zJyGitm3chitPADKlBetKii1UYeMRJDd+Izj6M/O+c4aGeTrOQtuL+QbujYU/FQF+1hGG3g
/EU2pbtvcdie6pEa5zkb9VKb0a99s7ytQDYLl/QqXy7Vw4h+Uw6utngXH11Q/VFAAkC6Zayi8IYZ
Qvk5MhU0KD6ZnqNMlrT/V8IzPwTV1SwkFwRgMqaeKKvSEKceI1EV8n12Jof7kJRr5T57+xgcFvpG
pS8kWMlmFiaoPyi3uD3ao/KkukEfAXBZ9DoDJxOHr1mdgwvhKqibSvwF3vc+2F/zgo1HcaB4QdZL
fiToHIQ0VnpibDbD/bYFV71qYaXQ5Evvnc89iWo4YDpiDPWFl5Lh7jNoYuM8258//P1yfFEf+wEw
/FqliXK+d3EOcJhsm0zeHnipBYUjS2zkUqR/Nnrm7U+yMLYOkbH2BtwECHpfWLJY8VcOANLwmhKU
CwOTz3spVzuY876+UGClxc8gRidZ/Fdlkv3UNkPMVhCk3Jhheg1D6Imo0XTaHjrMEeB4tAX1LroI
cTv+fDKCLMEADqVpl2QABJMq63EXTAwNTDDML4b6LFfabn4+/wl36Z59rsBaavTV0vBC26lA+gc5
NJtk+q5Kjoo7P6L1tGfBooeR2r0d4spNRIzSwiLGrZfiSuDIFUJ7f67lY1IMBwArV7kxsBMuHBLB
o+N6abhRXhkBFvxQVWlzQm1zitG7f7+PUvSilXR6D29hDwlFcsRxgVeP0hr2+UqgbNYIeX7yUxM2
XGhZWlX74qeIWBhp69oS4NustHspiVGPWZCF5qSh3coOEvPEZChKNXpfg+Qjenm/qr6tuvRthY37
kzVHkSoGGLFzhYo955vqOnQ8pKwJjhXozqeJq5TT/+h5yU/uYikU84yapUWFppDBZZfE2okGU3AL
Nrwb12XCaxuSe43b6UYHgM4pdV4JqdG6R58WEuLJ8Qd7r5jojNVw0Dy+dQYoDuv9Jtl9SSrIufWj
lCVLJESWY+kS+4G3rscDUMfY6Luuc9Ribw0ap3XFTi0XZV+IqJfJrLH7aCMmNFPpianyINUqNbdn
zSMbydcrdPfRhwBrH1Q/zXymp/ZNK/6Fhd22YQtvv7ygLzaITURfButu89zo/ipZ9XKT1Dpc67XB
uAtAKZ+/rK92zu0lX4dx4yEIsXrsdH6BD9R/oxbRpXcjQOgxnLRMd/XKXlO6VOmTQQ2hCO9fMoly
uniHRCYO/3cEWzA/mrSQWcpyqwPcjE07Rvup/ogY93YwCVNCdMftbns7aQXnx25M4pv3KAsOPUqW
4kwG6CmCXfPQ4TlRD7VvsCB2aAGghnZsmh8/mPiEYZBXW/y7c8g5t3QuQANv6YZftGPGTMkRBMKh
r4t8ZUw2vciNhSOqeYOj5aNqHrKzjs4XkqcSey8td35qeU02aj4wJnBqZwfhEg/9+BGzn+0LrXr4
TCAUW0t2nKT82NqWN3mMnUTDLdiRN5aG8RRwK63zs38RtgxuVKorrj+8qdASbrBkKeL/VFJaHQG3
oQTo32pFjwHBPQ4KKe/+xzC3tf2V6lo9N0nAdK4l1IL/35Ba3ALf94ZbufEzbuErArH51bXcoQkR
RcvfsXMZphANSWY0VMg9klDw3//hij+3DhEXz56sEBvmMaWfNlLvS6N4VWDxZCgBKwoiVpDZlzbT
YFm/+cUfj5/zbMuHYOG2RQqDQgJr6kxHCAwdQDefC9OT49fK3ykp6dIkaz1IECDdMgibYRrZAClF
W4RMTPuXJPU/tQL63M+LQrXRdjPQpDIY+zzIX/5yTGw0oOezpHdU3rkGMX9Fpv3EfMtDYVOkpYXA
+Xg40FjTOX89XdLuKer18Og7mukagtLsQyV47XIa4rn1gDQ9TNIdiwf/DnSYo/Q9KxYBDw4KHXrd
2eEjVb+jk3ULg1p6H5uqee8C/dA44wdTyhB7sKT4EOJnKW1Jf8ISIdaJjxOBCopeKkSrlzvG+v2y
Hb7AwR9mI76tsYwDVbbaCKgDMJv49oYVJt8Hxm43N4FkJO+OvnRSxdJ1XMmD4R15twYCnSqMyYRR
mSc47lxT5dHYcxu8FGsa/iV85WKDjnweXdLXRRWe91GvRWQk2lEKKRnzBBgtSsiJwd9J04HxMOH1
vBuT5NDjCZeQ1cvyxJkF4Y3jEkYdhKUKm4rzTk8+Bo5OVvLAqrVEYgjkKg/daW8NrcQbPZ2JTcKs
osJYzGpIB49ki2IDpxuEowCjfKk4INaCZZ/GoJKeE09XddNp8K1TVo6cAV0jGuJp1svylaWepMl8
UEmQ7mnpRxydkK/o4GHSdMuD2C9fAuijp36IB3iZ+lCnfusYPDiaD3yBjvlq5DYdUgLCM//N0L/Z
/6jTFdUDoT41H/z5k6r/5Ku60NzGKRkxXVRwZZd2f0euwh2I/bVsZYPSsrENMd8sjY2Dwv7fRgwe
HsXv1YXMGS56DPrsYseIQlA5mabNkPHMkSTkZK1z84gipJHpVTY6p1Cd24lu2edaaaPo8aK9kyZB
EryHEGlKQ+FoZynw+aJNpuhjTFhhxOolTA1pvikUqz9e3lwRrYwMf5XtWwsDKiA3oqy31Mw5kcNK
a8psrdgipBvI/lyCvDWe00+gWL3uTdEQouZV54X7hTjQUyNNE6PP3hGYFFzggv3idCmNqxZSddR6
DgJttThEKanU4l5q4VW+rNbi7GFBbJkQUm+ViUa9jw+lCrSgCzAq1fheQPs0M93dghOkpNX89SlN
CxOX5sCIF5TQpff8cMrjf0m/Sywj5iucC8A7HeH1w+skl6LhXJjcWADzSaPeW8X2uARM4qH2unA5
VqjEaRTQucFjdq1P9ad7GCzoD5gklnHTjPEa4iW1wxtCh8IZ2XqIpbrNRaUgv8s3YfuXSczSw+4r
P6xx3U4Dn3OX16Pg/YKYcgJP/MG7+c9dnG5VSsukQ4iFSd+NcdyT5TojzkojlOtNnbGaaV9yKbbI
t2JiSShtaj8kOmrl3VIhopKH4RnE7Xgl39nhuxEo0cG32bEMiTjRtKLQmgxB/LbNTnyNxk5EUlxr
BNBK239brn9UpT3E4Vg0TEhBxP3kdUdyyVatXVQS6/txbopBX6an3Qt3ExMlBmXMgeAGpnO46d41
l2BSRmJXgOkL0e7YAoCgo26Q6dIv5PxWAzW5ycMIz0KhACbgxWobj5mPR/t7DHvGDCbONXUv1wWX
t2oHa+ZbhfASOzQJHrlRgBn2V3+rE0eIV8Dbp1Y/+crzJDLj2vdAxAaNKK4SQHapngvqduX9t09r
lmJG9wx6BVJpKoDOXr6xDTeRAlX7m3DxAQI9w3SPjgcCBLzzbyo9qDuGcJ4C9emt9st5tGN1z/c7
irQi5Pj+ju1UkUlnhq9yWhIqOdKOQF8pcUjlOEQfC4/nbSY+vLWcOxDww3MDZkvNjj+4ArMwNb4e
69WWMHCEWcm1/003sRsrHX1jQ8yl0iAlkk9lwHf6fizuyGqGbSkivkDNX6pfdoMEEDmoY75qBmGM
NXEIeosERkVKTaaISt9XlCaWdm2hg87H0D3Z8zmS4hkCqlvNzbQlQUNpkpzNtc0uftB9rsTasjMv
QNnxWVXZHHkQiKBrEAPYVZo17z/2esHAJkczzfZxA6ilONb6sRNGxrnG+ME7kHxdxeNmoT+W99SW
mWi0ERQbM/M65QRAzlGe58HzYcX9Qn2vnFEpHnLnFsdJYdwWVP3WFx2geMzALeuWPVq/ZJLr4AbK
GPfNOQ0qpugAHTRoiZJzDvkREq1sEjmY/j+NvSY/nyNNNbPtn1lHHhdDtbd7s7jfkndjK2cP42EQ
26mOXPu4r5Fnmj07P4ZU24KjPubXNzEyqDZJt5IJ1ydoLKaq1QDO/QHFgMQNcQ0kXoKfUkBZ83el
bcMHpug6Mv1x0Sl+f8ZwhoEAqO4TozpO6R6LMG9jNhhJUYW8a61LM+XPmyD35C/EuSQUb3Z38tx3
P4FLm+iu6Phpz+ifHL9eWfiNpvUfaLd/X8fFOSUrqJKoEWS9d/f+88MbgPZ6pUQ7oO/9gSgHy6xO
zDtAShricJ0uq3srVGtmFca3/W8DGp9xK9ku/0FxxsGusExI59qj+XLTzrqmRNrRsMJAk+BVw/l5
OVSF0e9FTpLuqT28ZwrPVNAd5gtR/ZjqHWa1A8/vK+3cA1CCszMiH2uldNPh/NQiYzbZCmiAJvUW
k/mVYzTfN97hVblPNKiV4dLqJiJWsN1tw1wsbkqRzkcJHN1CPUmGmTb/uTq/DrQGq8OQgqijuURr
Wb2T7moBcshJlO4kqBDB+iT9zgQ174kK9IQRfQ6ZzuAY26SQSzbHBAVoUVnX0Opjyzo6V8xzuQJI
iHVeY0GUoE90FpC3DbTIXjiqCKpJUZT2wMDFWKHBsIGcozXRj3/4R/7Q9UnpxiWhOg2hRzkicpfz
cbyy2+Xex/5Pqql0r2dbhQ+GmCezbWlZH912ivCEN1qmyEL3z5b60s/h48znOGYOw1gBBYzwNz3k
GE1hty/PNfQa1vnu/yVCLJGAdy9MP5V0bGXQ54QB6T3JWyrrNcL1BwhbnLcADrm821XQf0qVi3rt
l2PfTYZAPv2MNM7rALJf1QYG8uczvNXUWmkVZT7QpQTRHzqCjwtV+nrnJd2tpbHe6Pl3WHw2JvHF
tPf83+X5JXwYjEmHnFwM9MfN/8+xuf/5h2fyxOq8tZqWzuwzbg76bZcG38DlS2HosHHIgqTdfi8w
NW2fJ0x8bYj4OHLZuNEwR/y68wT4WvxbA6PzZUPnF2aMc4NLVt6BjioRUi0h8rwb4OlL2iKvaASR
mRN/E/kFK6sknEZ7O2i91zni6m0MV4My7AOJGDq7nuZTKbXDBeNMHVfKWwJc8ZPBpUJdpB2fpg8T
x/2DedfHPpS0O396xL2FSBdGlUnQigjrLxQKILLbuVFTJWN5bWeKHPjzQ9D9UVOEUPPoHZSJhsD0
XFajC5jvt8welk2ZkNCrVoBx63v/MVOGh5z8fUQEU6h0I2n9sRCEwQfpVSCCBuJNZuyB1LQSD25Y
/oaDfaSHmFdMeoy2tuCbS3/Go/Sq6jqJjH+bhTYjh2nqYot6r/u1/p60PuijpdaS/FLgBzp5QOkf
erUHbojPyP87x2ButKaQAWS4Jnnl8i0HVPm7bWvWUux1D3LrRsIG90w46WxPR5DGr7g7KOF2yhTm
zGv41B6GJa0Aq/mD5Z30kwNjD4OmamlYWAPjouBSej+Bz7649BmA39I9HrHTixfeRO10X/TCR1WO
GywP+Dp8kN0b4WlRzzIiSHvIJrf7tK6jqmSnfNRnpuHg29REbF+ZANAMAPM9/asX0klEkUdptyBh
9SAWirlp5oEDCXUJklJo+h9tD8/SKbkbk4Endwv237UgJpBki4ha7IVqouaVfgHZxSjtB8PvVcFP
QP4wzNuWLOgYhEcur2OzNdbru6PojTss5QVFgAsLJgQYexaik9qLDvXKvC0tfgVyXrqY3k//iX1x
Y3yeSrlSH1+CtBhgQAZwc9y5Ka7C3dvmbAgAU4EmE3a8QYkldcyqgwWxLw08xUCXEfEF2DsjdH1x
GUgkSEXY47jsn4h+TAlKkc0EAyjp/YNFglafckvJaLFQEWMOM+XjIDe20164vFfpjFWoQcn4fiB+
KxfsJ3+F7aKZCEDshHnEwrLPIGYPipp4WT5E+CqqyIeIKEgTKHTdKYNWh8zeH0FMD70IZc4ScM1Q
MFVZZVTLU6Id/WgfxuXEcn/tACWflUOONm6zpG0sjO/A9QOoqmx49TRcDCp5hsKxWzhfV5mhEJKc
WyS2tcS/h2/pyJmLziIboHEg1f/1TJDNTHOB80yAaLADKfv7dkv2Ryk/OQih7APJkqZP/poAgMBF
mxRewdTlF8wWPQf/eJsXIPY8EcGsKOOLtqlHWsbBBp2NSmW3BdAEZSp7EhmME7VHePuWeE9eLeJz
/RctejKJXCix7kDlvODVi1TtvplK7qLnh0xiL/ufAF0fGwgxxVYAxbXRIiz1s+8WFPa2DR6845i6
ayMFfsHT6i1w3h+jpIgy3qvjwpFHEe3HUdQdmdSoUpOdAE8WSpDeU0LBkLUqQCgHB1As7cfB0w+p
pU5HIJmrbtuCVU/mW8lP0Q4AYq8w1mup95TM0gazdxdMU6gtOWBcQum2W2EtjPu2ueehD6EBo0nz
0BK7lVlis1z1JYWvT4cTaQl+eaSeD+9JY97mZmtCe/c5GaEGoyYVIagZfevzR8G7tLqLFGOkKFXf
uK/ZzgV9Y1pzo/bvVod69yzKNYlUHj53zqz/SijJ11caATK1Ch1ULuAiMowy+54veTqW6t/Xrl+k
NAj+sABg9O3FVFFjDkHZ6vW1/JZEOuU0BoHNH4YSjcOPnNZ4lxkiw4EkMzsTlsO4xKu7Hch2Mg11
5bUiAnqSX/lCuPSk2u9jFVpTvdFMz72g4kWHQqekX7HuZ3bjAjpvW4CFfVhFrcmAsC0MOejhqZuq
FwqCHnehq4/EwdlZk4+rnKMcPqw9I4U+3PNRp3Irzl8ibbbXIM+IAc0DXoUiPu2xAxR2OCCRJxjt
5/UiKFGK4reX5mu/yFmrXLfAc0lAbfykWXXHT1vInlR687IoU02KFDjj+xVtStMsCSFP8CMI2SJj
bGAPyB0ka9lHHzt5/+PrjxriOzg+DoVHZq7r2+VhDLfli/4QPzEFgf84Qhw2zIi7D1tEl8cAwijX
dJS0zVdBUp14UJjyC+4NQtJKitM68sARavwaCEmEX3e4zAlEmyBi/plZBwBgglW9ksGo0YeCR6ia
gowrnO4YuCf7OTIyhktMWLoa7sXitBE3wTm9t+R8Io7MLaueNhGiWeE+JtE1KjHXitVjjbiLiAme
KzA1JdkHA9iZqWO00oenpW0DqUo/5RTpRF9R788pkJyvChDz/M8ZuhiPwH1y/Tcaf0RlXYiTXMll
VM2dhFhaXJF3FdFw6o3prLOYcccxanC8zUDDIU0JDQ1x6vPW9XOJNVjCIpuitqDVbezcUQnA0oSV
VRDM+5D7+bRtnbzdWPuF+MUiglarfLqHx+5q1FuzdFdSQjjiT9zDYmv2ktPf4+gOJHb5LMfdHVgl
mbY/Vp/2powk/SHfVwnFqK6O7VEeE40zRKSWc/YTCPZX+ixIHNnR7PMSl7gY9+DrmTXIhJXUB70L
Hhe2L6W/63BbU+6SzdkQGs8tgYuLLJgDcrMxLanWX+Y2AS3o1zrFuutouEU/HkKn7aUop2nDBZ+2
teHEnAXQVmlJ3ZzNAz/OCDZeYPRhCgty1kzDHzhz+0eUbSxkONz9Ot9+1NYf0b7vmwdlabsB5Syk
d529rzS66umzWPi+GIfXhIrWBneisdyxDZhFMRT86x5Jc6Uf0h9QJ29ooWuhPaueCBc76QxZy6l/
bF8fOMDdp7cvzgVvpMMgq88LfehKCdSMGceh9cN2vyBjj7Vd0HYF6lzXAD8M/+Ibg3o1qoiPDgEn
gAEdxeiLg0hV99fCyNJq5ejC0Cx76cqiEYgXG2busnSyDsBTRQXdGum8Ecyy3RFpKN2OiA3rTPEz
Gyr2+8OQnbaEmaveRT2CKOq4konqGMQQ/YljRjjkqpKLfH854I1Ic7Yhx1Gv9CPCrNouU2zJr4CW
r1l7zIcyPhShIvy2OWM8CdEN8moc8gXhcVwmFKln53A+JzgtWDQW9cXWsV6FTdrBHfn0uuf838U0
TuteG10rDJV17etlU5qjZhSoOkN4sjkHpe1ZiQJDKvnx6ktr+BSNz3UWYjI/V38Ijk8qJSSyyfVA
/q/cJ6syfkxfkT9MxM3l9nEFqNx4BDjIi1b9/OIY1qpmMkpLTzZxdUVEMFFj2EYQs3EIYQUb4rfo
N1z/IbeqbrVe8AcibbYXWy8OpRa5sf6nqBbBrRe529Yd8hEuXwwQXr7I76FmRx+9NsZKi343fmWY
zYcK5TG7LBdHY6AxN50InNwsmXkhSEdmh7ksSZEzzfCWRhJioV+aKCHZobLwWtl1t60sU3tEmIl4
Mt0V3OIVEYNlhe2W9IfEe/SobijEWpEnl2i9RuAuRtLUoFXfjkkrM3ZPSsy8l/PRnYQojW6Pt/gl
WfCqpKTTOWcZW6rkvbr1NSV5Otxwvx998k/Gat0jcaRQdymlMo4ozrOQaqcxB+u7gqUh6yA6D3M7
FJ1BHBA7bRi8V1epQxeB7HRUbnlGUBTAvO0TdBQASMkPCJFYGjty0SDGuqt0Ai4azEVdFDAu6ITq
KSz0jVTbTDVBdXFriDI6BU+RdJsGRMcS8GXQYufXrh7C836zJQ7uUtnEq2S/GGmCquixcPpDkvRz
PHM4zpq/Ljo2R6BdWXndEDb5u8QvGws6l+WXG2VU2kRPKDf3JAeZTCB2ayz7yEx8T/HV85bXHMva
rZ1nC4xBMxTEyltndJ9zZgIrx/tsbi860whsPRh0QcqyIeM7a9khD0A/R5DwuJWhfpiOz5OZmORs
j3MSfYhTyQKtZrovRr76+nqua2lX1tYOf8Wk4ugymzU5j/WYCWEd7hMk/LA1rmcvh0Bn0y99aDpd
Wp1FO0nxAJuErYwRoKI/14i74/xWggG+805VHAfonk+VY73NP3Cbbmfyysi+6wKvMIqtWrNPDmc3
2YxGup2r7nrU99N+MAmNEeveH+xtB+BKPq94Ols2pkwdeVbruZ9Wd1UMBOQdjUrejkPK6xS6I8zO
gTtxXnocjkyOpSrjuviSPstBnToKRvLk2aLYxqyPHu9rLsW0H9D6mmne9bUM5IrtWZFFSOhfLFbd
AoCaIygPeP24nD8fR0XH7GN7ncp4Qd7WVXR/Ga2CISPQxhEqnMx9oQHHFQQ737d9VuzS5fzDiibX
SWNH5a2QVZurB7NYBPiT1emkmelcQWcJa0J5vmZdRoBPKzCT46tTxSOwJ548KMys3BenmklHEkGE
NWMIAEJkrHsgbVaBkaNYchahbHr6FpMS0U9huZcMcbpUI1pPbMDUxU9utiLp/wajNHLh2mppNWxk
ZmeevuP5GGoXqjh4YaB4dM8oonpKGR1hcKPO8Un80FBHuvpkGkhudmIVpPdGBxettPpnxvVgQs1N
juXSZq4KmVN0Fa7yKVcIcfxDs0yGFDVNK1k/nc/pdmdrqyDls5OxaKlORVwBVkHYoZ2xw1yW/n1U
6s8jGCFsNF6+4XVOtEZGYCsfLi6cr/uup/slLNKMkLFzgiSwk4RVoVsu9WP0aVLGxWr0ZSnyZIs+
2Raj5O2TfQLZiMTpM/VnkwhxEcW6BXvaudY3d06kgjUUKh1Cg45QRs68ZpPjVjOIn42yoO64S3ok
i//cEt9cG/wNB8rSIOiWX6ptSbsODejyq8+aZPmbuchK70PQzqSoQmPYKqJ4jeXb6Idex19ULpbd
WN2MZNSpwY6nfHYLzDFgv1ToDqJOLD2mOT3AJbOybsRbnrSm7VP7CWsfR1Q7MVACkTZQtzfsQWkI
aWWaz4XkLoO29Ue8Nd3qJm/aGqVLFOZykI7uJPm9fSu59IXb+i9+Z0BAXMlBP4NG4YgsNldeS21m
/w0FGfzTkqpNaPGlEk76e9c6HmPqPRAnLm0eG5QDhopEcPdziYt+AAuxLLjRttBuD8KRCPUX/oEL
9FAK58PTHjaXvaoAmZU8OymtNlIP2RP6PtM2yYbBdoOJwtrElP/JijtgobYpStN6kE33/yP7GHBL
QpbWKiBX2VhhkkZkVxXpaN3zdc2qd8uWVOaH0TCa/ON6zvllUhgYRVpH97OBp5pDfM5yTWF401el
YmKHJvMy4dY+/SbR0MsrNVaNzN8M+FSDBVaK9JbJrgUSfwD6BaRhJqzOcXKspDyfqi7q4fI7OLTY
dPyJVi92UGY/qg9Tq6QnmkbJZtcK1vlyZm8cbtjstUujnz5l23V470kb/tJhKpP+jTqSOiXBZn1j
/lH9MylOx0OTaj/KXnX9/4l+Fc2JwmG3o4/2Q0YjKnmS0etAS9qXAKL258RV4DXr8W1SlXvxeZu9
OfLiS0WiMYycV9jlOMS/jKfuKQhPPNigqDnA8sb4wAvj9jfhkYyqg2b9hIeXyv2cTil0usIjBCy+
CkReQxD/FQjQfGcG0HkQYdPUd3NivpFoykugioAOnaXPbPkNgQ7i6DavD/xUPPcTW6EjU4iKHclA
2TlcJKsTkP5k0LafJFUTRGcWY+K7EsB+O9cjHJM3ikl4eIufxDkC9ypcXT9ILPtSoCHNgUQAU0zg
nZK/wew2vx1TAFh9tuHcukaozrdvRg3HlTtcQ9zRUmZIHntpHGmRowqz6R1HhA/Awh0cVC0gwLyg
94CG4ce91M3WgBHx0Tbnit97Y5DqPmhgYY0SrJLDhkpoIaN8nKPJ1wYuCWemwQcKRsIVEnWmJaV+
29jVkhbo9cbMoaxEPTXW+Im/dXZex4ulYl2tqmoox7e9SzKZtORNYpMj5B9G64eoc/Cy6TXQK7bN
78S4EsbXVFkdoZe2oO0tKlk7VejlazM5/0oKifLal/5ZDtdbTdhrJcnYSkDL9Q5BkluEB+y/jyRH
/aZ3T3fyOcnNMylM8HSeSnCoY9iNtQVerSwxK2EUD85XT1NWq2JCO+/5tDyu6NZdANqGx/9ah1NO
HONT631SvWQLN6v+gbGJUPJsCoATp/KXcEpI9HSl65SxjWq66ck55wHYPH3b0cTaJYO5YIZNLTPf
SLXsvIe/xLHyXdFxTmQQNa5QBWbnwZIWIj1f7IMQ+KlBqukq0F8YKOGGpd4rCsWgv7KehR59/4NB
K9x5M55eCHyyf0NMFzawcNAkXbAdgul9TUwuvn5FZAAlXtfiL1iz2mKfrYw5n6W2oGXhPluuhPj5
4ak8rR2rH92PQY7P2O++n10wn0SsiwvgnOcfoJPw1jr86FddesWCW2q6mLXT4aFSqT2qqbn8tQM+
UVEvKgREppoOKXxtRsGKfJOrc6EXs4dEauc/H1GQKZ5qgBcKyN0XLVsZw0Wbyl3duHQRpJigHICh
Fkub+tupnL7W5LODugFmVxwA2/QmtJVm9SWOQ1TOwDHtA8vMfFs75daoTuU70c/ZU3tnNzTiTdW2
L4EZDyCWxoCyFYTDjO3oNcDgnh3P/D4b1f1KJ/si9OPJim0G5paB5UOw4VWmcir66uvT1KpN7Rxy
jRxmwQhiIN+8gFz4Mv15wyYLX17fxso7UQRgWibB4yDOxGQ7dWqQpnnE4hJ9wlNjwBRoPmjPKFRr
WJpIu7mlGt9Nxqv5Gwgu+k+veiWq0xFG1gjAznBsrbUrM4TbIMBsxtpoklWozMy3X4f5sOGdqbPM
Qx8TEqYAxBf8RTS/K6DakyCsrnS/tL7zzVVJ/zZQGjy/OQ95IbNtiCG576o5EEjyTRHokxYkJZWH
N5mI1Y40JwRTxCLng6f/FNzexzKJWa8czDh033I2Lzow4cR8Fyzfl9Eluxx4UvS94Keqs8qK20R+
0SbaxPRxb+SO6S2CLk3KRFR61B6xGPB9i0pAsRC+5JbWNvLIeiEnQds46u2VajMz2WvGufALsYeW
JMvoTknaRQNk2TTwcK/EC6P0Iwu6lnnNI70Nbz9ni0QVMZpm64h4WA3AatB+K+XbQEXvSO5OR5j0
O/P0l1/iEfmbPsAP/+ICTn+UNs5rDcKrcpqrgvLgVn524kbnXQ/s5R8wg8DK4zqQQSzpFOnzP2nf
og02Vfa9SlGoOrU4TQcxoBkyZqRG/aUj4YbBlwxTkYlD8ina2Rwo2XP7k1N4Hxo8aJt6El9I4nRr
9CucGfInrjoDMXIsPa+wrUIgLYB8xk46158d0MRxr5bAUl+2HtSFXosb7hHtG45k1OxkCVDZTFo1
/ki6Vwps+GDjsVYNPuBLyR5s5uSeyHPO+WvJS7Cyar7CmUxOGsEnQ/vfUftC7BwUjeLn4fisDBRB
V/GpWEGmvBl+SZ4n2yocHcsyHexRT4BhsryEAVPwFglo01Rv7RMb7ZBhF3gbVotrxzfyEU8QvrVg
M0yiX+bAN59QK6m9KZVmYBQNXC4chTnDQ8UvpGEsSef9VkBjxzlrhEWepLmJtJLaVdUDJ07cpnR2
zLsEFv1NZWVbAkKdpwjmYmUr8KgNLaFVlKB36q/SNZNMGOAVZkAGkjKeswdhFdC/UGB988vAD708
9EWgXKnMdGAjdcqjU3XSsq105ZD3LiCtk8ZhO6oZIcoPC7YIGCkex4clMYQtVHd6ay9BRNK+UHfI
r8CQjdlVgWbqNyf5drIruM0grT1v6jagOijEyKrvbEkpRGt2LyCYNSJqzvEJPlFuRwskRFuympsk
Dg6BXWPQMDg9ldlXtynH2XvbWoYUXk3lwIurVxdZgy3Hviy7Je0Cpb8dvB0a3ZicriPBpS7Pjj2M
EA+sripSrvid2rwVtrYt+TRZPcU7iboIxsoxfzBP6ZT8j5nHZd4H/bVl17V9l+pgZoe8fSF4k6SA
VxP4S0hDyhjozr3oJi6QSRSBmteP+lSRmjOHxoW0u66XA4piXefGMgbqz0lX+g/trNBwNze8+zP8
VbSzChMWpob7Hk3IeZbymzAeMpseZxrTWf4mmXZHTvaC0OJRasaKOCNm1fYUqzernakNPVs3djnF
BMR2A56ge6DOHCkkrMSQFMHorTnibktAuGKUgPo3G7zXwRYOUR2kfvQBup1sKPhpmMBPfelws1hs
eNeObCUvboqAPwqQjDNxi5UcSRuMqNDIdWig6/s2dEJb+uW8/XWPP+ZxLJ9fTzxn2T+dtmhQmnnX
CPYR3p4G4JGbrRfpIz9taYoD1VX+lWlAPvMyRmpfvRvdzgLO5ADyD5vm4WyB66yR1voaoA7E0ilg
1h4DdzujlkZxzB6hRRiYDZ1aQsZk3yONUWlnH1XkkTQhQHBbEbAaZFKfWt4TealGRZNSinbqLkB0
r3EBIs65p4fsD9+llfyzBpTHz1CBxWzn423t8PPnb8PZgWsFTY9dm5bLUx74MyyETXm0WK33URVl
e5hUC0qUeYxtg2DT+UK3x8MwZMZwDYPDHTbpIN2jxKnYYw7z/MYoVlwv8kouV2Gq27yn07NHUAqY
a9pwAVcAFXOZ5yfMTYJV9SQSGmGqxJalfqTJK9nIJbbIrJwt8OjABnbNIXJyyb+OOUvUh6uO1a4A
P3bj6LofXOUBD2uD9zsG11MeX9QFxfDqedcVkog0/eOesiBQVWxOojZ/UzLHw/zLXR+2q/ws+k7o
r1wAZjwUyZLPRzr9lAUTtbiSkAzUW63A3iv7jG9Au5ABEqttn/vtS31Mn4g8WboAN3Cx9s6ASusf
5+EF3zY/jg1ZVGqYgFy1U1Qn0LidCoJMr1c7vo3BQVQegoarbyKdTzmW29PRlQPpjqS/arHnVHzR
WDYARBOsnulX7DRof0UdGL37xq9EOj0OFaUCMZoCpuFHXSF8RYvLOnKXgvNNlt9ivMYGmZiHgeMA
3L3a+QKgFsXItIe+fcTT19R3a9Bk9GimUM0+OAvo/zLuyi/btNrOOywZT7GdTC6g+McEkUEYxTta
d3AH5Bu9YtG9dT/6kh7A6E6lNfIAhjyg7Gbqjg3LNMb0loa4nLABYga4LSTKPrpm/Z4k2VtfXKtV
8H/py8XX3nRrPf0WO/Rsvo4WFeQJZinICf6zhcH+YzMpQBLWJ62cQW3ZEWnEDNEFU7DlUcVYme5Q
IOJdVxxNoWtSCizr7rgazxZLUpxzx8jGCuL0Td0q5PlKcz/XYWHRx+Po6Pg57XFN8GV0vb8KXvFc
nbe3e8LNY3Gohd2XOD6UTVqAyBj4eJ7uj3gROncs8fkezVY3W458cz69aOUJmMr1pJi3lGlHnm03
VqUHugYFQ/83xl97XFVArf9gx9vomjReyLonhBnHBGBJ1xXJ7xJSYQqkldusyxvBeVwQ1R8d/17c
BIqDuZO9MzLwZDc0iOZjCSD2B4q4rqvebQJXJAvKMQbVzGKJG78aOCUbijzMwzl+oHlujupEheMT
21f6hbza57klc/3mG91xyK0ppFmdeCX5tf9Rnru7gWsCY0PK59WEeMCVKFtCom5Uo3HcI2J9q6nw
jigSIzHwJcJ3gzyHuImocH4mH/XoB53VKPmOD8G0tVqFupexyUm0omh6T17KqDLdnszUq/0EDNDH
1QQzMSceSBCSkDvBp0oR9mg1tWNoPsplaHo5SnPfycisRtaRVd6toMRwRhsG7Ve1cu+OAz8+hRrV
HLaleaqjXcyX0LUcH2RmWasdUinKv0EAiiT57bUQS0IECV/gK/Ker5CUlkfdQa8Tqb+rBz0rXAtJ
ZuNunzVBIHJ9W5qu+iWhugYSYlEndQalhze0rvCw3M/VLsJs64+qtCyMXmpGiU9b4DO2tbF/WC2n
TyrqUi0u8ZCFelSNR6IeqSdYUK1R3c7Se5hmJn1b2UFS+Ru8Mvt1AdFaoMlc/27gBH0Qb72Cz9T1
gVnGnFvMiLnhD7qytuPIhevCg9pwEogx93H+tzCH0Esl8q3tkxWgXInN+FHPBrkztC1+bCQLLgfs
TtXGXDzPoKJRb9hDWmd9781516ZuBaDU1YgGotlOXie8z+MK5nenHfAjwZOz1cUgssWSiPnOgI2R
S7kqBMWfP6tcgg5i/gtL6AHaecXeyOPn+cJ5502FvDXI9aSlelViGpcujeANWRi3iKu+Cn0UkUPx
hm8tSisMkiESOBPq2Js0qClwAJ2+0eMj2gcP2ESAg4fc3Mb3+HAN7bh3JYqifVw951FDfQxYrvLb
VSNgkPBdEWYW2tL4E4toZdi5niLpkznsLs6t8ze/KtqmfNZj77HM3Xf/v4KjXYyDEigcwlA/H4SI
vI5k2L2+ZgiJ3saRg6plRnX40N8aGDeZCDagJBWTKB+dlfIxr0Xaidtxe0Nl0DMoQyFWNK01CWwk
fdCVi//sYooMPMLpHUIa3BNcF8nwp7eDGGUjY5XaowolmhkebfVl6vb7IXYjB50LBSprdQJp2Q8g
G2OHnz+QpRaiDdNfCJOak6pnjTraIDiVqbmz+FXssRG/o/Da6x3W1VR3Rn/YtxrJsXaSTPsit9SP
aHIpTLi2ucKfsh2QcmoZSwhYAvATj16PIsnWP8Y5c2yNRYvw/grJ7ehHJ5Njb65NZyntsOrMMZf4
13eH3WkRpj9mW/x0fdcj7SUKQdopmDyBMMliFNsBabRjuKQQaFVU2BV1Hyvas0mMTc/X3GNZj9MH
l3QfIoce9ZuxbBJdXILHSiG4IEV5XZ7WRl6IknMpgwyQgc+EAM7vNIt4biT+j/AlKvDd1xWJ2u31
gG+Sp3+5rgMP5D40BGPUKcQEzBl5v+S2aOk472o5nLEQzSe1afLEFQPOMkowor+xuV7oXX7dcB/M
Jm6g+ArskI2v4/o/DB+EO9sLALwMYysjTiFL610/YFrv42ih3u+fzEhQ0TjkGm6fZAmekrYIx6RL
Tqpedu2A49Kz11ABBL777v3JfNcHKHK5+6P6M1qFwVf7uR/cx2RtSDscY+wqpJkVocwkgI2oQ9J5
wJLiY4M9QA9H8bM2BttNfS/HU9PMOO6XotFDFXO2rxAmt2jtiJ/n6g1YEgFJmmaHFWNByerZl+0t
+EpsiZOwAsTxhvENSJGk1604Lvol6P+b0SLcKcMvXhnJB0dBbZTGCbb5+dLJKgZ2zNlScu2pybw7
7d+jhhbWko7bm6py89Wn25proY6cE2xCbzbX1XWjG9GbxAUWeWK/9XDqkDRt1T6hLXIi59pxsvHw
xHwri3GuQUC/f0wE4g7X4Poqac4lhxyvqtZvDL/eRLhmDobIR3qfL5hvTr5bLEUH58CSgDRVEnnj
xXOuRl9/jZEO+BbLtJSr/hpmfuQLRJcxQNlpGb/KfM+0O7MALlieGRubVXsPaBMhBdJP8+jhfZnX
q69QGWiFWQ95G0a54zYeG8HzLfMiVbl533uJH/AWNzLf3L+sAcy/T+2nzongaT97oWWzdvDaZOAh
ePnyq9i+T+0JXnSnSk4C4DBUNpwFAXZXW+hr6KSR2xmdAtgFkG9vTPTiyHGtFcEpLC4HDLU/OvNx
d9iiJRoDNjNryn4nuQwLNOb4LPOxxHfUKZX5wgt4DgSKh+X5/6m16BZC7/PGejsnLlhYopDGritJ
Z6nS0oJ6eW8B2938sjbnNpuaF1ecaqKDxenNDRekWvODo8rcxX43vZYMac74WzNp2m+eFngho4MT
jyF4VWNOWL1VEL4amOX9DRQ00EFaRdq5EyjJKuk3Fuyybrp0fWsx82HRnhLz4eVBq/EXgwkpPh2+
OTXE9UaDvwQJu0Au5D5oujReAJ3Qasl8BzTQVCknHfv9Bis3TJO4QCU716giizUmhVCGoKS9d2zZ
aNd9qXSEWffVcxegj7Cxe7+Sn2ZC+3sxeWJ9fKUWUHHzi3STY07uH+D/9ac+4ag99/5JOR3cUMQT
lGzrND5u6npKS8DVZWVfOXXi9mJZP3KKgOcY3VvyU9SjC74kKKJ3P09OdMQEhVN7iz4HjbGVmLga
3GubPtVAaJXzR0q6IIagNPX7x2K4epPbR+fWTCrztdRvG2MZqRetTmpW0pUALzYlZ49u5f2F5d0K
/BUCYkZxhqjstsV40NtIh3CBaaO7aY5J7z7kLLCJib/uKLbAFbrXW9DyU3d3X0Du2JveCuiFPyTJ
d85GHT0U1XsEVx57D4iGNM3AlSLvBNr2ryyBTkTQnTixbzfrafaMHMPRcgkgr1y0OoOl49jlliXo
nHzFNfSwHxNZoCrJFnHdCBqJ4bFBDc5rzDPuABmKv6zCt7Uasck4HFyHieRClSGQU3eu2/5RV4kB
Bva4nlE+Fa/g2VdIYcu5vdOpG0KA9pznDhvfeR9ai1eMbZsvd7FseiI/hk/vZBAceuXKLlIWQayI
cIOYK/KQ/zudxHKAJ6eQVeJK140VPvTkw9ghw6E5E0LO09AAvFsZ7auyohA/Qf7LjhzzWVTJbG1d
hyaCoCW8X5G1NIiMKKnI2x0EUK+NAsAJN9Ks1mR2osvkjc9fX4HowhZ5CNcGImOkiJOZc2U17bR4
M5TP2pZHPRMIB2y4CuMsXo5s+el0otM+5ylzCGMcvOVL15PBVoifUqaSW94/316Ql+HHQAuvjX+W
bRSx/xGQ46WB5VTgZEjqyxEl/vKA4OHE+tVDuwj9Bl078KfyOgwzl/xSRpfSGNHyEw7LN7wTioo7
n0bVKJ6LWkZl8RJ61RNAp5uO6H8/fisGUrP+CMAdZBZ/sdNA6sfYBdLsXW7dvEaDtgnnJSSUAe4u
CGvfe/eP7GpHAb2z5Kd/HMLjHgn7BQqVDrgxv5PFnmHvmOxrExhQqgCA2LBjkwtObktdWgyUwcfD
eKaSssCrrKyiAdDg6tqPSTaJIqI0Cr/hr0l5NIQPIP7yUvai6ss6u1Zm7shFKIOd8PHI368Fkz+P
bew4FyUIWENHhyZe4HoHcKUHU75fb1WwjCgr7OrdF7s8y7Xw8goPqlfxTyrtYuy0RtKFl7YrKMgA
V75tuvTQDVafhFTtQsDyj4IzvFc9uDGfjsx3ZnZuZVYIqJRtDdehjTg1eA0hfvVz/HEwku9tiGVA
1FQITODdkWuUMzdEy09/SvmDq82UH8YISgmC2vi6CBcphseUsMOUzTGCYsB2KRTbnkiScMVsREug
mTeuy4pW2SoEZQ+tyjbqYEqxberFAkGWkp5pNf8wmfQ1hVl8taIYGpklDdbW3gKCR+p3+zJ11eqq
wbW2CwCEOXO4SQ1W1dkQkjO2aXXVgyPMKDNQ/YkE2tLWmZUOghuAgKqfGyLSLsFzeFykNd9z2/90
jbwAQU0/QNuR/OTPQ3+6qDOlMcuBDEDgVxfQG73ZaEWHvz4Q77nL7+/uEJ9S3ZJHSdSIF6w6690Q
vdK9tnVvP53ZuTqkDA58Qj1DNZ2ozzUA62dddIwcVV2/7b3RjAac5NPgk+ghma45LIvDx2sNH0lR
QQqDlnWkP9VuKaNS8qsYuxRiwY2iCCvMwNi3NgKy5HxW0ilMMMRjT59Tx4z89/jD4Df5EH7x8Ty6
vSTcoZwk9mq84RRe4tN5Tvtt9PGJFuXQONBZBnU+OEOGkZTTMEhAV7CjtZDFOnRDLenm4J/RdMr0
s1QVbEwXIXOVMuL8BERVmdULTYR4nPyrGp4rN3U9isoj4tIYFOxzaVUMXnurGX6btBm6S+Bgi2FJ
enXd6QDyF6w2oygoiOVJOWR0RwSFSKOyFB9MOnoNwn3qh9rgUb/483hasyKIQrsKPEyZsF1lg6HA
LB/QvOVjRo9h7MgY7ENcVrBbV74wVLPjU8+zug2Kd/JFKQuXLTrXY8+jNDVmwAwqj1dRZ7eBb0P/
UYQD8UVu7x5M++vElocz4B6ad3M1SvwXOzKgfpRGB8hzhvxNDZvzkon2iV4jWvEJ/ziiQrMKPyoP
qIRtXVETIjTJJmCkfKTuObTaaKp44s9Mkeai6KKOCQ/miVwtxjPJDlmf/QZvXzwOrCO+YtH25Af2
Wr5v0XllYmvnBbCN2tekg94fFL8rqXuJRx6ru0B+IKG5kRr5Dx+PTz/t+kNps2zdSPig0Hb8hfex
2HGuooAa39OSpj4QgSZG24Ob8EB27N2KFcO7+hOKB/IaTfbAO+uzAsZ90nlfJnNTvYAJTxm70nst
cGcXjw1qPPlAFm2FzeueXYb7WlLQieDTmPYoYrU5cxCQm148eG26vmkPLAyPtrQom/U1Nnvii24B
QkxoPHq/Xkg2ced4ICImn954QKAHsVFuwNrECTCwqzdGKxAIohAcgIk9L6JwLamnuNPmyku+Rt4F
VzNjpVVpvhn0ulCFh7ac3Xb7dnwVioixbBAYe2hrdY+W6yqTrGSiPPxE+fdBpX3n4rxXuOmfEChp
OWHckimrOvJP6tJ5q6A6+pVvepNNHBtPUgZ0Yc4GkzpDaTeGn4zDTY2Ey3a0v4lDTyXyYiZF1/5E
aW5BJyxdbUjeSk8whLbabaYYLajOXmQH2U/YogLiGc3h8tTrQxZ08vYbg/1xr6H+K02iRdirR4W2
plV59g57brV5bnWq72hjK7z1ck1sqeWYqpAB5Z9YZRVmoC1+3P5g54N8g0Zcq+FmrGF+tq1PGewd
Z7l2gILU5vhszd9JAhceuG+dnfJOGQTD2H85tjC1JBbJaOFcl2cxZbJ7ij5Eh+g46O3/OTAGfMqr
Jz/vKlYJhb9oS/L7iPlQNt0jTSBFNMblqG2fe7RRZZM+mNmKlZKhkCIOYPooN8DWtim0/K+gCM1N
Aa5GdufzZyOPwwobuosCLZIFHqv+lo9MrGd1SUM2gxaJq09C7X1JQz864FlSOo8JVvhb8ixVU3ZZ
j4g0h9MLOuk5xPtfqlFyF+xP1g7W9MwDuDPFOsA2haisrxZrDtx96pVODYfrhYTLKbOeLkHm53ir
8pWmuu3edhRUbm8s2fjaBusVoB0oX5waepreGjXLm+L9nlchmP1DfRvNeIfrO++yU0I5Ly6DI/vI
ybp4p8FZV+OkaRB+u99JzH5h6MJxH7kZtjYJaSeAp8CIZoZW5clH8t70BbnXxL4gfKtUbXgUWHvl
b/bQQFXSe62R8UYuXGO6nhJsY8EeY9PxcJXecNt/JyxYDLNrOeCHDtZs8IfsmMQ9unLxRVx060U0
8JT6CPZLqzbFJTvNcIe8+o1B5GmZwt17Vcl1YUcisn/iqlTJmo1BCFsr04/0HFVgGUfi+x2k4kQx
01EoXAipJQ6S8fixCtFTnlQi3Bz97DpymuRZZR4bG6vL1OtDJ9zou3duhKCkgZBLDmiNnttWRyM6
ZKDaMmqKR7UzRI0DFDAOEVM+DJzeoy9G8c/OPHZA3E4rIvwpFjufuOrvrOOs097OdbYOpf3n49zb
sUjRIofLr5IDy0InBfW9qzYOZlP4z4i2h710+PAYQLYFnkQVHlcCFML0X4xwnpFm5IxSpvZ/zaVc
OA6wU+Uf9pLHeT+UAGGZorxv/5yX4LSGYoju/1ZDy7dHJnzIpLC89S0+T+WSSNpE+J+hHilbd2AS
HiufLrliCffHOJFBTSpDXCwBRlgCWKvKtIF60tqB3xUJdBnvDJuab728J8DHoDL4XZwlDw7kRPsy
bGoyFu2AOzTjuKSsgO23ZposkHwC70jT4QDceTEk6Q/WYSDY1N08nlbMwm7Tp3uXGwUgRcDRISH8
AM4LZ6mG/2nk20Lockyp1hLAs4UgKlwa62W6ViZkdvYwP7tGz/jTtvyRFsyRA7puf4XQA0BfUqG9
lxfICrD+jAuASjst4M5kNaHRot2jAMSedtV13l3qv+NDdIMO+ZOgE1C9sntfXyvSCA7+oMcZ4SbG
Gt2ZDlNvsta/r+vbvfRD/jidHuHiAPqrdLow9sRb081bbKiXLjOCYJM3SvVtBI/DU1Z2xCP2lrvS
x5uWJtcevfEnTsEN4JLfYS73IK9EGMVTdj5ZPIBAPTy1mZY8I5ZKeW+mcQwIauChAUf7Z7wVN5HA
bAOOU3ocppcPTxWhV9sSxUdQJyn01xiI1r7zHvREAXCmDvXiXlTR8mZFCMjngwlE5ZRgxTsUrOEt
PdElk95HqU6qNgNT6uDtKcqfeSOiExWmZlmKilRzVzVnsk4RZ8gkxdfyf/reKhITVQNXSE5RKq/i
smU15b7jlmF4qXlIfXLjG8S1D4bugcDRAn9iRxRDt5Nfr4knJBSRYJh1L7/imxGF4hChVuhPS0aE
FPA++8makUPWRenddxfh5NWiVYi7zUKm3QLnHPif746I0Dkkqz8/JvXAoTrH98ThgTJTS4IuQNCc
mzUHeYQfTMWmphzLupbbMXNZZUsHUP/V7B6PYgFfTr88zHMtkscxcBfn9rgbPd5pDVjzK/hDWtJ2
+quyG8fRRVBas+NVhiJN+hQWzHXJvoBzSgAKIyCzstFgkA1DY3hWRc8J83p2lAgRt3DpNG2i2m8z
rW5nvKmFmR6FD87/Rwk3zIEg5bwQPGznnQwZzWGjaOYwQkxc4BWzRcCzBvEKdp3HxgifZCYNUjCF
lKWyMbTFxk6Qs/aA5uSaXoNt+LqRP2J1FqDJYGwRvX+22ntMni5E88SV+tP0SiyXVqWHEgxdkqiY
vdf2NlZ108u7btfcKTlPNA/cuzAUwpWFCNfGmnkfXiP9fuIGd9Wt5Ye9Vm6C1rz53khdO+fN9VjI
kI4ahHhMELpV7276WmUt1QXqD3y9UuNoMBDMYz5FHuT2O7UKR/p274hmwJYReKW1RTez/KQ1hjDF
Dx+hlIogkyCm8ZOo1GEMz1VDKSv5GrX4twkXkg5ppq2OlPnxmDbXxFdPs+poQZgk/gktHsKVrfj8
1hbFJJPzGM9DDFNRZZ2MBzgANm7MjL+S3ny6EfzN5lwL7Dr3dNKl110aMRxA/y57I1D4XpFWv984
tPh7xaJiCKxUWtoZQRqo+J28I4IjApRD3OkoHQzJSMkj4aj8+w637kV0xYZEYIpJH5s2ilgZqC1n
sTKkZFi+cX74FvPNyyxim6xFNSsDjbDN81/1xOHh84MShyAAydx4qRY41iXCet2uk07TosIpXBIO
Bw++NdDZPOgc32onCMOFjulxLq8loWIXjzBOyzMl6bZZFClfyyLJsmGVcIeBrPFxYIwLwPuEl0Va
Qixc/Hh+wuXh7DLpPd6WErCKthHwqxRsMqy117M5Clif14XUCgxH+lQGBHwXf+b8Ne6rAkYTC+44
NM2vPtahyOdSMVX92ZQzFUwtbmuJ3Vks7LqCwd1PqiAddYTf7G0E4NASCBs95vsd9uo3ajFZQpdX
zbuPOQlu8USpN0l7CszIsnlh5HPtXDMXu/Jvsh02X51LbXHhdaONgzM0cSbQYM1jFIFHvwSs0/0d
oGNTq+AmzzGfjOozPOiimx1+E692nouKpGNzCkEVCiPufKJJfY/XpOShPkCBcw1AzPkW0DC6FM9k
Ums0ds93/Bw/RZOeKI+49XESPdyq5piFsX1G3s/3J/K/B8KeebWEZp3Zxi3eIPneOVnsmWfnASUF
tsZ+p+zIJ2Mpvk/t/ZEw1UrZZ5ah0bRZfqDMNizCCtYlPjDywqwey25QdX2bQfx6BsgoTKvQnK2m
83sqavi/obT3A+nEp9vJl0XpKacbFcoNxgrzl5Aq1d5GMCiwD4oiPNZUBV14pSPskgD8UQBUXNS/
8MLckBTCOI/DFPRN12Sna9wZeVchcAUSaPnuKBXAHKRqbw+bZh3KWy1fbL7QuiMmauFr6j8MfAgp
qveAbCZxgzREabiuXOzsAjrLVUSWwxNBS5yyScft+AJobTuPRbuK4AZtSJCpcvFJ9cv3TBTr0OFm
W5LKOLeFYQrMHOJUxV4zjilBqgl7EsZcg4WLMGic9z0ezFr//gMb+V47o1Pt3cp0lH6YqPNxk8Ho
MJuGNLRPaNUg55pv2GQ74KImx+TmhuDdXGTXNF8E+uf6FL0z69vKSO4IBpCQUZVEnGh2lHYocnm+
fwooC8KJ08QLvaJiSYD5qkr1uXlPpX+u8nnficvyvUYLD+YjQiS8kwh+G3MMYupYIR5AAojPYWEU
YH2vWfGJMtwRn6XkMLFC2mjcKprZjL2K0RSNEqe2ApXe0KNRy/1IFDZIuUe9SZI+suqWhSFXShsZ
bYi0qosVjTjWTLb25IDtK3AldJZ4+fnbqSwTjUkvVHtDe1M5Hr5IJw1isNKu6cLG0fIMKoPRGLFx
pzT87VIZWVeaWsWgB/6kIJFlxm3n23MCitjs+uWek2vcKRP6Xb8VOBD/+yIqub1CF1c6ANbZNJYD
ZwyXoONkhrSJwKd9ebpI3tzHjhAbsvYBcygOeuINyM0LfxNr7RvDzw2I5Qd9evF2BU1ly7C2jRGL
JQ/viGXBouOi8spHhOg0X1Gy0duIo3wPQuvu842+U/t25Fl+nBMyimqboYgQB1BpF0j4VFllc+qO
JYl5yiBemB0mtlZYaGdy7vrNQ1/CmR3QT2w++5oHz86Qzd7G8qXbuK9Rka+oupyK3Rizuo2p2WTn
GRgMXTeQtfn7bBukffB49fe11fvG9IXOw0qu4oypu8KlV9WsnIwqzNNnGY7U/IL17rt9/kp0WgGc
OT9hEa84TpStPMgnzoOOtworrRc3Zg/su/G0ElQJvWULFOuC6x5tNI+4ZfjrEdQirJJcoq+FfamK
kE4IBToduNJYr1iKXtHDxnURCmUsIuiW6Yq5FFfuHSreR0ZlQ3IafYLOx0BYRYGk2pS8uVPzMsWC
fbAYeGrE5jNheWTt/vgn12wdUMxtJntpTbN7CW3g4gXpR7NgXYG6Cdp2K7bMkahxhrhEZ7SIO7We
+8E7NaEyc7Mvf3jtHXm48GPpt+0gr0UQzVt2LqNmGX8ws5Jf9VuEbhbTZl4pvsyoKjtiOYXg06s8
tHs+p/ihuYXMYy7gFUHz5W+AjfGr6HUvFQ4w0vEd4q20sRrG9utJvNFK3l3KhQmypDEld1skdWWz
VqhcxrmwNbsCKVzaYCpC5Io8vNq+5gDspDh49G0yq7Z9HIAo80gkghcEdBxy4+EJtx3j9uK2f6gB
fAh2noFLXUq6nU33MuYWUKMSc7CBjjE1MbYVbiR2RpfNfgr3k93EpYDck3KFfMiZTKncufW9+Ytw
6CdnDLNDCVHy0zbx27GkG5f/Hhud2TRB5/jhXoSR2ncyRpm89S4ShUEAt7FdxIuLIvs08k82Aj7q
MdsYjl8PabhWRC1B2F7MSZNaZ5LPr1ukZ8vNGxs8DO+zwSFsaZWFxAOP+VqByoRB9CasmX9T6/2/
g3XicmDdE8+E6Eh8d89nKG6bkTMQMudH+qpZPik4GhpaQY0r0DEyE2i/48lp00LGijAo1o/e7t+N
0tqrKVdMyJWHd8zwQjczSUzZUP9ff1Z0OEjC0PR7UsBaRq4c66bOjZj4lKmNNwsvQ1Qpw+LKLyG3
58V414KfrbuqAkjOnlWPh40pavN51MTQmNnSmqGeHlCLXP3zfPpSoY2TVNYhdxWI+x8AG5fqHR9G
hN1X2fx66LiMTuDr5tgvSS2UjHXsFrMs9ifqQIJYY9djapmJ5iHpMvDbIPB3bV2rDH+UMRft+A/P
dx7PtZ69oa7BP9Gt4eCLup1zuAe0Uh5o2r6k/a6iEHFw7dcKePLI4QWmifw96TUM1HK9dQD/92Ff
2r6d0K2VyDcWUgXmA2W80IZ5ZnUCmNd9MmWd5seagZMfyNx2dL16HqYXGYXs/8RvAk8uiqNzB9SH
Y3ryHIJ1xuCjSE+01e5SOUC5c2R4p1hkC48q+HZGNn8dg58ot+WFqbMzBuVKZcCwbDpVlRstS7AF
tyItBf4Ol67vIbI8KFjY4iaYrghCIT7x2vsiUJoPEOKHgtJn7lqAn8RF1NFTyEv+VImx0601u132
ZzCe4Ghwl5pCv9yLSuoGpIj5LKjFtHaM7Wf7Vk4LaF965ZIlCi+EqpORl6E+EnIBpIDjoJm0Le8r
3jlwWROdEWLS1ByrJ2MfwXEBaqPM5OkgtnxXOIAS6hlmVo7XXXaa7eU6JfSy7cwpByH/2s/0XBoo
VCV57kmlKKW0lV1yVId8Dt8VVHwiJ6Hv/E32SB7m2tjrurm7OmRhyl5jrphYGhnNQa3mlYsGKBrj
nO5IU/oyDIYXWB5AiuscUF3UOW+qO5fmrh5/2jI1eWKgjFAJGWktPbRCkSTiL4gtRI4r58W87iSb
vk9vxrnxWsunATZchwRpbyciFG6PUstD0g85lGQ6dzngtXZrbKCw4NXuhOpvDKrrlADCTzMILGy7
mPUsVVoIz9K2zelC7ADvVlJzBobzQSL5vpBbfAT3bmAJ4qGjQRyazvK0VPfdlCUp4IdUAos+Okbt
y7IVMvoKIYi9ACUGZzNMRtnCs98rFkWOemAzNNq1BvMFEK916kZlGqH16wkesdDOu1ilCTwTNFcT
Khils255jsdBF0OWdB3yGUOeHBmpds2dkSqGnXZzuQHb1Od/f1wEYTLuBU1Yzhze9lsnWW7qtsOt
RAHFThzfJiJEseW/zSb10M8ZWQPqROiSclGXSCYZ7g2SfCq6xBYxWnim7Qb7Irekg+/Khlzj3qU+
mYOxXlcPJWJA62fhtTtPwLi4cSnIA6BWFi+kk3qFTVf39NrrHK45Cdg0U6e5PtJJghbu1uyinCiw
qt5mx87+5puZ/3CfimzSLftI1oYCgqFGzkjziaYqC5EOIicc06ERgpNG9Qvpx8iQd7WdTIFm7OVW
jwfVCnwzXXzrALjpPmkjoef+oC8ErXQUXKAJtvfdJryIH1F1RvIhmbRx+m+jqV0B2t4qDK2uNS4F
O6KnAns8Uawl5hIX/Vu8fdqjOhdyXUagOCdgpTyWQaZeKR7tv2HIzXW3LaVFkcB/wh0d9kzdhJrp
CMDK+M2z1wkKq0iR7ByJ2K/Y2iv2nUZkFBoa2QWzp6zeqdIOqUU+WqZEvbvPouEHYRW6NMUpDMze
/SnukBJdpsg0qZR+Qpb/4LoAAteAWjYwlDFOlgqcR0vUP19ADNqwLFV3HiKyDDUEdbEEPCPNKgi3
6eDIBaVHK974YFWCYVUyJ5elHtnk9haZXzGe0rUcR8IWY3zFHRLAemzLEAj0HtyqdUcb4VVQDZJQ
l9h07G7S2h6JWKx7eexp1NYfUBZVggM5sdiMLrX2j66uy9/Xv6aUX+gEEcJ14yltzjTXudRuX/PW
Q8TLLYit0XAneMgKTtMlBE1ZI0vTbKWL7FNShi9PYRtRP3Yg84j8OBpjI7g3Y4pUnRO0yS7A93s7
ZvRJtSDi0g0gi9K2+K3CAGempjY+qesIX/V6HXUiQc5afRY+dSSwgYKAPNYB6D+V2KtN7ExVXc9W
41PpnwfA1JsRdQAbN8+1y77WffCdTbChQetU/jb33uCh1YVO6+jAzC3KhhKIZJNCyBgxu/E3A3b6
lMXWmrWpCOtMbfNLJW88j5F03P1Y5nVX7+BsC1KAdNNUU6DJLoA08OpdA5suHMWJOs2XpFEtoMVI
lbk8FwoxmupWJNsLhik8iujUhIiZfC5UNpzIATMpo7IRemb61CCJ6iTJq1Y1/yZgEvqDt8wOwwgD
oSVdZ4eUg1qj0sFkw80SF7VN/ZyC1V/bKhGcnrEuqK7PP+/QPHaGYORuW08GEQ0olEHIMZ3G4AH8
X1o2VxpYBkXJoOzj4JHUw2UAb6oOfSZoMGsl+NOeFGirCy5HVUYZGcqKSXLKPoK/YIbLoRILVffr
Ul1AAmTVbfH5nlBHsb4MwzJpBtC8bPqidgJzN2SYQ0KpVtQzclXDz9Ie+ocmCNM4fsfd4uVEMQ3h
M2IiMKvHCTYLSa+rbRf3LifcVmGbayeEt7knuGxTIADJJtyuaN3bSLjhquuc76zFs5wBs7vgaXGI
/OqsgdDtzvBCoaFDRtmnwK0e+1sTN1O+oFYmlAvZcTFJTRNu+5dwBPf3um2nDHv3ftQ8QSJxz0vq
azlqVtDDb7sTd+AnXGNVTTHmSc4BoFo47jDEewdJL0lJRdX/H3QPlovzVPs8x957Z+28fZLBayEM
RLW/xwpMfW1B8MB7BcF/lD11HJX6UEK98zLrZICaVYt6bhM6aCg4NCWt2t1tyRX1rwHOt21KyM/y
axZm/fr/J+2DMrrbGV4TiL2WdLFTWp3HbpKIfUwN7OuITyZuSMFSwgO5d10/19BDZXEizK50VQi2
F92h9011gLWqhqa8ucX3FyWT/6e9hz7a1A+bCnTspPV6CzPHqvVPLLDamG4KRQltFCyneuaNwh+R
d5hqNlqTsVix//bjF4RW/yAc7zWaxUDfe+p4nWc9LwVuOxZhklFRWkCpr3u/3MpZEYqL1YygnMLt
WXUBf4RQTT9OV1l3rzYPdpBY6Hwoi6/be8LXELdIQb9ESqDKqW+ozDI78DBWBWy3l1O4ijyWMjFs
dK60r2GTtskkwdy8nqXJ5Chv86LOXKoV1UzzB7ad+1i3OqtQ9a+u1tJqHe3BE8wnaxWKYZBVU9yt
8pWccYDUNCKAeIXmeyRm96YHM/fiH7vkwEIbmAWaX5zf6Vj62PhIsYO1th/5pNEF4ZQirmz3vhaJ
w1Hqbg1tlsteXSh+7LGgMkKMOloFRhoM6qFlXVPRwR8o2bb3gDVfm4JeTX7gqmperdZwhzZjEn/2
DYGEPvOJBQTwFzOJCJzVfXAZG4eyhmKRCNRAh3dwvfflhQvh5NZ9Jvwv54UVYR3TaXtJ3rrRBTfe
S/Cv1IQ0SZ8em6/UFIOx0rL11HbDqYuk+UqiGunglQ6mJ5yXIVUyhJM1YWP0YI/pLlEPIgmBj964
1WZkycTkp4ZjXFsxRB9oQE9wMSB0aYUSmrfZpddscMYGXpGd1tYGUqjfia43F6nDgSyOQN4AH2kY
hCLlze7h+iF03jk9uZ5OpWGQZiKcAfEMRYThjeCHN703cz8XlYfZCKpJSzH6zilxjJWYuLsasu8W
3N9zkmiiGWwzG4sp6J/EIv0F8uRARd3bAzn9rkHNtaReQW64uNkzX3rae3UpfsbaPFNF5Hhzbuh9
Rs7P2jLekOnNVBpBuWhoRzaaZ6zxSliuoR+qmhySedlIQpdmxkq2oleS+Y5FTde/I9z/k5BVGeRD
FFwokXJxAJteCEDR7X5w8GB/O+MvP1BKxdrkk8TXEWwcK5h5DmOcr63jWRH3z5KTwZBXH/6/Cdc7
ZJ/AS7NWSiO4sfoaQzoIvqDB22KCR+KB9hlf+g15bQjlseyX9R89VCpC1ZKqsFfp6WOBmYFMQ7db
nm69ugyDV8wLgZW2uA+SISwVrh3OQB+xY4buzYRFrvaWT4ERKZfXIwSGljJMVzgXTZf8WJmY2kih
zOazxR5M7vIzxTEFtyXyZNwwAEGc2npAQiqQ6tWscWO/TqjmXyjaJSrhgGth8ccuAZ/S1MbvXT2l
BM6ltxPMVUyiooop84faA13GCVbBeYnT+PSZYzcuXtn+5NqZh+t2X0Swpn12JQdrgD1rn5X4Fon1
ucQ7UyzW8SkcOgrjygbpsuF1opYuVrnV9ZgHSuB+vfwVgimOO8sFjcXHWVz+LTcMUn/FeAWvVNlc
+EqTmojPZdQmQkt/gRxUBBSXzD8ONcSjmYG4uwXJHfrXeuWiiErXtPW5HrfbrpfKQ/gOECNYH8Cb
5POKLnKiCJt68MmxGepoozKk+Z1EH9bd5VNrFAfPWY2751LFTnpRJ+abVMdqrUB+Xk/rgJ1ZGxYD
kZy4z6e6xe5QOZdvECA1Uc80LD6PELrxQjQN5tQZPR8RXs1o5sPI0ahg0+HsQulae4Sm9MICM2hY
Vqrp9kpXJ198DsQUNpCBos02CUwhf3zElB8XsuNfh3w86bDeh+MzKsuJkuyKmacIV7JI/Ctdsluy
ds+jDT9tnt13ZqB3deS0ePVvco4MDNy5virsKnRUPWwrEu+GswoErKy403rbjCJaNSiIRDsELyYv
jRGFa8M9JGDPoQsG3McG7ZRoTYRtQdPnu8hTr6AdH1ThD5LZdgSTLH0+/cKckPqJMGt/7YzkC+0B
qdmczykpfJ1ioVYOJUYOlWsM9RJIgLyr2dSjXK4t2VOK5CFlSOcb8HDwFUs+o2jrLLUKXeySoZyH
5dYXv6juTyn7rxM0mriVoJuSciyE8c3O5SjTM2d2duH639ElnemvN3+EeY+Di7TTQmoO+NScDHLo
uG2UVWLT77qQKetuzFL8Zw6JenI+ikf3PUGTBFc6jvCelbwiwH5H34Y4xbk8y52m6+ohljn0Pymo
pEf+6oo65Gambrh+eGS6FnYfOO45dyHnXpKsD7NjZBygf3qNhDfTG3rgi2QvWOhYoSeWvn25TCEN
cA853PxmNiJKwMzhEBAwfJKvAmwTbMvrPIFyaN1LVlqcaM18ES2FEkr513U7THwY5EWRhuZ3noPn
aNLsAtTT3Ql747MbSW/+0PFclFBTdJALzsTWJEmoRtukvkblkSIWgdvKBGSepyyH4n5Pjrig4waM
PeKxAEsmkl9y9YBM5vqnFXvf5TF/6UWReP2/HgI5Uk1TZqvhNQPRhQh+ZXzE+8h/467GdNB1Jp2l
gi+Jq+C3hN7v6frE4D7/yXAeqzqU8cU2xRTYqiOszm4A81bmw4as6vSDjzrWnLFi/l2g06TYDNNw
6Ah4y5yfCqq73wJFbGQxLC9QYeBhfkTf14brwlFNyyodUAjOX2fqDzTBhT5AenXZmnRTElKJvg26
93BlaTjgQFf/qCOAhors2Wc6Ifv+U95l9Qm+4ygy7Woze5DYVoAy37r4nbW7dEB9PFLy8zyx6+dc
ple87s6I5nhBWGplsmoxoOrZls/HbnAd1KbxNA5fHquTZhUE2Q3KZwgD3EU/RzCUSnZZNxxic1UJ
nPcGn+Qqryzkg6j7CgUSUET1ktPLo2g74UQLDFtX3tuRo03rkis08UwToto96+9DBQQcCBG5I0QL
IZq8aE/K/+sdDSzi83rFzFtsSfX/br1CI5pebBk4Qs4cGcMcj8vAamWypyV+zTTT+JJaqDOtIP7J
/y4UTM+ahAlNFdOwSWVY/mXznSM/8owdWM+Xd3ELMGinpI7m/bxO2OOY0TqZlBz6R+/2dzbeF/+m
MdU6BgbQ2Ys7tVGaJ+D75PfNJlF2FoFiJr31iqsEh3bv6A4AS6iIq4/QpSATVWwHQTyeWcWQ0QS+
+Q3qdPx9Bx81LAvknIj1AQ2qeZUDfZt7tUPpgRfrWPhiq68OupVg2YrHZ4KlWjmt2n70HOWalDCc
o+uYtRjbwJRtRdtgArPE94AheoKG7PQZTGNVOMhoj4+SgogA/WGjuKJjaE2xXaWPcaz1YCz9+c0o
ekYNVlUVZDmzn1Fmc2IGzFyfVDJKu2I+3NKUGpBuJ0VOhn6iVKaeqkqWTKbLFo+Wdbw8dkUJCzeY
7QsPOfZT/DRuetcNInN+SqqFILHS+XgWxHpmR+x8iAqq7XT18sOISrMfLA2pcInE/ORR1FWZ+GH+
mZUHFdNe4naVDT7Md8Hn1bSpnDZZVb1p/89ca0Zyu0kx0euGPPxWSBJL55QZxXx8zII/GXJ1DR9Q
BjVm9EW0vj3NO27g0H03BSUWV5v+YYmhHJIU4s+lgxKykgJA4ihkWFvt64skDa4uhFH2fqDevrFF
fXr0WizLzU6UxXD5x6lNsU5R0pnhsxPo1BrymIJGgKXCLvY/PcBAy/bcjjRmlWnwOyXwRD9yV2wj
WAoxCRQfX5X/KCfTGW4an3Pj9dr+kkSbseX+yZNRhT78lcQeiMstH31P6JjyA4qb/p0YVw44P0L6
nc1PrPvbnGodeMlF+VbHFhgLyAcPjNMPHTdJ1wqHmtzFYSTRzIBeoHBZKx3ri2kk1fQj48Ptxt4q
fpH97iSPO46Hg+xTU4IrG66IUbVVKjomGMAd6m5XbnkiqrdFQdM299uf3cg7WCVlv1oPtYTMXasH
zakcBcj/KLekeDJ/ubmSmmdCwoXFFJ1Er+3uOIVKu0IAzn3ef1Bj5EuEs10L/Yjr0sHSnRsrDBgr
7eVx5MXoO9rSSh7LTgssZirWrY3COjrHiFcWbbjTTk9/Ghtm3HgWBTvlfKeJoe2W3YYwU7X3wtPv
o3hgKlS5ObsGzfQB7afZJgx7ipsQmNcI63j5BeLpVNBcKk04YpJ59B7sWcDaGOtKpshTMns4qDKY
Z9GTm/Ox7625SguQc/7le4O7ASyL5DAh7FcGx4tFntIb5XKQ33yNXZPVwo/fj0aQK5CDRg4vWZOH
hqjhLQWDuC9aAeR4BfVniPazonV7/b3zBgyIS3YDaUgbFybofPEs+KasmI2DtiTZLFXFft6CQQl6
yQ6x+fNSJv3gl7t9ziHNnVL6JHIrN74ZZERxzYcY6d06C+m1ysyVk76zFopMelBcAHl+u7t9/zn+
tc/t/I6+Y83G1XkAi1dMmxqYWWiykXaYGajxl53Fa+MaGRHijybi9derlN6AF3wipCCIxa1WmGpq
BOp1ulZH9gZQ2ICqhlkhT8PYN593uOhKwvFEYbx4IT+kC+v74ZpejZJHERs1Tpel4vYdblpQq2/3
1Ir7Ydnr/cnQ3fJkibmQwONca1t7dYgpyc9APbPlWs59Yzpnx29MMVtYrL5gK9RniYD/qNd253Bm
8mve+vJ3PmK/4VfhShKME+5T/7rXCKzrlMy7KaImO3H1uB6WnZuiNOuoJnqWd+DS2ynDSG+QUnRN
s/JN1K6rrwrsg53mnKBjZZ2EJ3MMVD82PQSbwpCUm1jP7/X4pfQK4rI63zRlgSC87l9n6saMqz/2
HbkxMA9MjRoMNrDEzJE78Vin+zb06G0zvloRVlzI6uwLK44KUvF8Dd3o6PHhd6bBVzCuSRSWjQ3L
gEumBJ6IY6Bt7hD+MDZ5EQYz/TZtWajHZw+RMIvy3u3I3BJ2LhnqEpLUaKbGyjikBj6wrx61l2UP
i4T0uUntVqSdgYgA19fo7bNTyUeZYi/yN+21c+zAISwoSeUjqP/5QORDzLgSODP3iZZxwE7ASjgO
+DbAG6W1zxW4DD4o2oaVk8CUwTPsge/ccrMmzozrAK34zpTGxrC7CKYoZ7QG5Z7f84V0dvbaQgs1
MBJXPZOs/DnH72H3IeICcWec2R+UcktgUAg21848wV6ftrg8LYSnha3lOAu66vtQc93RMiQgOasS
RGA3dBNqIjPs3ple+eIq38u+jaXWum7jPKACYtp6MHFFKvCTf2PrYLwgxcZ0N7NHRMkMeCB92XsE
t3keD9WJnsTspV8PIxGlltj54GK22Vex+9qBG6+LtRAyXVW7rL1xM0Nw7zE1sX4VhfChhQugLUgH
1PRWQOee74bF3IQjLFhyCXifWu4iJ+tFqPaWNvLOJC3/Ojvr1wqOPQo3ZA4aaIkp50K8tzI1bwSF
SgqDoZWDaGQ4W0NdwcVUL89NdAygfx3NZ815KB5ghqSEw7brLRj+Xlazqa68910vJ9UvmnlVYoyA
zkBtW6CRropLRkntJblqmbpmcSq5iObs5LuX9XowseDrRrBtWO2idekLRM007QKVAAETS4ohIYJP
zb6nBrBoVbb7AINqdrL2IrlvGyzkUC/Xi0PjxQ50D/xRgGgDubGBz0vwyU3gnDRpRmUnAzfz3VJY
9dmJZdOIHk0di/tAuX+JZsl4HFCpKmOsWluU4E8T3yGs/CNV8UdMEVhBwzRyjsM0HF2dSbVrljtl
xfH+pGJ/PAe5kYJ+tPG/dMIwmE5VTZ9KYgvYLNoFa9vLb3pkTBvad4sbLYFQK0SUJADMp7FXcMER
+X8iXAh5hrrlr1OSxz980P2za41tr6u6Il5F6dmUz6Ey7fERLE3aqBBFs6t9nQVKYuAyqnqsgGL4
uPxE36QXjqIXcwuQCcy3iNhtm+v1NoTtJ2Vn0GbMIZT5j8rI6y2kEUoU/s11u5M7zmYcJx5p2o4S
VT5ZkMQE/IUPUoJZAijat/LrB0vzlOqj+btbdpRJpnsd4ktCQDjGqONGQX+lDSxSpCp8HUE3uN3s
dlA7zIfzyKBVg7bZiXPLqcAo/o+DiVFfw/Paxgh1KZjk1CwK1oZWzPvUTOK5JJR3IPE2TPZ83ver
ckN9KVgZK1p4CzvSgxxO2PudLEdx/AqVqiJuvJXrZpRBdZD+HVAHe941cPHW0/RNU3KUGHXDPBUE
KlccA/IJ2Pbqadr4jwKMB5RY3pXt9fSCOf3qTSU1/2Q/3TLFK9vDESjIMrI3YFa6mfWLCkBLrAtf
TU+kyns6KuKwoo/LXgfyFAOHFZuS+XxDAkJH1/05FsEs8Qk76MqAWufYakts3g9Jq5k9N/8VoRDa
p9X6ixQP0AN2qxmAGxudgpFTtae+7iO6vv3oaiy/9IwFQA4JA1la1jj6A9S3zOt6gwkxDwYlZrOZ
jSjHEieb30GgLE7F7sXHbNlad7Usbm+Nf4GamA/4Ais/2Q+Ng6AsJMDY8reWalY0QwZt3XJLf3tw
W6JMH8OqZVyDQ/pp5bvLtf7CsmqdH6Tgm/7aR7VTr+ujF7om/KlFknRZXSYVfjeeKqz9GEevymH3
Pfw9DaCfiB/98ggi2PlhffG+0J9IdJeC+kT+vbHt3+mmQvD6HnE55gag42sg72ZF9Fet1lF/VaPZ
KluMb7Si/ADmawqlL4QeS4dVy41r6FNtnzsX3i6Y2zgejBxKTDlxay3wt91sV0sk96HSGRHAiuzs
VCc/a/0oKch/ukFqvRtl8x9UlB1DIRNek5nBPnZt6bRWnnbboekhZkaQc0MDp7GpJI0wWZkigfe+
6lNA/0xUfwGLtlOvsUZPcSDP9zzfxO4kSVCQoQUz09VJVeWfAB/+8PPk0r8kx/o5DcTzGVx1trW7
qfx9bRdfdK0BclPCMv/mKDoJTOIueNAR/rHoZfsjS7rvJtcFLBJ8gbmTd27llQOhPL9DouNUx9hr
EXUVR/lB5VqUFisOpjs20t3ClVAkcYvZa44Y5PX3pQ2ccNxY3XBF2tZnNWVz55MczRHbnUQpiIys
ROwV3ox15L8cP7l0hBmXRXdvKbxHNZf1B1ErdoPp/EkyFmpo8xI8Ibzrcb3NvoTCChckHiZMsk6l
i7d52QTB5zd5lMOnHkqiywY9AYYX8f0vMsj7Lcdii9KD5MMWvQMtjuhRG8e4RtFtEItX/bUdvuhb
OE1B/KMGI0sle6o9wG+wHHQTazWBKfh1jSgY1Q8v/Dvr1yWPZJP3YgJ5g9iw15WjqloARliKjaYU
BpMl7sc5EvQgwV2WrdFxY8Ww8t+/7F2JPDgFS9WIzpN1gjGFn/fcHK8d/pDKZAa2QOEMaTlVV2Vc
rz5i22T37FIhUPfgi7aDSLtZPTmsJja+bW33mxlecAQxCo/SELhnyW8q1clzBGFFdfGbV+lT3ZHE
sJbaxt/LK40YkgNtaZqydIVOmvFlGPd8iu/W919D9PEJgfJeruPCwMF3Q2gp/zgav+VK5LMsTg3L
hG+QL+CcvNuk4G+K6B6Ni93sfkaydbeyk3/ukdOyPvvs55GZirJdbJlpxH2DsXup7Ti0Lsh1t8uz
BrR7ysP0MJaM7j+yrgceP4xdc7Iqzts04jb3m3ykumKe3jKlRH8lYQwyrHyotJoSTybVV2Pt56JN
9tZR7uMsbrZPyJ1wI/AJ0K7/4ryxVbeF3GmvHocPvmGV1GYU4DkFx2MYLRfnQh/6ZYXC5+a/llpm
2JQzzHAmkGUHPxoVoMOT9QNG9T7cIIU2ggElmxdIc2ELQATuZ1kBHeuHZZsBqc6OAgOegaRqzFRq
ADUOYFGSJI4ens9rJh7osdzAyeKKSh6rpuNcs1bOGaxuwYK7PqRiIQhZEs8nCBIEuAAoT2p1VOlq
nTxTmrzOOGYfR3lFZnR0QTUwmYN2evSH5N3P7fghjJ04LLXS5rMlgK0xXK8AuLz1jBekIGTCCyBm
ZZEUadTFK9nYf6NUyJYKsOdJmQO+P4/AaDVJmF9ui25BlsCOtwZ/YDCvDSMB14RMJTOEXfpKuWkk
T/Nwg39WGURG7ZB2w2sh7UcwbUdPhu1D/tM+85aagap+u2F+8OMIwJLLFaocJpa8ebdmK9BPcSvn
YvV2ckfK5tDZTLq0YUOh4lhxjV2h+Atl1gF6oJa7uSKAncRe84Ub7Xq3GvKvVxz3YZu/NGYIOhQE
7L7ZeA5N9w6fQsYfn45X7XqAomy4gtvBJkyy9jQiSamH7wyvXUXWJD9Z3SU4jInThjwUPO6lE/df
uTBznWCpyVKJbGyQ75seM2cSnMJ6U2UDg8JXr/k6D5HEFMkEPDSmda8xqOBPoTq8nhyJzF+DBga3
KVr5FY8RY3sFvzQB16Ul9laxN1yDf3Zz9d5rUd/mp9A116Y3vW5u1Gu7nVWNU6ggRLZOO7jOfs35
bt2Fle6ZosUbd2hepF6AC2q8gXwOJFDkHef9omNllme1N9rpx0RfIdrlqx3S31x6AUt8ciTo6FWJ
me5Uk+eO3J2LoS0AuO+nGzpPC2PCUr5Rl/eKgZ/SLUzwtrLVEkAjs5uZXVau4T/mFLgzZ7Vktp53
+SkojsJN5WguJTfvoxnGYHKpXsGUcgkmdVhdOvcMT9LiP33iGf0Wit1BMieghabkAIxB1Pdqrm5W
gM7oCTgPjH2DPtdftSR1jKX49PWxgyEVFoDSGz0N8L3pL5/5dSV58mYI3He+Ce6a+KtUKYccdRei
85Cu84myin9sFB+m6T3/K0cx5T2a+N9Zd4zlqCWjbswC9g4yeTtD1+KiCs6X/S/ttp6Pk6KnB3gY
mnDWpf0xwkgRKoRnvyzjEOc8vNDPohzHgdRSdiKZep+igsvW2DGfaVYRPkKA7vFKdNJ0KooXT9xg
+NY5H4WteWGQCFFSHwN3+wPKGuPvpBYLSTRBelLWq/5TmZUYzW2Tq4Bi1Zf0DJNfJJuNqXhjcQ+x
zc+NFwZOiwU9DLPOo37wT7ASc6/mHGaNgsJiuKSuJlmo9Bu2zvWUO4HPvYLPZEet3r6pQbk1Vm1C
a21Srdcyuau5dtVzcAMi+BjZdmO/IaUZbGwLfQEdfmPtqD3yzj4Rrdc4CSfsVqpfQQ3BxsEzYl5v
xGdZ8PKTt+PHfVsn4bjsjF5PgkTwT6HVPG55yF1WoNaX8Q18gYONLYdvPWYUZJ9zebl7IXL4duwK
t5V3hQUaKDXj/nXBaosHfGePtbX3ePuRRRqlcv/Y54Mo7oGiYf07PWs4DTfYa2bsuDdQ3V7IdQiB
z9s7H2Nh8WcTIjpQthHbHs5+NMeosJshxxzJY8n+i95SihNssI92FD37Q0rOUQEoTu5WNGmZcnaP
UerkhANNx5cf8Sen4GmRw5s8Q4QxExrBN89KkEy8oXxDG0u/GOOgzU7eNbxZaUXCIr258DQGnCzN
bSDnNvs2DGxLFsxWdcBankB20txXKRKmVAoJPKg2q5leTFv+J2xE3sM1b0LzrVETfVk9Ke4TK6Am
f/sE+RVAygUf0W7yEH6sl6cDsCaOyBz37EmlxSjrhdU9oOUmsnQLpn5+a2mSmTmG/tPW7TcyvLKZ
earIdkO2GqbGTd4jRfg3bzB6YW+1E4kH50ICkEUWQNnPv+IjeDuceYUSe92U/x5631Cpg38i/6//
wnfWMnczxuL60xWTsANOFqEc3sBFOcZGsnaBgez23AjEiETj9n8At3LNCQcEJKVsya9lZVDDWnQA
DoeTH+YCHXVLtnTmJxFqAkFX/R0s5qs+7s2Va67n65wCzqTSsjvMGIMK4dRyKY3hQJK99Y0ZEqti
sqZuN9iziWYPf7zBALMcHbBZjhgodYJT8+GwZB0qxA24WYp7PGcB6BNBKgO1P94mpgBZUes//zdy
KUfb647DtSqluvEXiRO+QKPMiNFa4t+5HjPYU0hJFXDA4FglJX075Prd6yUeWnlHN/WTuR+BDhtM
zDqeL0IsTlbAOc3aDyTlYCxZXlBcMXx/gWpgVrz1Hj+eUokOSSntGKBigFPsPS8NeDnjY1WbmZrh
fFm43uz+8Z/tIxxb8cdpA+IBeoXDlJf1mnpp2hMx3pATPavPNQ1KmsUTYblnGZE96d0/nOjU99Ys
jlwcVAw9vy5TBBXalTCDYiJVDshsoT17h8GLe9USfS4d973aVPLbh3WGveVQLR23GSRPLvzPfRWs
6lpsYx0FlN6BHqgTmoKa8+1jpi5x0OpWo+0KTKTptDESAMDnAOTpvMtljMebQLsqWJUMJ+LIgIS9
I7VFRPxvGR56zvABdfSi/HacVGfT0I9xKlIIDNnmMcPGT9CZxgGE1X7uJwoH4jlEH3q2njzrjeLj
q2mIDUw1eV+/OX+6KcgySmbsOX5peHSB98pwkowEXJ7ioKuXI4A6UFWV7YT4N/yi/FZED0qPBaau
x9Oo4K47o0lXMO0mRkyoLivV3qQAowkJr0cIjK+e8j6viHl34UQkr5VtSh/qmVANSmXFPacdR1lT
FFErDFsgYAPAoCt4t6terYQkq+V4U0sTurpPwp1Ojr0hMUsYat8+KZqklHiHS26/6eswz7hros5e
QImSDSh8EjctvUFEvF2GvD1AC4dAOkJ0uY+ZZHqGHnmOmsQy2LP9WQvJLu2zW7C4exPmj6CBfr9I
CTaKsBX+U2jD9/CzTcEMB0Anq5OlQZZXGFYbwTi9znG8tgJXH+vdVY8Yauv+wZkzOwzYLRbEHWwz
/iCi8S1UdACBD9p2fZCKOKPciJmIqM9aK24u4FyoBVgfQKPXB/iN7fPpxjJXu9/Vcts2vYfXlvf+
+OXtObk4+NhSPlBPb8R4WK2iDj4VywegemldlBiQEaPLuXkfo306AiFd0MgNkfeCV5zR0WSH2mvP
x5VZB1jeAgzhTlVuwRawxUCps0cpVzH13e7WxdRvbtI3Hzki13qyQnNKh1DusQFpAN9uCMvdYCRC
CSkr0ZlPLloZb5wVHFMAbwzEanujr4UElEfoKQoVDlIgwseONb7bGm3zeIgSSub4G4srbJJYyrj2
Pb1qyJufBDF8HGSSzFPEIhY6ed0CiLYn/eBwOaJjESKb9rWsP+ojjxcTHrx993jKV/Z7cJxB2kZQ
6fZLBx/gOJAxIQlrbWfkkjbAk92ov8rqDxPzoALK/iWcT6GdkPCjPWCPhvG22Ftl1ox8zg1Jh+pt
Cy8FYwhvZ1O15DZJcksFFMKyI7r97dihHs5Cm8yd3/Hxyf05IFSr+pSYkQhl8C4dsBMywz5M1TCt
yRBJY4ap38Do7T9WMUpai2tCeM26Kq7BaVlFK5v+0R+mZ5eefS7Sf91hjRh7FUk2gG6K2hWA6XWD
WueS1dYjzfYHFOpUUS81SNmTt0xFdQ+2wfBp/+V2LXjt6WWenaXxm/5S6bmpcrM2rSpt6p9AmI17
NcshaLgBfqq0p8YKLLX3x4YDt1SjjFPpdaCmtntqXUdFLNwD0yXdbfmryb69YRF5nX5p2mhHV8Or
EtWdhgrt4iY1hV0BXnI4goaIxOH2YMCMOP/sEN6x1hhM3PajowNXT8ZbRhB6qiQp5Uj3UIW/SVVj
YMhtP4agzFMepGyerjjvVV65HcQ5XKyen+rNFKHda9BYbs3btM2kMpS9a6WsBCgPmedSGEbEnSZH
q8pQemPfydjMQrLvF1p+JMn1JoqcQNK8q5V8tmXSaxiDkNAcBN43yLKglgD1n/pxg/zP5D2FJVFx
zbDUs9ZQTQVnBpts3xwpVlAnaWHtyiBQN8fPXOHMtu6wUoKlvcR7TFhqDyCnDDF8gXGuXAK6+KbX
sC1UoSZPCW/c/OGjbUVPgYfpHnSonEHyLCMl2nQrHeYa1WmHrv2A3I+oOClQ8j7Nb8QEkOPDVdjt
FteUMU9F5zHnNkjZSOGsGQaYfmADW7dSm4OTLEPed820rFBTM3u9Rys3IEUAXOlndN9Uo3md50Rx
0EfpscAi5JNTi4Gj6lE4lT+rASHeljOOvEMVlaAUYtvofWMcz4qIXzhjqprJqqactBnvK6CXk105
cNalYcVttaxrDXpInvVweYyRFL3QM7/cxgSwdLHC0u1CeZDDuK2xIEez8Cxb95Cam1mbbZ0zuepR
djV4kzdZ/T0cvpZpoCu0pTgJy5SD8Pco4cym95EBj55iEzzmyYipSyuZe79MNLtqXXGXYfUu+Oln
5j/spgE2hyO9LbPk+RGJD3QAXMSo1OdQchZTgiPN0hCvPchoLCMJ6V/x97NpqsCESvCmOA7sm4PZ
83PKfmz5jrZmLpR62kZEaC3iU0pVWz+oLjvgASZegC7NQIkryGKS3jfcEG9auzv4aYFgHcZfl5C3
BWXQtlVIG0Ohk4qgxcDJUoB3Ek6sP9k+/iw4bJcz9dcO4r5doUc6HPnEuPJJ/brwex5pvYD3h4Ts
yhtJ6Sjh0yHSUzKmQYdsxl1Nw7VczL0iKZNw7FUi2Gl5lsXFbiClxpGGOVq6E4K3XlVJx8m1sKaM
x1QtfL9+oPnKEVxjPk+GmiobTTnkekdYdxSUNsJ79cG1q4Si7MOnC1KEf5a4tkMHsESKdg10fS8w
G1EoVpbUC42Mx4ycRN5Rx9LLNs6H3dHUmvIo2+PTNJIO9CHQwJdVxY4xQ2JcyH6xs2SiBKApUPe+
AdqFuCZjTfSaVchdr2yVGgKcPY5vs/Hs6ufohdTRrZgs2esQ+cW5FAIfY+roT+qNFBVWe/g8TtRe
PGwT/noURNh06G5DTQv6dbyJGJBc1MPQlA/pAgHEZt+j5zTyasjodNgCMzI8HYkFeGPquXCbruts
NsY+XK2JPgjaPKdEr4RctFXG6NFDFlmwgwSdYSK80rRRPfnfrqEa3tSyHesAFNoNDsstdRcmgVBb
BTVj8IbjHNTHSN3LHQdQF9+5tAERq173y+wVAsl7SnKCapf/FiFGyqmSKa+f8xwprHTqIZw+gbof
X1/Gs+x/1BaxzW+EB588cdj5nucMtU1reD8gYL3qrvknY4P99ovPbka6CdtOOWSC0VjgWYd5EdlW
tG/quM9AN3igChiwtCB02CR05B6Nho+a8lRNasvloSkICz7hcRWN9fOOXQ73x4Uovs0ZUqHtdwFK
JF1aEPjryN4QN1R+M/HHA2UkTdMBbm38lOW1jn2pfRDiy+Cq5qAqltGUI76B77LXZMN+sjrwdrpJ
bYpp15MhcBwyjP2Hxedt62HHJeu7CGzbqd/C7dUj7YUGk3TgQpy6S+Fp7LLArdapQxV58oA0wDHm
bnWKOJvdCXb3jXfhd19H5EmG21jd4vUi6k0Q+tqWIX+nc2Wmki4+gUQfbAG/0hHW4rSaau/N75gO
KA0GYyxblKbiRmhIp8BI5EmURnuSninIF25uAiPz4SO4Ql1ZScYp/7Yk/b9fU+W5FqRiHPNezZsx
ZNhiReQkJutWMkzHJ5wzsaFO85pS8Tktme3gatQqYlxuMaRUesbJQsIMLg+rGXWpI+neSXQfEWRl
bRXKWAKKl1P+GAzZ8qvJtR32PgXEMI2aUCSL1Q12KuB42Fi2gnzaJUEEXDU6cvlTwT3PaPum4JRJ
D+514TRM4qoNjexMVblE03dvA5aSinzkzPJGp6Ic+STnfQ5N/9N0NXvEd6AxgrPFWsH+4ww+0/kh
e/MUwr5nZMp9LN8Zzde+Tx9zvexmPIzc3vTucYj5BHAtqxveToEyKDAiV60SBXuMZ64IYpWEVAof
9dkJnIU0fJfuAA2zYo5OAtVOnfFTAHWg8vqgM65iCx3dK0SAdO25gO2vYYMoxFtECSB95T+4BuHl
uurSkLZcKFOv2PVbVKzp4RMUOwUuK/LglGVUIIbWLwR6K91Y+NpseQFb97zVbDupbPxyE+Gc8Lk5
BbV07zVfvk/8IFKwrSBrHti7HUvD6LLZPPs6+miFPRq7bD9B9gZRQk12d6PuqFiGDan3uwyLxa59
Nuv1K+eKzjktIfwIKrUyJUYz2bZrFZuKuLdQtvNGQYqrucVzcxNcal/lrpYDdVtC9tYFocNITWXz
qoy4y3XfhbV5jM/5YyzPW1eNMNWr0dVYQ53Ir6J0ioIxkIgK1j2YHoOENs+N006v9iHToSNa+luW
kRmkHN+svWqNRDzTbRmsbMOh/mIzYHfkka7nVLa9D6g2oJ0iZZTFKQelWDJoZYRUY9o/EFjYKe1G
zR2/5OLCPp6bH29i3dmf6lKroR6e2YGdOPXkR5z/ZAZVMitSl/T8EqzORqeqdVpN2EXNxD2bnlap
0BQitoq24N2Qe4Qa76LZn5e4E0E7bu6hVjMrDHdsEmUQfnxcv5bWHkSQjVYcd8cPE8eVCM3e6tTN
DoJjzJgWBEGpca7p3RZMdIqDpmpx99Ch5ztoAAbMni0NVBi07t9l0Lbjnj90zULWRIN01IcyKHgZ
HUpkgU12vPhrKUTqYQcgzh/BOvCF+mTgDwxgXGNOhsCYw3GVhtjL0bXchXq3IJWd6vNIu4Q5KQWi
ubfTSjQNWpw5tIp9nRnVeXke9cenbQDPfYXJadE0K2MBcrhi0rGdTEJx0UPF2lYx4DGJzYtkLpLR
M36X4VWNRs5GrDiZe/b0jqXVxh80JDAPj6vCqhmlt4Ta/mOp79SkI/L4XR/VJuCMaMz/N8HfMY/C
Ds6RfHHnBg9N85K9TXua9XLNHD/0IVa86/pyiULf1BB/ec8si4NJ+RkG1aa5uAAKx3knSvwx5tE5
EyLSw0pY4EAdymFGa693iXUaDa5lb765hsSIk81ltWnC6WvMdoE4ckcIXB7XAFhrNoNXvNpg8H4E
vJ291biy6jGf0CH8rDmR3sWv59vUlb7mxzYqOcD+ubM6uhL84Le55o8ZV3E9zFbNxZHnln9nNTPt
AnicxTn9F4eQA9FRvSmFYzvvWo6rFXAcFxgbnNeObHgj93cidDP1K0ggkIk0clpcHARAW/Qk2NmP
ageX6J35IcaF+95h9X3Ub9vJHhPL35wZ8eYJvtVPIjq4BGqRC32Tc0dqA9jzmIALpkZaml9+UDhj
OsOihqGejHwkQzus/xZwVaISk3DJFRVvQz8eFHO9sHKwQKQAVnS4m4MgEYSdrJVzLfncn8xBN+Wo
hHHiunA50AbO06J33eLRE7nDNR7Al8Cn9zaFF3RgiPBE5r1+T+mml9HxM10AlLlB79eL7tDn0m6c
VcSgf7fCn0LQY8K04nLbsJ1qbbghSh3y+JKizq1zuEuK/3XewlfRZNR8EnupUeGVquQPf2MX2A4s
TkLAb2UoLj9B2TDCwhHHcZCOfmuEWdXK8PWtQAH5pylP+nzIou6fRVArHyNvNMxU6iAOz1DL43zx
wz2Xe2GuOVyG7+LQJVEW8b2G8pCiSpQsjACHtv0unaWIF5A19Nv2RTNryKpyX0rPLeBM4pYGmQlU
phN6MN7ixaFhOoqt2S41+COmLHVnFFIMz1WtnceHh9vZQCCv5ZLBx7cLn/8rz+l5C35rye3etHYY
Yo/WJ/ogx1oaLRglRbD06F/n1BnsTGCi2P74OMgukUO5qheEi5YwRWW/oowjiUYpv2kGLb60SmlF
2miBHYYUeXI8yGIg/1Pv9YBnSsCraM0+SKP5vZVdqI7E3jeVdHU83P5uFDoGRjIoOrkMptJVHwsm
yv6eLirBDnoPDDv7HQJkQgrXzK4BEHzFcTWriMFLB2c7Lv4rOYE6dBeyOE71mSZ6WZh1C6I81tJG
NL4xgvkSVi3zLUUxbjaLVktStE03lyK6bzzXoh8ytG/BBF5kjj4K0TqprFLM+c50sjbYKATDbEon
r4Xjc2zLy2urBZl6g4XASLnG8QE6y9FA8XrA8WitHo6B9r9ClVXwTocnf1SpptPri68ZOsIC7pRe
wywDmce3klD4nxTwi17l/yP74SnaPVMCQHi1RDV1TAWM68xKDQ2kfGSvcmdy6boLHEghi+BG17I8
jvVTGJsBuUXpP0NmYGghOI/cnlxB41tga/MrM1496MeTKCot/4qDcEMuX0hNSYaGlE0b2J2Ou+0E
bPj0/771VaHRsQaLchRJ1ST8n9+QjcRBzo9Orrjf0hKelWiTP1Q4Uww6XU7Guro8Gm8GXu36RBWc
VBnlUmBDGb9BdRs7TrD7ZzglWI3PQoPPm6hup7PnxvwMTzIvUJplQV9xeFvByBDfgJ7xN3y8VMtb
yg1Wjok8kSJYshHbWwtpYwsw3o8iHMsWENTASOnvCgBM1ABK3W8HfIfDHHRwCUoSiOiJEg/VsEl1
1WXwDI0b0sq+JZnvSUrgG9xYR8MLxciM0dcVV2ut41KYtUrhM33Yf5KqZOYpk/rkwkfvHM9z7EG0
1+K7nLqvnRK9VCIkbCBU+AgokhmhGc7h1pH1imvV7iEX3GQbLOqsnwfdVy+jSDiSHYDnQspVoE4s
+b3xnjEdRqIUvz5AY/FDGldJGmq0YDOTubgEVsxYuw44iDByQIMHgKWePAv3nKfhnFhlDFH9DFbV
tY52ZlmiewELEd79GLjvF99ytqbcjhlm68nyD9eaDmiJ1VWUkvVmCDQMpipYAaUDBT8jBRDdwTl5
LE226fgQhuvyn1UJJG73IyS+CcInYopMEGpUBLAIcdWEinwqnQp3WbkaF3r7qCrGyY9YQew6l6tz
fYpcoQUbtKUjrfVPnqCRPsrUhVG4OHFms8jA73IznRdVH5ipJ0TVQViZodYB3ryCIxEmR+EwpAoH
LXcPFOzozbf1IQEmvzzYHFVnFqR2wDaMjaa5kN/9GwHeBBLF5BmI+O+A0TIJTl/HqZajXxjY2xIQ
K41EAjErFYSShFfFzTFYrjaQcjxOaWqPvIKRSAqtN9KI3YBvqI1h2AT/o4GlanYxaNgMgApYPvOD
6QDH/O+7JjwIdbFGmARdRCBQS+EXxcWD8eGI8Uy8MhqMP+JFYZM6w7aaovyLh/QnrxNCeChx2o6L
N93136erqGuWafnYzZ2WfZ4DPxy6hhLImgG+8NjLsGX3VI2GcdF4AdwjT8bpWZ0rtzVF1lZ9A+81
nuLWPRB8L9YjwRma0ISuV7SumrelDrN+C6Oa77KBLYPZtXC7o8MF4ihIaXUthUoO0zSdd+qSoUYD
Yr5eUlJ2bgS2STZmwyP6B+kU28wcvwtNKLAEyM8+biaIVu4E9A79/zoMeD++c+UHneiOh9Vmy9g7
KgmJ+YP5op1/zLSCDzZeYW/MfktKfoQKU5nxhP+g4xvxog65RSaf8yWsRpcLiXXHhEcF9fWFyqiW
RBPKNNuek4RpXNcjfZfbNECJDrqqMLgkqaBvbn386elSRsAlqA03Inczwc4g/rlJHO38R4HhfEB7
gXxdqSdDUYLVdJYv6cLacdMc6f27DgMx7yjiADrV1VVBrOAjQcRSeDV3kVCyC7Cy7L/4qrxCoVC6
GAXF2aCvgMOxM3HpOvdxRlXbJKSjslExH12L0uSg+lydq4z2DtNoMZ6VEYkhPVm1v88C8xy4j9Ew
dBQYkCgEoVmGqg6Bkd3MwW3ZoY8oP8P5xKAOZEG4iBBfd47W5SEV8rzBnNrKnAVvxwynCNWezxEQ
A9zD2QrkWcSa18WQFc/GpXOjv+59GcjPySiqXlVP6Qe4scr2XIxVYtKU4vUrQE8StwJThP6YXXFY
9ME4wZaORUVQk/4dp502DietFdg495tvOeFXIHTmvUV+YDE/ziFra/lcsTUdRX4VtMKC0mGP7zM+
SFfecOxD6hrgruqzqM3ZuDI1tz7ZSO2spH8P2tTgESINEOHdDMu7I0//v771FRaw+ViNjc6RSvMS
m2gvPyBlAftPkHei6WbUXxJhEMdNYJ84y7FJaysEBWa8cN1YQKNwxc30HONNyjm0Gz2OrM8My/gE
glsPVryirr5uDY5YUp4owju7I1lZEJcFdEo6WgayPWq8qLtyxsXd/rcFvWGVPfyNsf2pqrRcz00w
jg2bcpfSXsReNM7qhcYo63OLYOfe/m4Y78wkc6f1mUV7FlHnxK5sGMBHR6krWocTTIv+v1jflE1l
DLpLFe0+J5To0pxfrlQy0rwt23FGlEdVJvk82dQWqmmGMHN3Olgar4IsXMSIK5vIZf/9tRlT9Oe6
Ms1RIkp9TT2GrALgCZcFnh7ua68x2LMaFiihAsgOh/8Bcw4Wsi5p//ZE1gIsWOKQg+oVr2QbOZ7F
yrK05OU1Na3H87q7JXTJbugnYA6dVL0U3Fdw7rOoLjwUtbb8EVIKU2bvocaVrfTMhGR/OykSn0yY
/sB29HRT2+TgZXuEtrPyehivfjnGqyzpus2z7sjOnu4zL8XF8n+Uj8KiMqHC1vZh2WbgEEXMa4uj
BSgM4fp4YGxGKYMgtIaOjsHehWNAksjTpDcbUzt1l2N9HuxJ8zQAn0BbH/vww2A/+LUlBMVaEM3l
m3qGle01yjeI9ZrdIMjQraEVHQBO/m1bqbnQjQvmy1HboBDmQGu+AEG+JGhQnpBm82vFOkw0gnhX
ZG37ZvGLRwuYgdLzX25yd5vNvK+GpqwSOYDJB45eR8za4JGkerg0Vxh571frNhbgtvPLJF7C6Tai
me7aEl4aJHmEavjcHbmqyyJC6PqcKlhwWnvJg287isQYH98LsG5MSwutvCy4CmUm6uUUM+hOk+jK
gLhkeISbYjnU93AHtPBi/pXBrfrODiZPJInBbtn5//XN34ZeOCmGmI//H+8AfS5KqD7qpSiJ4Ktp
xs/ft6ruGGGLpCsSsIp1/KUzkKDdtXi2t9Ls82zViFn0ABQG0IjIRbyKsTZablaLTwHApWLBNbGF
Gn8whym5N47etLoDKhnzr+oGd2vDB8texC4NaYuA+bMEPTZKnssBbfiiL6h+zmzG6v5qXJJFqDj1
6uFffJoLbxl0HKE3GAEjW8zCwFsHyLV8W6i6z2KEoxYDcNVJ9eMQfGeFfnEGrlQ+57IN/qBj1SPH
25hejCQP063X0K7n2werlQl5tTDrwCy19uW8v1y+Zpif/t42Zyzc4vxIg5a7pO5na55hi9sMsKe+
/ZQRgN9V8pSCwd37qAnWd9w8V/M3uCaUqGJCoNTrJ4aylt5/uYDIyU7gDqZOG1DXkWHH0N9gNjIx
T6elo2JSpFNJ6e/MaODAISwxjT5yir1V0KU2qbEdt0s7BuXDNUMkBfNv+H6u/dIslKX0kdBcBrek
muvDnliLAk3VNk2M188/vLiAcNLS6x27LZqx+ULwacgFx5EJ8FewtdK5GaeUHZx2tzDc4TfyXqCl
CFc82qKgQz3QjKVcN4aEnUa/f5N6bQu8rZeHhqdyhSidxKaU+/t1hpA1EaZcYeyTcDf7d1IdSlM2
RHdogfPBbjakk6FaLpQqyYNAggXie4z8y89MhdjB4Hyiq8ixgE3vsxkbeinB6N2i0x+IX+eIOa9i
DA9LXW85vitsKtMK58tThJZI/rOmOu6fysCAjdpC882pFE7jeD/jjH0/r+pm8wEDUzp3qbBZ1kAv
TClruupoAKhYQoahCjhvDFDXv+VgrlsGdk8VSF2tddgla7Jjc1T1X17UKmoDCp26DC7dgs5AHX7I
QWUXEgSOSOFtE4Y74tBztCpMTr21N/l5DrQnHXwNWz7iBAiDQWZOZaDwc5jkdN/bSmoWCJ6BiGrp
zemdqlW44vyS25UFxPC7YgBhmW0TgvKCzAAQrHeEOT9pFwNqtlYCFleRWWPXtgexlTT+k05qH14z
yiCoNrLNsIH3VRoihc6YRWjpNCZnbzdlv+D3+V+XN6iO+xP/088KU6K1jeSYm4CnKLWTN9H2vGFW
X7uLNXLZ2yaMijLL4OXA67JtXTLCwF6bbwCpq/E1GDIi1aW3ZJ74O0XPbTFgK+Sl1mTZrxi5nBu2
lARsu5+zxj6EtWj+zrIYHD21eF7WlLUqKkdWd8CbgZH5WB9VVA7FTU2H7GrOjdrXVu5pbYWtdXuW
Y4YI3ptuU07Hv16h4WyzAHuOn7xmLCMzlngui8rozUuXk5yyaPJVpun5wYWLP0EoW7pAqU4wUN+c
fSxbYJU+Tt7LcIMUMaxNfy2TUXbdNInjxBTHnZa0LPnY8vjm0bC9rk79OCKlbRtBIgi4hY9qoMP6
GkHr85sZJeYiNRhjctxKbxJWu54Fbi81h0xI2QvHR+ujRbvBQashXIw0Q5P1sCSR8j/7SEz4e8W8
yHv7y2bmlDsFEMDvtB1CET0zVc72miApIShyKap70lSlwYw5wqRsTAHSIbtaxHa/e9Dwecrf1wvY
4aXVQ/egoaREeuH3CauwsCXV5KjqyO+SMLtfLZjzj3OZuMGfbKY9G2FeW6/BQc4sZ7Bh7xlC/kf6
gVLXqbts63MtVstpZlAuIEzxPHzUPX6nRo7GNf8WlP0G1dfmM6YcCUhczhCVhVpIPPHb+zuAqAbj
LXcuCwQsQTjSi6wxnT7L+S7pb8EMaFXGTomysAM6lvzaFYWE5vey4OQz8Vvwpf1RJmTbCC73B79N
wScxOaaTIUiD4h9d1ufIjM8Bk4tlDYU4AFpCo8E8A9yvQpOfFLWETYtndDhb4dhwZnwDxDYVU0vT
p5sf0y+bj0XGLz5VvMaQ7mJSaIi9swlEZ8rjneJEqf4aJyUsuxEhJJCygAR1FGtX1fFFTuuYxPOK
ErrC10QEUhvv68Vm8igXeg167hytq47ivUrnTXU4nrFsyXyH4D7IbdqIYbyTu2V0xg7sKN8wdt+q
cjqBD/Izz2jxOnOK0OpYmRsdzVjvTTZmkzl0UvRqw0avwTKBkH9flvF+l3K0w11YfhoLyuL2CZIN
wdUj5Z4jadVo4hEOss8duCtUpklpWNw7uJ6yd7JtfeqOYVegOglVZTP1zuKSoleHbsM4WQsZvaF0
euinGeZQVBYMf3cQ5iOpfKHg9cMg6HsfA1ipPE7r1xJ8tGEzkrI0QK1cA0qt2dTnZEKNEU0Qfa2M
ykxwnYpNwHAVJxXSLSlsSfcZYugi7SZW1/2mtQqbkEPGNDTIZXKReVYdW6fNj5EU0DfXZ+HUvV9J
/wsyCq8jlqbVJ1+0x6dDeb4fOFS2RlAZ9ju+GWchzeehR1zrk6RjQ1aEJFu6fexT0P+qhLzej9cq
ZME60rnqzAI9jlZnyCSkSwU5gUGHcBkYcV1PAe47SS5q4m14qjhyKHDZMtb+RUkQDFk6e3rah8h1
vGSfmbyBlVUIfxM0CiZ4GZQcLu9+uA+wZqvRMcbSdTmM0FzP3yExPay0FdiTenjuJneac2UzI+xK
bAB0HCqBm7T5etNpd+HbWdS88xPREkt+DY2DmcK0+TNay+cYZjmlWQg0TzPtjGg/eVoozqAyi2DX
gx1ynGWdkVz/+SPoD0UKlcutDI7QuN4psJXfxvTK74XOkYj+BSBtwO04Q6p54s94PzEY/8685HAq
aPbS5qopgDdnVvojb8lQB0ZjRRaicYGc5fqJc4K0OxKKamY4Lusz5nudt+8eF2JQhpClZtJlsf8w
jtAPtrDjTSpIddEm1DfPl4ccEsYyZDzOK6ZL9QYQn3BhnAyTHyjMXowjs7KueOYH6pOuAmhBRuyw
1Chos/mzNunLckhCN00WsKPW6oEmTRY9iJZEPYsRHMP2AHMN//CBr65cQULTQ/SCXdFN1Eoj+mK+
1CB5lHUx8hjWdPfYci+GEf9UU7UkaBFSYPdFRLSKJegCb3ipGDr21reiexATM6cwDoS2yqEzmJua
ARCe/HGW4w99NgCcpTvKAk+PJl8rviM8jllQlraMpX1EDpNGYVipoIVx2HFjLghESblGsWtXmhVZ
Qgr3MzmKywegD//IWDhYFBIlEaLai7di8VM0eALUQDGHFf8ZNbBqB5lay6AkhnRkj5JIdyCCQhTd
WtZ3c4rtrI4NP2NpQnUcpXNA6PgcRD/O+XGbvNxByV0x6PeP0cqSfE27sE3XgVi2hsrheSYyjxLa
hf+0+jQjfHHnH+OoOVBQP0d60UIbdmN0JAWlo+o9uN7dEkva5rvuWjMQZ690UQt8ZyfoMd86KREz
G146fO0/6inK4GYwfqkXAR0tI3atzXClbKqNDozEFirRo91Ca+at3NoFGrInx9d5f7/0IMf5fcLv
uDewDsZPXOKlkTLhQdN2nSkNZtE37JesJeJcRHVDsEUW69vjs/hMQPUgZr9ZfKyUgfRAkzgG9yGl
Pfs6GgL4v1VhmUF167QGB1AfJfNNL5RBSf60fshMj7H9ys4a2/C6i6LmQYHq0Lb3Yxbjkh8kvOJy
eHbTmdD9CMQAFk/QES+0OS1GJ790v0Jtp4twH+EhHIevqaa4aL8R2K5nGT5f7apT3A+w1LlIxurh
7XiOdY/pKeA3mswnLi1SzfWJfKnClHSV7FzOIORyK8FVd+oa5UF0zzhqBq+iDQSci1V+8EPr4HYT
u+SxQTTPVZJXKnnoEKIcBTYAUViazpGxXc0O1kVsEuD6Jd56gTdaKR1Mfe0S0+DUeJCNzJrQ0bL6
ZgRSCSdz9u9nRiRMtdqamgcvRlhZpp91gIvZfBYDiyeKCJ2fFthjGsdaMK16Fj+ZPtd/pxFWvZtU
pbYh4fq9/Gg+aXDTLw/ae39jRcQTuUjOzR8REOSRM/0fcDZOgl3JFjFGB4SUrsZn45QQhl3IRcHc
MCqBgW4ah5eISivfszx7SuYudOsEu0dDy6AfKCJ1tY9CX9hHP2NFnyAHPfl3U8o3pse14fURHQaE
1lw/wRJnQ5FTDcpPS4V0V/O0P06B4QPuJ11JwF9oO7GXVptF4j52f/YTG1Nl4HBcU6r27Ok5Jq1v
ZfDM95xaBJVjWFCW+iLZeq2HgNdsobUHvaVVBl1mtrseIFQwYqeUonVtSo2iHYGGBF0KRlnHZda2
wNGomt93+HX2lkPlHI+MHLSYhqT4M9ZhRAn6ik//ue7aSUao5hZDaoZQ6+frOmzP73iISRmH/+MR
cEtcGZpYEmpu7t6rErUiMrh0O5TUrexZ+UfZKytB0OEdlOMZw0PJj80hMwi7HJ+XdA7JYmzVtXEZ
PcRNaN9i4A7Xfn7hnuyaAKBIZILkBID77+4eyxI9dHrXcgoEPv/ceDlLRJjZdRXRAV4KY5a+V8V3
EP8z+r4PHVefQ5JVGY5cBXvhCkTgNaLARcAAgkmRQ++eHAFGiUYuEesZ8O73t7UoY8/pZL67CN24
6yedTetL9nqC9LUNPxN7RrhkhkcehTAOlwqEam3nClfHt8CYaYRCl9cXIgCUZ6GXb1wLwIMxgM2o
jTdk5idak4hB71W795jXZCUwMyNJbKLrYAiifYp6gc2ylvZ00YxOv17pzYAaeK/s3Y8j5msOEmJL
fnLtOsRZrXWk6CP382htwH1WgzJfTQSqAl/JikGE5AszSOi27MS/a8WNBwcBzYGCHYbevPOV0Dr5
TKgzXt4LcqMVnIDISQ3ecCH73ivmASMm3zPbCiEF8nlmN9ZlgnrvrqZiVDNvgPZYwnd3yuM4/dY3
CB461aCRSLfrC6oUvvaEAFNdjwFKoxKJEPi9tmmPu3BLT8XQ1LsPKLNiRrqNlMEZITYMhywGGq6t
bd7hXI+jVKaXdIbVQ98kSUry/LB+goIFdS4Vr+sB0BRNoRk6sr3kLbuGYCrmxZH2+qoRUVj2oFo9
pZlYhZVkvUKXVzwu0M5DwA7VpAoDgpOVeM9OTguI8tNqjqBuZVmGgt3i2iODtWfsvDwD34YmA3rL
SM8nzQwNR+xpaJVQZSZDz79mXFp7Mq1x1IjkEDNWK+qIS5PJwbYj3CHiQmuPCPdhQYQbr0BVQKgI
rgPIyipwj2g8B8cRCXzE9mXY+9k8UxsOibmIRGU+Hb1Wppg/d8SnpXhTj+/U6XDGsjowmiVHojAC
zp1sgbGQcqnme+/Ufd3gnluqwfHAbeEGbTtLDBQ4xTn1C2Tz31GMvqvfzzmXkoILn8Ib4hsEE8+V
LoJt+f04kzcTmo6/H44eVQozPa9KeHRYm0j42s4JowPair7AyR+GtV2To746OZv2dtsRU5rxClws
nr77Yte2N//1QbPUczjzjWO+ESNEgz1RLISJQJ224nJ0mPMlILE6+cjNrfGHHYQkpK//rwI+Imy9
nA4NETxMsMzZLgdjhUNQOwO2srxTdC+GGT3etJoMHU8/AhnUyb9hp79nF2QcHNj8x4wKHFAR+TPB
RYSh0yF928k+5x3T+hAYDP/XpKtKYt/ii78RiAwqGifRvQaFdRUiGIm7iHnXBA18BrYeq/zTw79n
zAkk1j+stRyp8ytcpQThlYCfcnKn8LWQLwoA/PNLWLrg+SO/8SHdnjCv+LcD2JrpMidS1UB114uE
BwuL+ZVRUasKExX809tFOasfLIYwEDxjbb6EKJilAy4jhOfrW+CSSqKsZGFhMZ40xlzLuLLkaFv4
6lMpE6rcZxuDHpyEMotXnVXaBHGLk6dxGq6LyFxThYUz+MTovrX923RwDKUqmrZFIGeqrfL5pqx8
UT+qUUZugDjSJqbaWvhKstik/BlrFfyIJhdr0YGOYlEeDEBrwJ1xyoQnLZ2/hrOmkVTJi+zsruku
SINmeda+IDd6JhzBZ7kwIPCFN87bKRrYKeMk/iBXGT76/41elqiHuslMidGZhgbgvG+IlLRiWsHS
orFAH4CgEelJMpvveE8rdc8RFPQj2VV1rf3aigKY0kz57+cT18GsDwoMJOdWRm3SYvKdUFd+Rw3w
C0lUYK1YMWbEpCXCVqgCvnOaphC/S3WHVcvekAjRZwenRDY/fVEkajQKOVoUECf+3y93FD2zJ4ZE
kZh02s9feSunkcOb2iISTEk/dv3docdjFdJrSnpSdIK3WQPXU3PlXHUUezNdffkkpy6KwNGltyET
y96kGfFQMjFfH6Su02aqUHeZ75j5Kj00aq6+hjxCZ5lPjF7ExilnvdNgI/CBE1j5iq9jEwP71d2o
N950xj41fFPpkMvazyHPe9iinRcLMW6CCQ3q56bvWeRkrCczhGjOdNRnPcNl4i84vlyXbaCuUB+g
j+w0xoAA1/Ndy7mbE1Rx9I3phhdN6VnDTPLxx+W94TBejPzxIxEI3rq/q7LDfevRQi6HKKtA9s/4
oA7EfPHbin6BMO8yd28A/QtlaKw1yI2OVmPclM7IQcBo0VIICsKxHnlF8XP1rqtGbPr/K3njCYy/
p7u3W/OWk4V33RbZJfzzRxniyDyirTHnXNGLZojU0xCulU17pAPrPOiOZrBjvZWuwaF69hUcr6uG
dx4/+jb4XbPciMgcixD0tS5Nn2f+98+lwCXN2JgZOcwaTP732eAFybx7YvWThOQ612TLIXvsS0jw
/AAEZ0hsFRQw4w4eZgSP1biC+e+yoK+jhBqQBWigUwHOm1IXI1IT/afmdj3VI0H+YmQ4U+P60QrL
eQ3Iz3LgkbHidB80wdx2wfX3DKoTSW6WF70X8u21C5bwg006V+U3XOcrUXgM4i3GhjKOiI480X4/
5ajLWdA87QZCdu9w8Jq31Z/0E57lIy3PKDLiWVMbh7CEfqJi//NFNFfKmgkZZPzMcAI0B7hDSlgY
Dxxjnkk2VZD+5HoDNFL1xWRRSD+sbu+qdMYFv0z8mOH+Iq6gi6lccSx2yhzgV9RFylPGydBmS9WH
d1/+GGyrc5bl64nQ59bB9v3H6/U2q1oxk8nURnB9I1Bnv3Fr/so62lFT2A1fS+CKnkfdBzcD3oU5
O/SvPf8tqrP1qlCqAJi2zkvHHd+Ri0le84M7jyZBZU8A4EiqjGqsXWtpj/HL95A0CBimXRJSJtdM
JfzD9RR7NMYaYp2kws+s2/FCdN0qKUEEdo8HrlXpYEZDxixWOzs2wykONl01+ZFXx9GroJIq+3of
43Oo1EfBlzlxq8GBBn4zekPqrfXUee0z1BiZWjvB+08mciMWOrldoqc/9rH6s3UBxWGywvPjw9MF
bAYRcNIeqgj/knU5QHiP3K2P8D4sVdxH3fRzfebqarhjsj4iKJrX0VcbwAzaJ6sc5uHfjoR6M/A8
zc9VYnsMqK+pe2eiZGPnBEDx83YjEt0dmrcdwlttY1Kb2W1tBS92PI8K0kvUv8jgw9m4hJ3eUFN5
uDbUFCkIMieNxUoQXt7x5gJEc3lwO+MZysnvxweisTMCqoCqTfxyBfMAL4XKA7RJ89rz2/F3K4Ds
UMqE2IwBvygH5OVIywLQbGoeC6RgumSiYA/Qx0VYRRSySg5DO/rFgf2wDEm5x3jlsse9sa5UjKGA
H00TF0D0Jw2LI7aVJNaJBk14p3d2cmwcmxXMT26w8P/g/KwOLlJQIjelZ9+1ElAlzr4pCHDguDSV
/xRMxSrgyWhEdqAwajP2bec8iIcA2vtKjB0xJUqtNUJpIl3Tpm3f5DmHYSo1QOQn8TnjB3Gw+7Y3
9Qi52UAUmxm5KBm4fmLlrs5somN3PpsMxQsvpHW6YIJXUEKOOv31ToSJLuNiM+vDywzz6svOxfeD
0NiYhYUp2Z6UXYhAsiNF/qYgOJIDMMK8SqYOzuouXnp+9UtNsDaBTf9RPTgzaUDeYiHk7eMWPeol
+PYBvy3SMmPFDggLA7cTwethXZVdXUsNbfB9J82vs1DqXU9ielWTI48pP5FDAyVRjxKFiJYPbhVC
AygRXhvD9pGoav6wCFrToUysuFrxaml7xWlcacsRleu0Tk13SpRAkvPP0OPRj7SrQfvC4XGDLOwy
uPnD0JN5qo3LyEa/dvNR7oPxhvyEQyNClBM8sZ6TwZn3QLKlKgps5m1Be+Hqhc2OLMbNjsoONDFw
stE8gyKhnHqqug8T1bdHNPEIMK+BuVEulRPbYiOlYU40Aa+MOJe5nTmsBx8JGpYYWYgxdm6GeLtT
H49A02o2bZXw3vRes/UhTi28SoVtn+DjgTT6ycboZXJLUdylGiy7Y4uhmk2svjEhAuVK5IDD2AnY
JDTSkQ3erYj4uHw5JVq6uIV1xUTSCQ30FcnE1QisruOP+AAn5ynTd2ixxtEkggoCVs7j3DbogHdx
S1RMJHR8IlHWv/I/Rq7s1Yf8lqs19hnvq1lqRb6FC8ySg0On2AGuZXnYKT8YNCm2jh7ZWaHNIhAm
ciG4/yXeuL7oS0VfIj/xrimynIbymgMjbh+5PGwoa4WukgBo1ClFsa8p9DGZ3jwwFe8YWjSkXGL6
CO+I2Vocsz7NjZ/dwi02wdbarzS/46c8jMQj677zptYrsLhzFWI+Qe1BOuHJjsqTeKnxoMdoWKD1
KBqGnK2LblIKAT2Q+wLXnXUm2ILxe2+GHTFHacQ6kHPMLItrOmJvjhJ+pqUNhJ5DCOxkD6+ZyAA9
ATVz9Aa5MCMGF9E+y3OmBN/TarBCusOrpgi7hPsf54piujAqWb2uLV8QniYSme65fSvE/tPLk7Lv
t4lRIr5cGHAKccS/jugZ8+qaoLxTcZOAHOXOxGhknikN3vwEBrzguTdHkNUCd9DjpkafC2q3YYjf
UZe4viZwDWwC0hsy3yQfMGdC4Q/NIezoM0LDMDx/u3spEEnLToG20ZGDt6SAWfOZrE+jbmTnfpdv
RPpykJiYvwJvuoiIk0OIECM+cgJAaRt9nhhCBgO/EEZkQXjkTcF7licFgl4wvoh5kTsoiedTkzX0
g+ICYKarhwQTm0Yc9o75sfUn9HMehz3OzCF8ntNxQRiHmjyoyfeEx4aXpAWEo9Z0h2GMEGJXL9Yy
w5IdnQIL0miu4fbzWk4X9K0cW3sJgwC5mn7+0UNMs27a/Qm4go0ipd8WocfhjdaYl9X8fY5pux4+
t0fmoEhgNdhC7DvXoB3dJ1TbK8IP52oIIbyFB+xfauEeWV2yxtx+drnmTj6m0GuBJ61IwPHyUTfn
h3C6NUWL9BUHQygp3pW3hrLRnMFZ4hurSNVktwbobuY09p8fok8ysg9aoRnGngIANfHydKI6tT7c
ZQImWHDmR/YsJwKjY3qpgPV2cYy/XMXMbuSO2BM/GVUVgiR2UXahsx93SUXKiuzmhTb/R1oZ6o/N
6LCgr6593r/orejBdg5XmiitpVHrYs/unI1iMf5QbbrTeNYPz/jdf5PC32zJDLM4X8sLhWegHUp0
skuEjW5/xbdEj7Cdxqq7xbyAa1GcZ3HPy11t1BK7EF9FsqDcLg83UPJ4I2UccKgaVsw662E2BCxV
yLTLoEcmdAJRgwh0yxoeYpDXPx/uAfcIoK60qCOId9NGqiAXaJeR7FJ/HyX9qtCS9sBl03KuQoC8
H+2cqg/GDqH9+xkhqGOpMdjui8dHf5nQC/LKl3KZKdxlBA77bykGMytQTrSCABhL4ZmXvgNwaYw/
lFiqwKmdVAthZMRQHCuQk7mcd20Q7kkBAq/0k9CTEvQ9UdRL6eRywB6mWQgnmTia45MK4ARHm/DR
3nWk+3iMt6AGHo/C3xBWSALk+Ap4bAH/+d+gRM43+pyBSyVpL9hn8PPtAo0FdUKK3aPTif+xfnPJ
0zaEARCfnf9VBFAL6KO9s/4bcGKkIYk7IO67UhERUqFFqjm9qClb0a9P3Q7jur3MLdMe984G9C5n
oUPoP55blGRos38L2GmyOkm4cF/JnExaaCC6C8SvriUM5gZITX6w7n3OQK1HBGw4FFBll66lBK85
wI4VD3YMlvqZURg0FfayFssH7Pd7Ggape33nopP5pXolSJjTPdNR4bvOp7zPRGrpZwt3OR81mARN
HP19QRcYHRVdT/hqigTXrZdJuFytwybe80A3CCjX9PmVNWDB2IeUSScAptT6GhcG3RW+7ckHUXgg
TTaEILhPdwujxdbGHaMJq+2AGIke9373C50SGJRIhSMz5mktVWtsiEY5lWFN5sJerKxRCWgJ1Yw9
ygbm4dNKuB0bQL8fjpQqad6e7PEgleSmZvJL9e9dm1gVCUSolvUDOHaofY+j/1uLfAE9JaTmDzPG
G4oP8nW6tE9ThPMLCxeGOVF+3Z8Yz6mJo2uSQV/UAz9MnaUwNdXZ1VPmvpbwstXvimY0M9AaNmK0
J3d6HciTZ/DdMEhcr97Rf8QGtk1FFHOwCZZ9B4jBtosys/f+Vj9C6rpMwaVhOuJb1gYMLduzQk+6
PHnCuQsc1mZYTx1M+24KMDXkR5V4jgyXU+RUtcdfogKoVZPVUY+0SikgWjeMkQ8MhKY6x1/94SiN
FnZY3SeljKmwGl4XAwoWZtzzDLZ4VwOCq2WRXAF4DkxKZxrXV4po9RaOPGTLVh1llO3cqZhkcHY6
oa8CDEGb51h//iTf3YE2w2EkoxjaAKosXMzP+e6bHuJWD7S4wxwSp67dTDBBiJF0wV0mz/dLCPq7
TXXyvsBNGuJHW2SmKKw+LiN9yD/x6n5dQDli3T4mBw9hx20x6Hb4EgGQMCV+y5qTwVMtl9jC7OzG
K5oR8BT5o7523m+MuGs4T9CJPoBdnGNen3abqw5QmjmSyEO/eQp6LYrngdkktlqYmMIOlcpwq/y5
PILLtt5H5jPFQ6dVRwn+LaKTRY8jZv3tGVdAxCwIp9W2RYzv8XC2WZ/CPgKBFxYsD37lCPvbHzct
J2fyw/uO/G6mDnVF5/Bmna4JbdITK0hlu0efXNtp+4stOO7mT8BopC6KHUoPCMkXEambn2HG84hq
1Rrc+MlnXBaYZJQ+a/sxFPFsug4EHDy8KHwrt3td32865vA8Rppb3WEWz2RSk+6s+Twq4oI6NEk7
FcmF67B4Vdr8/aZH8v7Ywv6I4Q9dscuQ5BWYxvCXSlEQAt+/61KegSBRiFps7VF+xFXWL2sTUtKM
s17WX15DdkNfO5J3IArnYSlKVOmVOKefJUi4xKcV+DbBJC/VMLo/L8Xhre/PbHyU6KfuccXagpPc
6/Xmy4nygrZcmJBijX1e+OtiNKYpFkmi58BqTkksmq3sX+v0QNQxvmAVGNlDCCAOcXcgfsI2WgQd
Vld1W7kEWl+HBw1gFE3kknp/7MaDOg4kF1Y5UVmnodyobzeZfYuLAQyjmGDNTxKPFxcq7ICS4Rxg
suxEsyqwsW4ApPWnRIeltqjdbSeIHF1gBcmBZ1ICF12z7mVY3HulmKswICpFp9JhPVTP8BXQLeaX
zsYAewtV2wbvI4uaQTD6zFyQBZpYSst8ApIcItkloVkNbxHupXIboHHUufT1t4tsfa0N+Jsna7kz
kUeM9YEE1/mtjcKZyKDrYLJc6SmEL//iw2MSdlIeRCwwP6ySHNmue1q//0cgPSyhhxfxNahcTEVH
Xp6gPLegjHS5TW/dKLrMEEEM+iCFRUhPhuko0X/jGDemPqhhiJbo/8+xuHq9HEW2gU72e+7znkTW
oDmy1lkE9MwGAkLgoKuPTISCul2X+XfCVuS9grN//kRgo/5Fs5vNEdfhOu2kAU6sYn/O4gyCJ+zU
Wyq4VZLhaV2F5l46mZJV+fGAk+lLgwDze8+EpamEmRM0BBQmtCDADs2tj3NZF/6k8WAZPs4w5GBs
gc43EoMalzKAnTmnEaR2ChbDLNsyLKUZTtohBAv17zOnf8PQp95sSnR8oNbyh/wFW7foqLRxKb8F
EZ6bln7AU+NDG26OY5xSVTPPFY/2En0Vvf41GBhT1sn2kGDkKUf2mTyY/iXk2TuhpQejJ50qe+lW
rJ3usYwMaziCkE3/doKMLZWKg3OYIMKBmU6HKk0x8QEzP39AjCVelfcy9QhwFMi9riONUwzvedIR
+F3D3rl/TFpV5QBCM0eQyslHUTKGRmcvWwTJyvZCcaEl/r1ljaHK/lt5LgOelwllHlu8wOS4S7wv
I2bEiKwG/qETquf6964qOMM9hFGd6/m55jTBaXLv3tR0Y640QG6NsXIGtT1HNnjhrE5A3mGlxSoq
zxEdz//fnyVXs63r9LvmAShX2p+TAyR+1pzLNkoEPLLzNze0/yZgr7kObhUrXOrk46GDh+p26dTq
SFFg7tzkAWgSBaSf7lmmR7bNprnuJnuL9gQhJUnllaFKNBtEJ//MK+fSsJHclg5e6c7TY2WDxO/t
9JCfztToZ9x5sb8hEX75eK/IvyhlRLqh289i4PewTFuyDBEzWyqQQ53WiPUFQ+1M8PNRPY9jF+xE
bCPa9hApfNXBxt6s3MgpzP1CUvRtaI6DRNZr5aLH2A8pxO98BRFKlRKgowyeNObC2iOudD+4QbSn
dQCiprlDQFNxu0QmYnAjsf5V55D7jS4uCBZM491no42HrfiN9DdXVDI8PECO61MM6jqnUVZ14NXb
AzS8Psz9YEWydLSUvmumQHC8K3cQKl+inXD33zqfMmyY4C0NC6I3wKvp1yF6UMp42Gt2E6JPnNKK
M2OgNnAdlIM7kVRcS+EANeXcHcy4NwABfHBzRmICneCrOjqSR8CDUdwHjUg+erGFa1m1LTiExkkL
ODqaXz0EuAzecvjLXcix9VtSzjcVWesG29wI6S1keMko4zZ6XrOppraYjnkrB6KJKrR9X7ANh0VB
qK5TMT+4MenGWhP6gxvPFBJFcSl03B3UzRshoDRwS2+Z933Rk3y/VflseTJQiVBvLIuEFiOVfwHa
TBS2yh2bdNZ/Pmcowv56rW7pCZ+WR9VRjrLWArxi93U/1dLLzoeqqWsF/qxNG6DhysDcNRlnNTps
2K3KXT9xoZxroTFlqt3rSkXYzEKZ/2Q0EgRBI19i5CHLhCoumZuikEAyvKP/BvOBmng2Z17CptT1
tg0rXKx2ROLPpsYl1Q+0uRrxxiLAhCK3iRTg1tPkfmODYtsSc6EQIQVLVeftby4m9HB2qa8QDKSc
zKCxYO2ottdoQUt4sSXjLOGrHqBc5woJ1PLXR2EY7vZo9JCtDCWK8gZQvGHajGWp128fO9Z57nkc
7I06C1unPj+2v6VbMhAXakAixsD2GcKGiTtNw8Vpt6Juj/GjfabzH2VjAZLSyDKQ75SVxTCSPvYk
ra7AGnlUQY5cVhQv+BL3OQ/1I59Mi7Fwv7fJl/sN1ddafMqgyglavY5dKFJ08WFgM0GNeFDRpluJ
JEI3h4sCfAkU4kIStLDlyfCVExXJ942fFH/hUtcdK1D8jU3AALmCK7hAZqf7emQ6gfZEuVf8fB+c
6JFlO2hFDPYM+otKgVJ7qxdHbzGxajEa576rSKHLFPQIpnzsTaqAzJoa259CmIOTO6knMbY8DwDv
yBiexEWBK474NnsAMSAzXjErt34pgyuVDiiDhSXABhDqllQi0PgLPbr8dTsbz3Hpy5IpHv4ndNaq
VzG7i13kl7w1ADUks5JPeZm/yed7tSlxDA+n2C1jfMcDVOcbyFgS9+G+MdtwpZD20Msqw1l7720R
HpYPVLfJ3z1y4gzwDm9QBPBc9OhW0DXoSPxoVwrfxs5JamujZUNdVPI3GFM3kTD+uGFaU0qnANrj
gt/3BdEs6C62lhRErrQm0utL2Iyc4A5Il2alRFca2YWumZdu+wcFP+aX03vChZ8sj/QxAh8eSJLn
QPg2t6+toNsWGhYX87L7bIKHRXynFj0daqmRrUkROT2/OQID8u8sPBwuJZALO29aoiu2VrdEfSpt
elKz9fF4b7pVNMOyYirLPMtaVldam/MJ1IZE1N5ahj0q/Y37rv2JCvLny4D/NbyNrNaudy2icqx+
rQTO6998l+XmVxTU1i5d41vfSb6CnN9GLp91EhVK3MOT6pJRVWyAbpBP1SdAJRCRzdw90zYwqylt
HqkvS1Xo+jI7s7bsd/DFwArJkMnY7+ctcgLC0O6qPjeAYMFfBTw4R8xTYIt+csnAbt3XGnTt0Zj3
e5xjQVn+P4i6g1qqm4Dq4beHpAWI7Ai3mCSxMyk//Y6vjgguPwoJOlV8M5Ke1EsbBvqvuWicDO8x
w3dJOWyWECTtEz87ch0EdhFMBfLtRBIylfSpxlhFLhh8M4AWbVWD5TF51JoVuJVAsTRxXzZTHes8
UjiznQ2GVMlTTy0Ct8x1dc1gW9dye2aHXTpl9PdO8y+63rNpNJTGIWaTwj4Xlq9i/u8S8AjIODjl
9mUXL1dSFHgScdICLY8xSVnCC27cGu7JrfEOe35jp8Eq5q7M+U80hqWRnEAX6LdSNs4Wevmpz9Fr
BKfLrwxUWOclM4PNwKzrNgkx0DLi1oOhDvkST5srtmvu0f9bf1pad4BNv0dAllTdnqj3h2zAZ3TT
/YcSBXy0mGFRxP2j1gka+pm4Ry5G2BmUT/mXiI1mQjDw/6t3AsE3GzxKTVxjhNkwqcIcaxg1pJOR
GNj3+n7EeDu2nbadoKY0jpwXIx+SB7Fl+5Qzcg041Q2DII5PZHtmQkH/rAMPgI1xEb/sbEJD43Gf
kiBHcZTD5jRzG5EaJoaYHceFslgqZYr5AwY35/Clhh2l/Lyhl7CN+d17W3M/Av1KfelBNLncB8TI
ZlmmrpTRZuMNcC4iDf+I0nLQeL7huWttnBhMy1OI8BeBspdX1vCrRxdKw0zL+mb/KndOCZAMDVwW
BZDeoMpqXX5fcIjzn64R/colwA0S8aL3MF2DHc1ll0lSu9A5KbOJqOFhS5dPf6SwKT5yWcBlBoch
8W28w0E4uc65Mayw0DqHmTy+mgtGak5MD2AosFeuKikVaqOyP3XljUuaC5hdU/rhVUYpNOPkZ782
eJmI76r3Jhap6Gx0HvjCsgH2Oi5egecbhCOC/ZKh7ugP0UfdwdrDPezV6shsdPCUKuSPiV5NvAZw
Cx2qUY1Jns1nrzcNYi/SmeM3xXKkq5RCWgRPMtcXpOkDoyiaKf3NO39ssIDdlmZd1e+8VP3hBB80
WZPHWC0txZIlIJB9bRSWzYDJtHExvhHRinBVhJ7THXCTio0AJ1DbLrVlvO06wUPo4bnr+AlMl5xO
qr2gl6k6DpuwLvyrZlHtJRCBygd0pJklAZrcWjktsqCHsMPMOSWw2p2piR7UV97io/KCa7FaeAdl
3n2t1MAyCFoay7AebYSgTx1U2C6FIUZ4ExFdd7bdmvPovngv+1/A6pGPysdOFvZ8F4QxAU8Vze/e
Eq/IC4CUl3YYUCa5Sl0uae7LR10jR/TmmKf6RE7zRuw8TzShDWMr7B0GqhlcHcL0z0x8DoAa62VG
4FPCHMm535bc4IBDZ4Q87mBC3Feuv+VbnpNdES41/5ubz6ellaQDzWqxR4C0O0SM/d6j2Z3Hy8/Q
aUWPDLVMaiXYD7I4+k8QJvs95Pl4dz2x5RFbpXkbpYPqyw9FfBs5ONxjP/QbxxY7Jtctzmu5WVW8
Nww7LioEyT6xfIsBCtsvq6Q6XW/rLeAA+WIbYALm1nDuLKPeCawU3JJ2ZD6pW7jTMQf0177K6zAZ
8MKsilwSlhWBFrl8vBdVBF+Dyiqw88oaK+IkoKtIemWtf8kA7w+OHbD7D+jCvvQx9API7xqSorCc
Dn/c1/3PAZ0v2jk5jV4yRSJ8gjjVSF9aa//BzpE9Yoi12S43nMQD18Q+2tNdaWfW6Q21h9h4KG6O
ztmM2G0WGgsHDWuMnYjB2895w2v7hlFy9aJ3kiINCgP+5uM8DF10Z02lUBd2MaTmiDSqpMfdDk4K
O/J4Ep1dh0hezZoAxOtlEUjMW83p1f2t/V6uYEkTwSzXyWf15JxAu1FavulRbwQag5OC6mpp19Xi
2CuJuNGCDCLjJPOxSDSfquTAvxsviUSJdlDDcUzQmeHNfUmgUA6JsUvjuxf2zuOmhiAAh2Sniept
9L/NOOh/X4tDsV6wV92szVi+BkGNlnviHtUhAh62pg4cVH55j4NL5JEfvzImZ5VBPXofed5vgBEo
MRlGusZxYUQ5wf5xhGSbGYBW/06MYa68EvxHWE4pcP7lq0aLTELwOgtetqttea8aPyYXxIC76mKa
t51jCLcrveNb6PP5XIsWs/FLUQLf63hZf8ZR8rqETKAeRTyaKtiWf4kC9Kv3cqJUx+Q/ig5QaD3m
SF/nBBHfHJ06u6790pOscYMn8In3I+Vem3OCxXOwDK5H2tLxaebJ0YFDb4K1i2rX9ygX79o9fDZi
99C9LLGqowALIRIUAKjzeQEmfvFzOabb8tpbcRNuyUnox/kFFxgWaB70q1SBIZcJrZroMYp+4DLo
JZpsHZwTwmEnydHfM9MUMFACyAHgiae0X3K1P1GWoRjDfY2ZUZzN7Fyp1eJO9Q9LldQ/ChtN7oZi
FGwJ4bUtCFj2PjXpl97oUTiQnRkUcgCh/+NHWANAybApsOsqLEKra14hRxg4Bzt4MKsC2+f1cTG4
kZpAcsxP6LAupvSiyOEgttou+bWG3n/7yaJ9IeZgJMtA/pyFXtHrtMec1QB5nnFjbixjGeAK08Jv
voITghamYemGM/gM8IQxkBAQ2KOuAD2z+jCfnakzGlTLr3+vvakDbSWwuMH/2hhQq+dQQyBK2u1o
HPDF4WQ62FYtuw39dy1yft8nKhBDyJoGLGFHK0hJXthJrdcWAMcNXKm3GuIPgCO5QG/TSoiQ2Cbu
rGJ8pufukwDMPC50yK0258Ie+7jN/ItJwO8/mrTju9CzqCoJzDAoIgG8QkWJORKTXPkwzGVTXj0U
qF6A9mNIiHiOODOW8sUk1Mr+kIXMUFLHOcFyH1Va+A/xCBhV2Phu8uEdDq3092JRhUWZ1bn+seG2
hNKDAk8o9jCrKOpnMiLatVDdUcNgmdWQLnA1DR0jDcbGr1lphwnTf96JpVriugCR9exevmzaFArU
Q0JCZZZy94nW7Jag1wacU1AG/F1ebD/RemwbaA4lgjK7OzLj3w0fAil6wGq4KnJ1Nj8ykWZCLvAx
xUoXh/4mrziNhU288NYaP+mKU1VZrWh1t6nY6iEtXUv4my1cxaXCYHIjm0Sow2KgnXIMRqDsr8Jo
0qc2OQvb2HE70XIZuX4Ik5/WLLbW4ufFpYXXuYgfSZvVxENCQG4tLmPs2L853aZvWonkEo9CBRIB
ORQo4nDL2/umJqhsu0gZRfsCWbQ1HSCysB4IXLHDuyQZ8I9bsl/4hNMO4M9po2mJgzmlcU/1fRII
VkLem87Wfz6ioXzeKp4SfoGKz+GZW7YYiSJ5BJ5D2GXIXcIFVE2Ce5AdxeO6q0WZrum1vIg1KCaK
QF8OBqpbOd9+asfl3mxi0WKBy/v4pimadssf7h7bLUARukZFlSLvLIVBKYJALvAujNRq0u2er9uu
0DfHbWEiuYk4UGVzk0EYb960D8wyiGysUe66lcLj7bgmdgXorBbt/UbH/Wi3xzPgBSdWuTnSSk2i
VEZN/Z8mVYrtfrxgFiplCruyFfur7eveBIg79Y2rs0kUZu4OsnK1d+bXtZEI/IzVIOF7OqOKNJaq
zN9OOnvaMd87oGzlAAPKgq4xkICyWSYAk089hW3dZ3cjobo0fXbyxM4VDGENLphVv1Unl/Hympe6
UL9BpnBm5rad5/dYXfvuQ+U5pDDQMvSJ2hfwXccsHleAUtd9y4c9bEhWEk8BFz48aom9AvpFig6C
eqpWwZrocldmY5Ay96t5v+oD+gCMgLwDOM5JvcGb51jgdBfD0gZYkogPaIat8vHg/dnd9oUApxwr
zX1gI1KqJuZRFfLkGP7bXgjPxZKiDy/lpD65iSRgPMWP05w7oAEMQvKCx0dP9gPFt+auN+wOJnHR
fHjX3IHI1SODTHPd3lQdml0E/bX1nrD+HcUy0qKpPUGpDQ4FMas8l1WyISmRoRnNscNS25OxPoev
7Zp9UQWMP6NlS5m5WvQhMDzyWRynST5x8K+3Peon9ibpVSjhBj9RUC5pa23NIIv2BjzYvQ3h/Po2
47qhYhgI5cNA6TUpXBJZmUFpkcFRiBx6cvNUUBRtyeHSJAdY/Y9h8m7FGv95/6TW0cfltpma5wVK
vpURBZBkrRlctg8uJzyQ1ooqDTq2t7W7DQ2vN5+iYEeFrUUjRBaa9VWUanp3O8al+m1SYz7UboCw
aLWUQ8TkihNV0Vl4SAgoCJHRFS/uZJt67W7/HDt09m1nYe+hNMynNJj+9P46tp/9S8swp7HVId0o
ye7Y46aqJERpXuj1yyjVMsVwELbIIlCV8QIFTdJXM4OkQXFAjR+6VZn9xmabG0eh8OqtLs0KNE/D
vKaPsncYe+qsZzAeha/LhqlfhkzjHLcNd7jrHs30C5gav00ZO7znU23TkeJq4Eb+jWIk8popybZS
p8UVnN6l0NoCmywhmx5u28JLrf0Dyvz48OitOgnTdCmoDqw2FojcEJwZqQCHXdsajO4Qfp1GPXq4
bhhDs4EmiMsUkXTd5AMdA5FYhhwbn83gzMp0lDgRy9LUXnUnD9RCa69kLyhwhIi+vTfm6CESejfF
CDTdOP9V5q5G4IJgaV5OxuFXO9XTzMdnPAmB5N+AMUlCQMZ40HnX7xCfRBzpP7GmZbG23t70t41c
N2jCsnTJ6A6QWenhr7u2uUcgUATw8kKno8KY9ECTCw5h3aw9CgFmdt6PJwcq7U57X4k08Gfpdze8
UB/iK2FdcgWkGWuUg9JCm91yTyp1DtyCc/i5IQkBWpWUu3OCc7btcmBjFO+zce4WBrAzLSEmgCK5
kHSmrAMpb88y374C1JXq3YbBZGLdiNVKKT1AsRCjtdWhFsZXxAANClTI9aaW73vY5VwhguKXhaXm
eHo4+jDV+CqvsD2GdKcVWaqmZMA67nV03pvfNlFxF0i1/fY2PpbYz14QwzuZQWYpJqplhQyc7b6G
v/GSjm+7ULM2tiHK/tGCh829OJ6dVUVgZSroPpw1TvQzXU0u6ELeLzIvudSZXdyGVKI2AanNFJKy
maPLhwS88FQE+HmmU/9YidaRv012Txt/cJnlLXVYSZqU8FTjcNyq1vdBwZ5LACTeuVOJ59aD9K1u
NbXL5TzxdFnkt2E4dWnbwulp+0n6bjIH7s2W/j51rlI0oWUB5SYl1L/eo1UWpJR6ZiXsnyODPds0
kW2K9Q9+Se2SNwpfU5poamr2/aCNTocKo3x0zQOcGhBuf8NLTLPcZhUmIvTUfd71dx2mpmGw7238
HZ5FX3UX6a5TZmhcOb0q1if8fptRi6VhF/vTI9LXl8vyVBGLC9JOV1Qj2j7Tj0RKus3JJo3ZYI0W
uYPlz5qPhcpFgVxyn6kC6iWW5InN59RSrNlrHVRi5GT+0TiFiaQWOcBuei6n8QoClRVW0mRCB1O2
TDrEngGPlXrVW+txrCnexFnMHoEl1ffKhTG2fNeVY5FQ+oK58DxZetsRWJgjkhKRFhwzQO8AO/pZ
Pb4BxYH4ZVXtnfKKcMxeaDBtJcLcqrlaxG5aqKn9geeBdRLuDqUizexP7Uw+cui6KggAo0h7UdtF
1PoPF2cBlmwvKsOzEFWuwL9vu7bpedqN1d5BEhVTXH7Iu0l6jucv5S4SFhxnAxTxDB7EJsRPS1fh
wK6N/FbqaEoWArhflaykVvQA6kYd8EyApXQV92RJM3GU1DfWjcPMUJBWuHJw5681mrG4fO41nM/u
xxYVeSt6n6w4APN6odKqlQ+pQGgRK/Z0OZ4v3htwr+/X2tkdzQ4od24wiVwaDUA6/IDLNLL6Eb1P
FStCHip4V0/ynqjQtpVWQJ9TijcJvZQO9Fze1AcMO6GsFGXD7hIM2nbz1KOqNcq2S4I3Wzxz1l8n
ETc/nuFcK98TKlY2vSAz1gf1Ex0qs+WdYQf1BPSLF2Q1C+bS62ftMPx3+3VhX6A7GQG7yP//LzQ2
u1FNHqY4QpObHCzARNE1mJrL8wLWxoMtqclSBGJJofHWDIU1v04Rwcsa/g6pZk+REcdiOTiOOcTA
rn9jU1dz9x1wWLJZW2aEnB4i24WURS55ZMTloBgxGRb8gyBJ2vZovaNVOtV0ugkYZLHFq9FvNLR/
OQhK77zoPMIkOjQazaxaE5ClHtnActWFDpdSvHz2DlhjoHhrY6qbe0GwcTDtMG4O9rckCg0jtKKq
DbbmjC5jjDH7i8CWCNVo+0b4vTFkprEbkMKQlRLQlEFh80eAqVIa0Fxxj4lr/6sPTQVRDo1QnnnF
y2+THpQwAbeXZm0Dr5tR3G5K0QGfI7cxgziIIbg4JkDsctO+weqClZzvinvqVDHodnvg/2ZDthrt
TQiRhyK3OFQr+bvOtYDUX43VxGzK48MWG7P8laNP98tH+ZXaf441LueQjFWlxfhQYr7ibENEXObB
8X9ga0m+pFrMLjHXH3n8VZuN4W/6CM1uTdndJcxDc08HCAkcJLlcrV7qHg3iCpurS5cQzM6BmJgK
ekq7Zaf5hlh6cYCRIMHMg+PdDaSD0UOorXGdjTAO2IqCNNWy7y6jhGZwYPJzTwVkVPxxpXbuK9wx
ZbioRqX1AToD+RBHbWtn1BvFt2LUz5oXhjYssBslCOUl/cAOYUjhzQAZ5DECBab0JeoMuvLpEyUq
F5XWL+CAcfiL1KkjNQDtQuW+spDiB7n/mZTzGRKZCuzgIQ26lU+nKd9AEqXnVMrtjFTQN1nDYdNk
t1anaJ7K852lZGgatpK5h6fGMFj/Tx/0r1VCoLsnaQ6RScErQ5HYJeMUnaVcJIVJLwvCTCkm4T+i
6f7aCuh5gsbMsjke+bHGbqna+DIVF2ew6Hnw/UXOdxnM4bJBFMp4neCN2lVoiy0xPxdcScwLWL8q
zSkonC/OcLYbOQWjmnBMdbsxk18DNn46OO33vmy0jTJIzl0g5mf96598cqhPrCj9TotJHmiTjaY7
pqnaFX5X7Nt2Z8abOjflsfY6l3nYKI5BAJcj6lIQXqWtLlc0y5SnxK8N9glEZgkoSmo4I2LQEKfF
48DnLuuEZzYcgjH7EHXfcaG7OgZBP7oir1SH8EF+c6td3/mlwkKvFTwmGIYFnMPRiqmCJtgObR5x
yOFMFkNrwS7tgSeNgErz/bPgsrmXV9RRBjpvthhXGnZ+GuKG/g5O/D7dXKvH/zw0rx4D1iMnFr7b
VPzCKrYNyzbuQ0cschFdb5Ojjf4IYV4E4/HlWbzWQNoFmL12plRWk2E+xOCCn7ek8NPdZ5bE9YWv
Qa0vLFuQlSVJrJ9zEHCaf+eKk6uvKe3+ZY63hZjAXd+w336Xc+6JWqqFu4DNzkgmMvW77NOnSS8k
xEga8lnFW1lVJuLS7dDInxb2fq0Tx8w9VzJ7qd1qi0XlmT2uhgAhjl+2fz52nOo4n/KG7cvmXYsk
92foEdOhvSjiQpGri9H1nj5fyXYsGrKyqmlc52V0biLtk89eXudmLoqI4oFTe/Rmm7gPYFHWCyaF
udl2jA8kL9balbTrJbV+bwB44Fau/9iWcmlh0/K70pEXhXwLSEQ96M/8pHhT3iNArAaC06PmhIbK
HW0bSHd+j7vgqvGOgNdnkc78zKU7tBWVRhYC9YKaFy/e+XZN46NKhr4YITKFhjNNlZYLHduLL3J8
2aE+y8Ygad95s0snJtvYTHrry9DNHxi2X1KDbadc0sm3+hJ6b9emXdLtO1BkET2dRZXPnCL5mBOl
EDEg68TG4aWsMiv7Ku6wGem6u/uUhto7jGmdDxU7UB/oxSJgN6/7b3/NtsmmsMlTzy7ugXOaxyIG
F3uPFGPtGcx3TV4XOvV9Uzd0KT2nTrJAnGSlFbNL8afHUvZYntLR+i2wxKiDePCwD6YU51qf3VNn
r+SG3sIMHy93l+IUyLEl3bppBP/ZsK89m7bVRSJ9J1a6MATyADZUKb7zuavZKGKdNvxwJJm19qeZ
v9jdU6VpkpgFT3RCJLsbx9OL8NCdZxsqZu/CaATXI7hFtMdC84IWw344JpTA9C7a6M7IYwXARLoE
pOzyL2SvyPziZ/xii9v5FamFZr7gz7xPs90iU2HJtkoOQTzzbDIstbi/Pu1Cc7OOzxBASYqui1FG
muLsFkjFoAt0pvOn0pbJ9qN6e3UkI21zHrkcS2hqYq7hcxhMbHSHSdbv39w+jYy2/NmoezLyNr58
N99IAYIkV8PK4K7rv5+jVecIVLRoMlaJIhelXsKCsg/auPfswQb7HmcUVbpK/lmuBkX+LgoKG4Of
+FuBOBRYssbR8B90OUlMir4exFpHbTVdWe2KMObdTf5zEjOg4+Lkw3kYgi+c/8HO7QoaIU5VcDn9
OO9AyaMMmNPCHUQ6I5KNmO4iAV27ewovu0N3RkXpE3+bVK7s6vpnAdUDkOKYA3CmJrDZN4g3QwhC
2/h2Qes4n/QXsjDHyXXX0OIzJOwgYZ1keY+wO8X9y0Ad03PVWIJnuX+QJEPbIo8jJytaBM5m7IHb
YJMaIUV03mPNQgV+65DZzjHJTNptw3N3jns6V0VyS3SGF10ZFRsyc/yeFYHmfouDQR0uG7gufyHw
RkChDNsI0qIxg8sQQaMVUI+KZ81vfLBeiEY6uvYg8GfppKfUOlByEuAth3Gic8h7zZFbK9HHViIs
ja/p87UDOAlo0b5t95hFGkcgodOTG2ZkNtesmxyOvHESUz6NazZXsTe0jUIlxdryAuB2U0T/URaF
krDFolM28bS72vKWNIIMxNe04RwmAWiRXCIRmVN+dXz0KS8kKDyDqoTrOqxUqLMM67XOV7Mu6sFK
NKSOa0oYqTM3kTyJbYfPHpcYHkmNbtfs8ieDmgHaTOt/ppch7gf6kpdu0mrBZfHSl5w2NmjVxYoe
IZnId9p1E/6oli3o+MB6Cjx3hO5Brn375SXD5m+tjkCZWvfRVptOPs8cQdaGvA65DBWQiM0K5KW2
inGv+I02FgPmBljDmSW81xnX80sqLh/ZWW04qPasiCgL0e5rkiGm8qxg58kyOf5oS+MyVO4XqC8v
u2CONxietiSFOkbmlMiNeXC1/pMxD28Cna4cL0GCkHWQgdCaqdCHen4nyiUhYwh/zlyRMPyWnn/V
cFI+vbYZkYFKcCRW+KCP7/jhLVJjVndjzTGMsbJ1zZM7kvP4t+7GBLMAgbcURon2bWxEu1Np13fu
RizTtxmproVtpbonwPTZTJM9J/YDA8yU6bntIKW33i+iyOyUNKmmQ+L5rjIi2JBLPInI+TZIquyh
r/xfH3Bkzi6JSuNpK1hVdAsZdxm1k0f85oQzCyaHKa8cQvwdw/rDONMmrqHlba6kD/1+0WhV8rIg
+ZAL74pT7HHBTe/G7mAQeKnqPlek9WAxJ9DZ0hjAQsQXhUdkKi6Uv3uFN4f6RIcRJKKYIESHoDgO
KpMYIVTLqHWuttDoaa159g+sAFDcCSMstGBhV3izDcQ4j2dgqCPlTpyiJcbBEsZgRJcaZOLKIO5D
tJt7Uz8aLXoK4rfyqSV56CS0K23Vg3GBXbRQp9oNR5TEEYAHa1BqFE5EwVQAOsPS9CMg9czduV5+
CW6rHVOISaq6Ca1S8n7xfB9Tq4pEOIOlJAB6D9LyHJD3Zjql4+zvHcEJQqL6kvDlWsts/UZiQQoD
6OOzqIkMFMpCsEDE7wmw6iKfvQf/z0YmFEVIUnTspn7yE1GX/INL8kJ5GLDSghtyKNwRa085zzNE
Bv/BISzz6QagafImO/wGynU2Y+R0CTYTudTFYpbzpIOso0vtoe6n+ztNT2JYyykdxdcL3mnbX0ki
YhSNG/vOh6D9kfcXP6lEodVxu6ekCCTF+D28DA6jh3elCS+oVjJYzGDhj31WfyHCEkGq8ubPgeL/
dFl33CxHN8c5s0q/FiJ9aPEk5fOYts8S/XESfCwaFw2ggoyL3NOuA6jw4bU/R3C14Lhgw56XQB/k
lTh4NP84HLpoRLQQj3WD8fQcivZqDhISHuD4+hdvbsrSxu8i5vkcNI2aZ4bF6aZ5GKy1hbsBmQuM
dcu+X/r+SP9IccTB/DvWxmiBn/hjdj2QdwhgwKOnnqnRdrV1yOKVkYKUW49996CPUuxnXfjXN7Ul
FqkitLPytrDFnmRC+Km4B0NdkvYWFhFfaWuNPQjb0pZPWh4/mwbKCkYPYehOXvXTf7PXAbc8VzAB
TvscRkkxrr+qGhUbq6d5G9h4XOk5mrSoD1wzi6VlQ2+xk9hxQOcHjZ/IgyZlI6rdVQCxpGxbrlnN
x1pGr0uEt+CVGcmc7POumb1zyy564W+XUo1IYHvdFzIgvUiZHhPI1XFiHqDRbxy7q5HXDjb6z+8n
zzdXGPnUWEGk9qdIpufkBbxQSzaQOrxkm/AtROYF7bZzu1uODOQQFqXCXdGGxEGeBJ8CaDoBpd9I
SnzOz2z+Y9PFOR0JbwV2xvszA5No1WTgRdj9nwUIZWFJ9U9kuL6FHiBEofy03ASwbq3Or7RpIMi9
VfiU6Jm5yn5BXyBDTWNk/lZNbo3zkxZ/NYKR49jhkifskUKtDcISVrYetuzZeY+MhhjLxkrRO4zR
OY4KCyYEUe3ruO3+snliBnQttaRvzbqFBkl/2jf0Pikcy1Qp3eSG1nEWB1n9AGRkMx3P/sn5jctn
k8C80rKkbpGSV+8Cs05xp9VTZ8XT6R0yue8KOv8aSKG4oV9z+gyG95Pp7Yp4ViXXvwVXhPUfeLlO
cmpu0uryc2YyS0ycEpjOGszC7P4rJSfoJwKmybD2tD5pSNAkDdtAPhKgNnizZycugan9dDHwzxAZ
d96ZXEtftNU7+VdiCuK0wkQAXlHtpbvDOcoeupAJWegZKgVWcpYWHgtphqy1l18iD7ECxDcxM1kz
6RamaH6LztnNykvJ84lPpKdGhIdsYl9zXokrJVmX6LgjK9676p7LVkDyQxMnvdXw3FYGek9a5zB2
Maz//CFtZyYgaONUdZOs5y19R5JEJtisUttvPb3buz1vr0JTZLJ6F/H2LyKjZqq6vL60SLUxnHQ2
yA4p8c6spsKxqRveJPTqPzf5qPySUuI1ae/8PHwZHU5M1v8RODZbwHbl1cAsG6wO04O6D3AWx3gU
6Ak5wfUcrc19ztqnFKnC0mXXMRcahA7xyDbuEoCGXftITm4uKg6IjU51jOGed2zt0YKzMuVvQSDO
ldahkdlPVPTJEg8yeBm21Crc+eywU8onCVrC2/J8y5YaWP+rdFpZGanqF5mXihoT4g9QLLJBY3Pj
b9FKCM0h5W8OioV33CWiFoe3eWmUdBIWFSDNZjDncrkzlVWLXAXbAVu5U/Jcw+LBU5KYCLLecBuK
O2fft87TAhEucgK/5bB6vFHNcwRZ2rxYaVq4isSTheZdQwLFjw3/PGcEDMcUvXuQOYK+U/stpjhN
iHi+YydHEIqsTQnMJegOjQoVfCq3ZMHwt7iGw/WcI17lZByyvAfJ6WTULTS8lZdbKD7R5bmWz+lA
ZqQjUMNDAEu+zgfclmUODUkenPdB/iylnMVIN/kSSpWZTkz9eqs1bcMRUq7BZqCH/FwRBAJSWOTf
oKTpgIInQ57dUigUNcWLEwuQwZO+TnlFcLLumAnPir0lecvsJ1xTPlvGvJlSnvlt2z1w+W1Pzp6g
Xo2cOg1TAoPVc8nZirUymW8OEPlrKLK6VNziOzWulZqBGJigQ6FCSrYCOtCWnT0jqHrpqK9EIKGj
M9pvevwMhYDsqUWzRRmrEe8k6UfyvUwYKlqY0b4Sq5Wc8oYkJEVOFhNPdpsZ1FgJAS3lrqzgiG4d
d/TF/XaE83jK77DNC/dS/fQi1BbZFPsrqabIeiV8AzvAbfwGW+kCs8PistRiAle5VuAq6WZ60HCc
kSn7H2zTYG5BVPChoUMHYY+eNTvjP0+czXdw6Et/MxF9Qs17meW+HG1rRjDRTSIb1eTQss2/x/zp
gyI9dBS7QpG/X0tuKpJ9m65bzbxUCpFE66AqPfrECUZaTjcVcmyOb1Vltv+h6RI7t7cAxdlmZ9HM
n3lzLU3lFdiWPe1MwSS3wAmzn0ZThmQyW3c9hVIuIRcT9uvz6jFcV/79nzh3OFNVveYOONj0GkWy
XlkmgR9kdzgH410vE+6iP+M2RKyaTgi/HJjrzkdoIbq/29CL+oEODl0R8Tm9kxW+gn6XAJAcMRAX
gZh/6+xInW3UXrltQdiDB/y6LjPEqQ+HBQih3sQHX74y2IGkUdMDaVKpEcxGMwgtUIq6W6NOOXMi
zaoLm5HaZDrGBgZM7xXatMHcakaWIyFWol2YPBdF7Lpvd9587laOFG809dT3e6Ktjsh48fFIF1kw
y2uysLcP990/iHfb+1l4BQ8uoMUg6uze8sB9j0eHAVdfnpWkyrIDFpkGoyF7Ff9cFGSXnFcD2Fx6
cuba7b7R+8BKNvSgFLKfzo66YcIOddbyf9+tQAjDqacv53tVzIjGmLI6hLOVl4O/1UhIfZF5Wuiv
2Fi9SfPwO1QVp0EbRN/G/Jqqmpuk34jI7A/0pior8KBd0usjETf/71+Y4E63s+BpNpHXUASUG77D
Ip80qczDBXXnG9Xa0j+Bqcc2hvGTjIr3B923V8lImWPdhwxxzkW5ylKDFPWO3KR0zzzvQkX8/8mF
1N+aUPT1VyQHMGKe3EPZ8QCH+9hxhi5ZIVEWWgTgE1LSXSQrZsK1sFW3Nxs1TBMJ/eJHUij+8mHT
7TqTT2j4wJTuhTJI+g3IrHngZU1svB7sN/gax03fU8+SfLTjQi7a9eEeisd7PWVLYPRITI6p8K9F
6dlAHRGzHyBKaRvqXSZ1u0p48FBvCJdsFB1IKvlPLSI01clEFlo0lM8z/9gz13wHamYYzLtcgstk
hEamLnry/RoiuJDATCbtcesAxB//ZXb6rs+VXkLVDSrrdjAM0v3trMiUGfWitxFe/zfwLdjMcDMv
15gbdIY8nPGTZCHrhm7uyFPRGzOo4GNX5IJuvcL+RtbiXt1HxNxDnnXL/0BzgeHAhXB3l0rud6pn
+VkX/UAtEnbJJZBXr20wewTzktpRo9ZkXrD2V7f+oD5WZjbYOrcBw2L371kPwz/SR4BY89PJxleV
jc34BzX0Cwe3C7AuHCsMmVk7AIZeSmHzZDDVg1KWMRorV+N+hcVHmLDmMx8n3MtG0eiwi8d+oTDq
+bidBpX3ItyRPpOwt5le+q5ZNYwvD9szqY0b3tjYlDl6D07UsD60Z3R54aFH6ywGpdRbnLgEIqKV
HWJCH/N9RMFr4Es5oBK8iSI7YvickPRdbOa+8JOdBStza24jBvr1pX3csYcqMcCq0Zv6xNv7APMg
IDIKDah+ocBIecsIAOIfRAp6l58zfwhBZnlA/Osgeimw0RmiRg/zDpS/ktuILvPheU9ZzeK3YKB7
9swwEclMIWuVVlp4O1bN6G2G5DVDEMMa7F7NmqccCop7+TwhLpSMMR6oo12TQJ19AT/4pgzakXdR
JIYNWmnQzbnOnrj5h3xfBSXu1/xk9EQyyBT3qBz4RPagwGyRJ5RGEVjQ5snJNU2Fpwv3hsyfRIC1
ezrjdDlAyR9amINj1pGjaYb8gb0GZXN//xNk4TLxbO4CYn4bAPPKPQTjetV8vRAc7vja8h4eKdDG
FWrsfOkKKybyIm3MZ5ENF3n1rHQF4Qb6WmKJdMaZvuYdRsHOHWATLgrqRgNJ1A0jnkbIn+iMnBh6
YzB53/L440mnkxJgy0QMoI2h1+ru9PUeDm/CfOvf+KwE32Dx6V12nr/KLSjnewzBMP6t1ypRtKPe
45Uq3ARQiH9QrDfpM2f3YHBLs6TOZbuDT5VS3XMphQEPib/s/bK8Th9isfDkNK3VGZZ8fG00K+dI
Jkws5sQ6zub7q8cQe965ktULzH4NNaSbOgxxTTfW2PrwKfuVq9VZH00tNquCM+a0sUe3aEv7JLl/
13oa3kvuBRDwyD9Zfi7h1678V27aZs66Zk77+dg1kRgLR9QShJYlDlShG8CxqJ45tb9PhLnpoedu
N75zUOAWyFsjRpjRvkxJcTl4M4Wj4jZRAMPr7l3jYKtYmVOPS5OrsR7ZllCKRi3WdusDIgoceDje
acaOxWm9eZQq6yQaWAgmnqey2KAOKxN0Vb6Kav8U9g2EUTfHzK638gJrRDPdp5DkQfaiYUWhYhX6
ymLJ767W5gHrOAejhBfLxA1m2nIHi6Ljr84tkUCv6KMF6/5vHx/Gyj16AS93j28r3G2jc5R3Ci2p
rHoiPfeLfjEcrL+6fHMbJ8saqYxmpXNWneCfmYIlMnbJ+VUKKZxhb3BasjN5A7fa3/OY4r8C7OVk
8VsuJ8PN/fb5MFIskOjHjBARgDhwYUF6RN3++11ytzYfKVPGdIcuw2KNYeO5DBZjz2ejTC47nfIP
rcV832UexZkh/A+BpZt4oQv/CQ+NVTd+8VFkmznfC8kFE0OYO/sGfkASqwaRv1wvp6zwyaIR9G/O
0dYMcpQCoaJ+bW5U7Pv/r8jZ6Hyc4AnKg+MiYguPbXwzjEbv33cAYg1l6oH4L8H4fRcHyLz16Md7
6OPidVAG2aJfIFO+nuVkif6G7bIMg+y6oAgaQ1KgjelZwcudycSszqzVAKUelEjBvNrprBxuN8YG
V458QltcDJjM/zDDBoCeTxNvz5YIQDMSsB9ntSY8hJo1Ln3tqfsoHcVqgalHLK+GaQEpWIi4c/o5
4NSisCH39KoYITCVqVeSdEmxzaNL40QOIIyJ4MUiRq54jqp+SAn2/IP4855VEI6t7OwRLPkBH7Oy
OqJqx33oObjxGvNdBpmluIQnYVeN9Kh+NKL3JS/u1AjSHtSX6WKLjeLUDdqweut24cyjJ1li59UJ
aUsN8+0/4K7n1TLC/fwE2bUo9MRFe63WV2FsT4Dge7ylwHHfkPFQOn3XMJBo+HrxXhJxZoXxd/Ow
kbuJMIwoRKWX85aEynCSB98IiiSPtl61L/fdf+cTDrOpc493TwUNEsBpgkhNpu5NTirS749SMXj7
ES5z5xoNpQ4+2R+HhxB8pXaN538PL6wXESB7qqzieOX8ZbzVvBhdJ7hQIZnO/OPsDsoiN1EtlfQs
f1kiD5j1wh1CHaJ5Dm3V0axgDzEyLw/+L9JLOYSJ1qi6zmLv7Zcry2zEMnBfPkzxHGjIyeAeqrLy
GdV4MmdsWoRSY+VC/rCpZgKCyHQTBClDF4JBzbJ0OIhXonzx4I9NOayez+KkbDZiA+fRtpkOQxN1
SuhZqMkv2BmafTuDW5tdPB5Y6bEQKK3ltSEey1XcMXZsLqKVEWKxQsz0OgyPfNL5DS4CuQFRShoH
8mNwb41Rk9vVALNFSLCSXCwoMJT2U4MVUjTQ0HzC+6ETLq13MI7xZ1HEUR6PK4TvecB6ZJ0U+EDw
EhryP6nQ9ZmhJlmXMHhPon77smWu2SW/5eqhfpzk7cATUNddo+YnE+jyuRxWS/zrxuP68sR1nB0x
2+ie1coysKwOa3ZcA7jEVskds2cADy6nZOty+LwML602LytsJQIBySBU0Cb+v74CdKJGHYDOLc+h
Mn9ybMMJaLwZAL6iv4ZeWMC6NRNi4vkbdMpS5LONxII0nsXmsfevK8Jz7XCXGsDJCoWY9IK5kJoB
qR8WRl+DHp5Ji32lBjtqpxsmQzV7cwVZHKXEZ3pBFmzG1btgpHiZtpuK211Cpt4kNn7hwe5zSuGS
ipQ9GIX214RPTbhpBTgMhtRe7VMLtD/Pb2oJUT3UHiJTVve6OEBdEl6hV9+YPyjk69if3cl0YMp1
/WTLWtPzK7Od9MEqC3TndaztSBl/curUSbeao98F0fZAftUon9IVagsSFJ4TmoPxtKc4DYviDlsT
C/A0P0hnOymiZvn/c4WSDRDVsZrtzF8W1AuGAGqvAz2TzWmJN3VvWulhD+8qdMypKtSrVPc/HV8U
X/f1xsCHZl2/K8FZzs6ttvTxfibIji/bgO5iG3CP10enHuEp1OKfU7c9WMD/Dxe0uBNyS2Z25iv1
TttxSZTxeE0IzSvCRv5WcV6x1ci4mqIQZObldmtYKPxYXhVZa9ZheRbY9nTl4U1duRqyXRQ26M7E
laXUTt+pyAaKn1RF2GCTeVLUOqGKuTuNc9nrY/jC/sNi7WqmOltLkkZ9AClffBkuBHp6NKTr1ZVs
Lk8Vgc4gCnPjYDjFWu1EX2Fh6HxPNjALYDER1VyQPoxgcjGtqMAY38r4rb7HS2MYIlu2uKybkDZZ
1B0xid3YtK5yTIrzhIm/FAas7IbFDdcFJ040iCRhRF+4t1lzjCLnty5D3iC36eSq67+j/cmz65X3
kIbTPOXB3kbiDwhb2QLmeot/+LceGJG+L6/GGBYy9pSjr7wv92jdKvsgdjVUOnENdJilhQL7k67G
6cf/eanKxNTPKsSTm0G+ybuNN5V3qSfz8sWXEwUPncI8j7llNckyRFwN6uLKaKFukPcVbzxRmrR4
l75+e7fCMtsoA6WW2xri0QKXJAt2S0+2VFv6KUkjR/P0s/0k2nG+bFzF6YzHbUNm3Iqc9e3Darfg
YROKL974y4Ev4dILa+9dFlhefBf7O6H+781GRZ1lHqh4SGk9rFNEldA8TFN1U9XhVaFv0FMeESEr
zpMKmCgbECajABXIz0XKMKKKk/Jv4JINbz494ErQT1Xkr+huRUOzUSKTnUxDgDnckGmhYIH3XUjO
3mzizY2G7ioyoH5Xg81MhvcJ3yOQnkDcE19ghOFwobQ0oWQ9ZHMVtIyILfT0De9vOBwpcLOUaNsA
VJo9CEP6b7cPB663LICZE5cNb3gZ2cvZpziLD3+tVbJBqWi82n9H0oi+jgpvmuCz4smXWNo3K7NL
HVO/8Ux+nW9IcXVFC0gM/7aNXKIkp4plHY/oPV2NXWMkJT8hPBYPclxhN79q6iyRWgqyYoXDXS/i
n7bYsoObraLCw12MS7afWjrLeFRa0EbnFFVqoVMHkSGXF7Ba75HNHLsoOJmcHmJg6jMAjaJ4pxtA
tyXUC/HYTZHVzPAJCeyYn5H+AUmE4RXesO/g8nQayTpF/y4UglkA/4up2mlxIqoDLdRBYvIlgiMc
5/3aBIaa6o1zSZKBhjQj3u9DeMSnKDOn0Si6WERXSM3GFYSJ69I0ghAlXKHHzmKrh2eldzPenURy
wB1R8qKCkrSS8r40v1ewRtW5rg2cs5lfh2ZVqZX/ZxX/kdNFepNv3UrpKfLPqX0oSr21ivubh+3M
jaYNS8tNwYLcvZaXc1EkfYyRrQpGPd6CCAEq2kJ2b0BUDE0irmtGohCAW3dNHkjTOv8KVqN+rgT9
nGIrUhbNkw7GFnem07rPFUPxMwEEYP/0QBriVNEQX9gffZC5xjBH5s8VegDZTgINAzNwAqcLYibT
gD8NPXl+54UDMrWISHQ6qxlqtlBxwWa8QyqW4+h9y7a5NBw/bb46YcwT3cDSyI2BAadvCdhWvHgl
0TiWID/i2h3LqtK+ljkjKD55jAYv9tZYvhBXzT1OoBSpOCXDJDniLbo2M7fH2Da4XcyVvicAhg5o
3uSI4UPXLjgPLCBvFPVu1lPXa1Wv2HsgZD0pEkRc2CDFhRHOJL8fcjKIT0YP3HY1KHmw0fZIgI7f
nEKwFxZB7qYyW3JLH+c139NneXQBZYx9BU08hSIuHbM41XrimjA8ckbRh7CWI7dw1wX9ADJp6MwH
adzf8RcAMveO5Tp7L5pTSTD5Z7r8oRLyjU6RO5V82/b4UZfABbbo8SiZRPAwo0jFJOk88C0bqkP8
GMTYLreWGDPrPtAr/g5xc0w3BUK+qQLRl3uqj71VYqEJqbqhF9Bl7u+stBw+eqoLVmymc8iHNEY1
kPjUY16eszlahO6mqOEjXCKUl18FOWGFVPL8aP6ZoIDFTJ1K6OgP+IOsRD3bfHETOSlq0+5QkZpM
8BcBC14AK60SYjfmyjT6fWWDk5rmj1WWzhmBNffRBbyE9MujQ1YytztwMQ5X0KtZWP1DSNadgPYY
MuO2G4cyo3yDjvyYeoip68lzroh+RscneRTnkvCDCkVOL/6ipAMTKbPYtCXKi3gQH/4QYCF+O7NE
gVO2bApWP5kJW2J6fjfUTqj0BZ+3X7r/rsYAt/I72+MmX4F7icEJlb7fWDW/7Wn7IXTGTVXBehES
Kgw6v5ju0dzUpfVrD6yunCpr+l9eVQ4EUaR2pvtmtdOB4ZwCVXgq3LzWF9YWo8AK1FAme0TbvDTa
obz6lIDclEKT1wF2vLkvYK4mL6PDYHJeU3akxQ6rMhC8POKPuXVFGpXGitnE6GsK38iOTxa0kGhA
mki+MxJxXHMNQ+Q2BSjRC6B/jK4uBMFSLnYlUioP+nxrNAqI5QeX1k8e3QoEWoQFze67WUMvJm8I
KycK0ANpWactC8rPoFPjpZz2qsq1QKpnI/mzeO5GF6IgkTC49yGaIcfxl5CYwFd1FGteeKA4H4Cl
YfIhDOVhln3CcrTriTaIp2zLK8MHruzYqcnb1vJVhwd8zFzvpieZA9qUNiqPedrE6Mk9hhGvS2VM
8BaMy4QWCH8GyiKWCnmG28k6k/bUM5IiJ5sJrk3ibJs3PoZr+XmO9aa520gosuqUq02p21Ub55qs
L4Q24UgNW0lbn6alyXDNYpWALDugxRi2JG7L9NHSoYDxfg0JR3cRAVmucRJ5Wnf2qQ5ol8c3VwLx
lAwqi70GDvUiCqm5Q08xfE52wPI3VGzvVZq+leMRAHGDqORHhvHVrtEPJan+a/upxDglU5DnQMmM
jRfLQIhm4lJ2F/Fc1bvoitPu+mPKmEiXpJYGHurL6gS/MJsmNnJbzz3PiZnDOvFu4IhDCnurLpnD
ULsxH2RCBUl1vLYGpByk9KfVATZgC8J9L6C58H/3Kf0oQSFpMQqgNWvvVv8bUrH+QRKFHPblKQSM
cU2rvTa6vVErck4YuLHiiRQuVj2WzOFNMUlacjob8CoZj8iLw5mZ5lZMYz97fa+r3l/Uq/EeHoBg
5ub6m9aTDVrUniHriTC0KRM3mGM32qUISgdnypvIeLeOyHwQzlQ07dMTNBEvw+7F/9R1uPU9OgAS
z4gUbQbtdpDSnr2D6QKotb5CaDfDC7dxPQnOvuc9UWCjpy1EPUxDbxG4vLD3CQcFT3EdfvLrD0UD
dMW5PjKrODXhj9vZbLJWPnHx9tJdRbfnPfil9GIoYdBOjqzBkmiEVxz52XTbumuyTBqytS6aEytV
kNMK04p0f7gnyEtoxsZrHGcqBejh04NqCJHAv3sjl85X1oQUZOAGvvU8v6DhfRf9+ql8z2vBJmso
GK8dRYVMgHntOzYKWU1iev8zof7w3L5FKmakRoEiTZ0E7PwP6W7w7KVoHVnQSoydrGTQmtCeiY/s
RsJoSrAGPIo6Eu54p6RmlOFKet1+Bs09oc+y/Lr6tIxxMD/wZ07wdVIkPId1nAfn7alf7ari9A8X
98vjI4iMHOlRNENJ+I9VfxtwDckj6eDez9Go+4DtFkM3Ubga23Qealznm5em12Xsaq12y+d+c3X8
ufGo5KvWQaVqxLFcRWjT3i2sA+FjfbLWHC+TaxIYs5rpQfKVLk1IR+yz4vRVevOYjKMu0BaN0zno
NxZY1hYG1yXFHbWSF0bVD3S7XYEHFdmBKkBataQ8GqYzdXA9h1Zl3Q/Prrq9IsYR1F24sPtqLEEW
JbjR4GH5Rc1gmox7+Nja23GXHMQ1LntAvJe/5P1LSdQ44m7CyU3PLzpvtDCXP2p/uiv2rl2CkyIQ
6myytHCKroeVHNJV0DIJCQNdO4pm/1kICaWJ58Hyc/DnimmZCzxL3qtb5rXg3tjRDR6i/77q9qYW
muqyVor7jz4QlQn1REWUoe+7rD+OFPcBYKwk4/Ku8jX7jtGgXLFMxOTxtTb++cQoqFaRxFjYcwZY
/6Of6Jd29FkkedVProG5eqi+mBGYP+VBD/QFFmH8h6D0Vbcp849aep1VZ5+XvnruafTkLAJOhb2v
kjkNpZId5XJyQfOER0We3BK5vW7FUu4D1fJUrLlCvnaNOG6hegbNOBzUELLcVPUofgRaXOOucDb4
gI5dp35mhsqs4oFxjSgMRpBuNAk8fYInj+4eWOS121ujbuZgXZTHTwYV79jX0w9iPCYhX2hpURNl
YISwgF/LOrgHVDtfQPpRpEm/aVCobWurwb/LBfHgg4v3QPlAmMY9zzJFjHckSLPgOiyEFtzRuuUU
KMp0u0vW7+J5Kx9RHWhtj55kvbNDyzG+I0qCRBhQkuZ9utXmK+R+n/aW7pnRDOTqsACECuBYMKsP
RMPSaIqSQlFYMeZhrMf1p0emRwQEKAHgnT/yM4qJvOfCWMZz8b2GPQUJjOnh7FSAivveShI3tX3P
PYxhg6eoDnZ9wuVdUC7qqVUJPrFhnSz0s8qFHHmbKt86LBr8sQkQyv5XUXUZNlbr6D7BVOXFW8vD
zkLxQzCJFH5oIfiU5B6CjY58ljWelJfR5ePxUBzipsa8cqacM4bzIU3IjufXcblSpopV+Jo9BxoC
cCXBmk5GJOJ57q4nXq5Pj5vdwomDkS53E2WdMQAjdrfAO6qo9kZcy3qDl5ra1PVaClVPWln2UL9x
ZeobGqtkiv0dRmktIr02BCHojlQjJd7k7mTnH6o8UEIUYCVXAgLnzlr409dTlp4RW6x8l/oOBCli
8yQevr2Q/WVwaeJ5QysiA4yeW0yOUGXDr0C7ZG1QXflTT6jzow5fqO0SZk/p/J1yyXAZ+RYmIwS3
xU7Z926KaGU7znTIbqa4xbBFxvb2y+n6eQLYoJDvfCk+SC6KhiejONb6YJPAZFRVlaz1ebMT1ENV
L4P1KHvlKbYxUdsAFmLKBFlkEAaFhlHjaOh6XfDPlAotY2TJvSBNS6F2nwE5tCSqGHhpbSlenUOz
vRLUYbkpQ4cX/KPnJTg68MTq6AOBgrW5UOIGA+qPYdoOgaW79F6MBu50x2r0q7HffkwcwIVLHJxp
SwYVALhKqg7V1PpJXROx9+Jz7KsZ0teiqVjAWUzgQG/wckM6sQLt5mrrcHuCosi4cVajPOkRftNo
oPDoWHMTSIEsaNf2aX66dynwTrwE78vajYDgpZwv2DR6mHalY0YnkKobJZAnH22lp/I9SGKkS3uZ
0EF3ylu8Fs3dahRD7v3Fty3qXX3C8fAzRoaKV/iFQbTw5zjELlGJORgiXgcRaD4o9PCc2dKjrKOb
D8b62v1v7XXZZQdP0ZHOpVPgKineFdDqmGwlVRAkO9CVFScvty/dLn8Jkzk4SinwL8L39OMt2RIq
CFuj60KgX3P6YCiXkns98pc9Gi22q0HCiok1ZN0VvBloz/bMtLXK88786PdWDfa0S8dDaJ5lqCqs
BT1aZq3evTNh2UijecoqdSgeWpkoDRvGf0wX9HG8nNflZ4leb75RdvbCeoPBMXyDzgPpYbJrlRvV
3m+y3GS4+xfqhUR+GTWb/QgPe+utd5sv61FN99VKEf8EPM/yxv8llXLktEK2HldR37HyaIyJn2p0
D3VVqcv9QLxZuOeqHKhJJ61H28z1J1vjeygeLGONtieKDPSmxExv0Pyk2nZeO5bbxhAeEaEMNboZ
4G3iS8Opw++tYsl2BsZRGYsqfDQ3SdRvY3WCvX/FksnjPmL9ptqVMQK0WPmUByioXzMTr6z1FHOK
U2OUJ76LlSYdBZTRIEzSdS6JTbIzyyvkSKFVLv4G4KIe81SOiB5nnEmWmNppAKAuiIbW5IJ7wS1L
HIX8yc7GtgajD79k3yLmnU2oMA+c8zkVYq2KpNJ0fq4CsiIz16CzcUwWuPbl+t7l9/ZjZqjJsEwq
1LWl0DKum6pLTfY3jpAIIDE7oVtIq+X6B2NkUzM/xKy676wx1syPARoI2PiSLE4ekUMvWYGL0IB5
LW+v3k4iSrhRq5r/HdzbDLYUHBI1Sn8gwX7ZBQXbFEvnWArBwVs7BabkmO/Npt3v8lGJCcrep/Gb
+TzObKAsIezNT7+7UZwNnE04V/GmaCJbb1oNTjKyYa8GN0HmivCT1GmgO7cweREqoWlAwN1+iJfy
lkP49Ce2sNUw847YkSpxvcYQX5KPhm3VpL5UUFx20ssztHtjM8qziRlvGVeVgmtUyfyuiNoWVc1d
DhJlfHbTZ7CGhNSXjkCL6rnRE4D8bS1dbFB7sAcihpIxdyRrUPkuTIbSphgSyKeJbEGzhETzC6dh
DpI72gUfu5Erce2XWTvPw08MjtTQ3KWjqUz2p792xxyu2VkTtfP1BcqiSO4cfyH5bYUUgcHyv8Ck
flSPR5T0EVHjYDlFkWkr9pN99ZwbfyZ5GChcjJPVwsSg63GgXCrer8H/l/YQnfcB19reXSPawWdE
qIdH3cINYq5zu/9SEnc24RwICP7ob/GKUHt1wEdvP0Af4CWxYWUTExIy7dZwNIKu1ZwxigLU6LEh
zd6QZdGm04DAOtnXjAi5XPgaLzg+THN6rFnAzAIBXlbCnVlFn+tg2fbkotfF0c64IoPw+QAT6TFh
qJcMad7KsLUtc+LIU2+hr9O6M1Zzn/6Y+/Tp9UtAlwRXJPtfhzyqj5dT8A6uXWuQDBrH/WjpkNGo
FkdJgGimMsiTrpRSxBKJQZ2CcqWYDnYeaghAvY5RzwXkgrET+a0Do07pVJ762iUhKMrpJGjjuJEJ
emr8q+FBDT+r6c6k8YVxyRhRsqCp5SeFbBRRhALGqw0+3rdnCADLwCE94dMTTn/x3fEgQejmUtIq
JBnRQBPtGlW7GX5/Uon/B3IBSzTg69d3Kifr+vd00NZTexxJk85K+lMWdWx4EaLEaTDAUjtEQmdb
jl6TUxsKtt5YrC1nkpSJlLyU876iE8F6E0b7Jv9vXd0SSb26H+3N1ocVvxBkC/wZdweOap8vtRlp
8awUk4BOZ3NRVfuMGs4lvIpwmhRFbRs9OcbzpGRKYRHJsB40QAKoCUVQUp6hFgq8ZqXDX0M0l5gD
xPsmp0Sx0WgKU9EyRRa0pP4zJKOgYdRnvb6WdELv9PHYcT1Lsh/fzNPgHpjd4mX07/7wb3wmf3Hd
ABmyq1mErKpcj2/saC1vmUlN0OG7M0SDtfXn7h1mVjnjGo4JUnHtT5k6g721li1B2awKv0nGtEvT
u5PbdUx0ECR+MzhG5U3k7jww28snVulHL2PnHRVdhh/LHuT0vsE+BWGWS7LiYoIva+PVCUJ3Cjo+
6UsuGexxeuo0flg6Xf+M1Fdo3sFUunHJonOH+VADDYtVe1Oa3tHI4ql3HOsO2AmYArAGsY7RLxK5
DTG7vO0ACtLuUqO+tPduQgse4LsPrbEYIgcaOe+TuqgniSxbbYIa475HPgwwiqVAyu3W0YE6mSlL
Oe01GqbUeGVGHJ6la/yE+aKF/mo0G6AQ53ChFojCciSZav5OIRSxEK6TY3MXm95YbDPEHBkb0vA4
qzP8ObLkSdcSuFecreK+Dxc0TiDAYRqG8QF6qII7Zkgez2mNEBcKLIYpK/HRQXyxw4g8pv+l/yH5
S0oyybtEuz4DlBaP9yjeZkA2MbN2DWGRQFFy4SPrGi9U6bd8ANUszLVLIKvtMtU3K7D4e5FM8Zdr
ma/4uvlK91RdLjMaOro8nG/TIgm28lrmonny8hqYhfsdh/pmZh8+YfRNvm1mluqvJvzHtPJxCOGX
qH0/sY81EPPaRVwATib6lH2/u02MzqLeUKghTwd6zP5a3v0ATGfqJpGTmf9A8ZQSVoJyb5FXvjsO
JeuW/WcopuC7D6NKjR7aWu+na9ZZwFRA/YKcKqDnPPXm5C50+N2XTByUOYzqmulWTcvvsN6oyePH
lyUFB05/oGMQa7GhoyV3kTNjFNmSWMibm28xla2BNwNj+ABPKSPAa50KYF7VTPu7ex0+NlOvJsnY
cJ2do6v29Wwq6mgzN8SzMJuQxsijCPDgcAClMWOHONdm86jOciXDV3+3FjvOJqNy2BCLqatt1lWQ
N3xIcQb5zCTM817KEaKo381M70B7Kgo/yNxDQqSFFLASQDtx0yyMTtghHKEvv8r89Ry5sMOMVn35
9XwhZrMZ+fPmgJKvxBZJ/IoGNNq1+0tS0Gl0msFb9qvLropC1J92MzqqT12VWoWxQOvJ4gBL13lC
ZIN8valo8sMvWJFgDHZGTvva7RpgrdH67cMg+ZmGxbjEAggTfJHQwljljOl0JAQ5XS7OpNYfIVhP
vbuhrqxz361UIjkGlQ5DktIUgVgRS3rRdCLt7q8mSmkwJvNnWsNnECjjHC/Mas8dEjtIRe2qJCHe
5KaYhAhYw9uLNMPMiYzVWfq2kC4hjRkuhH4W4b156LhqNr8HQk8jqEwzbaoFoyVEfRP3fs8peJz9
IfsBuSqaezqbFBGG7WwziPKVOxN4rWNgKue/LOBTxerbpEOtMQ1PLqPt0+8m323QY4eSnuZinLIu
xvJiF08gkEXCN4FBOa1aAXvsWdJW58BykSYQeebgQIpazjPGRSyf04hp0MgzWbbkFQ7bz0vtSqGg
owYpoytb9BAOmtN2K8ItvsiNzlLG2ZZwzfxlm3zd2TDHMTaIn1H9dtoynHVKBSTCBa3Y89nQPEZp
eUIVkuCsFkYvzXtEkCA2HYqVqY4VpxqQ01kHQo+p8OcG2GIarR09L1GSnTpsjiqdKR2Xj7MxmKdS
2C78jdjradGm/rzyMSQcEMDfdKf9D6wkMu5245c2Two0nyMl71JaPUcagSAviL6volJpC/6q/pWL
8xnqHKf/g88h8E+sOxgryHqanN0RyQwU8AWgdO5Y+ijwwwnveF9PlIEbxLkfRSNU5Y1TVt1KGLVz
yShTsglEQcCRKUrLHJ3VfWOfiZGdVw3XTx1Jiq2OoUZ3qT2DuvkRQ7MBdLh5aqjL51UdyOjzEAhD
kc665UqU2LKKKkLfls0grBVimcq6PZh4npBf7enejHZ7dqbT9d8Q4kxJqYqOEYTUr5qn/LvbwINP
Z88ebpaS3c4pPWPRnpenHP4QxTGCTVc25ze7UZwCgQxiS2FA2Hxrp+0xIMUER7GDF0YgB9Bv37kk
q9CCtq42WOkrjOqgYvvmPmW1bgARnSgZDJRoTacVXlba5tdZmMAlT7Lg6n/3LKdi0ZPhDF5QuPXv
aarlB0p9YDwZxV9K542IqgKz/ItC7igUGMhGSGcN7QJRM1cvlRw1HgDJ+jxNa66PZaNyLDYrlGzZ
d+SgYqUYdl4c8gl3N4jHZPoEEOpGpRc5mMWdxLYjWlfbKZCrHK++wUBQdTf3oR+5aZBP7R3uMpUN
drVp4GOIMJIF5ksOIsJUMmzDHz5ZgPj3j309aGp00TWCIb3BOikdG+e4sjhqFV91rBPJeSwvUlC+
t0cnpVqB3NwTBvVA3/edHGb0wvV83XUu7ADLUJRjr1FpyQqT9xXrWvmDwsTawXaYyLdUN1kJUpAB
44E/4UXsv02kR4w891/9+8GKD4Wsik8+qnq5ReDn4AVfCrXDZgFS9QIEIqJCz2oDg1qU6CJnJRW2
lVHw90x5/WgqTAkrBmKDhHDXNrFGrCz1uGw/HGCvI5MnVglxsdbLPsuyjh50JkmI/1QnpYPvevtL
aa0M0ftqfw+Tjm8g+la/MJw5VNAB0FATui173tgt5BnWBhrLiOY7/T2B8PLFKgRoOPKoejid/HrR
NlPMTADalItriyNkoFntecE8tDDzL2CS9CicARXDomIyUXoSsWQx5ieRbXnYWPsnK7oqwIfmL8pB
D2As9ssZdUYPYIIZO1VLyD32+xzJ17gGzMJ3uNiMAOiYe1aGEnW8WWBR9WocCgDcGPk7KdU9GRT+
J1PcC5HhSVcI8rS3Nxnt3ORoYgD9yxUJ24lgrc+Fy2j7SoXnc0Ki1fFBDbSRHtr3ykwAAhep4kWr
Iu1yvqe9JACNt3czqixlei7ViibdXiMXaP85cDB0DfP5NlEyeu5EJ1VCNZDsSqibFJ/YtjEXL6Nf
0tqr6aqQ3CkzGYBaroE8rdJNEEuXLLQ1GDQGx/990fiIhPvAS7iCwLrrXtDbytly3lhRo0n/byyT
k+D8JGKXp9r/g2qWflDQmnBbFroQVHMm9F1HapbGw6Pbp4JV5u9/SwGvTS4z4pkqsfON5qU/fHli
t6AxX6xbIVmdmjphinsKU6xOypAihSp/BxLPlJtS/LHYTjJ52fgUpyAKmrWugYWdKT3f+BsHCRut
lEDwpmydEjHzZR9IUvZN6pwuYU9zVSU+kHnlFPKOoynaVlOd4ejBlgb1R3rlYNlnSHAfuW6SFo38
9JNxq9vgIc/JHjZ6NYnCG/MWQxjybXBg2GPwScEz3QnE0J2lBqsDBnA6jIxgO8/EY5jqVGW/PZwM
uNPNuqCf0E7M1eAzUriC7hz7aXedX/JcP8ZfZgT9j5E2LMh/LSu/D4auBWdFaB8TPXmTGlvcIHNx
pzk1t/7C8AuKu4ABa7shSVl5A4K0IMg7LDgCN/7ycv+/1Ux8U6+l6YuQmSXOaN60atH0Q7mMIkWm
cfjWhBzqZak5lmWRpl2UPlrkitQ5GueQPDeQHKG3M5cWwCsBJ3SOa64ma3fxpeyfiJX6JQrGTXgp
uJn1IvgRAwxK76NMwtmipRw95r36597RNb5iKhIhJCgZIE4R95hKHsq4+fxRYNXLHx1dAsuH4PKx
TBJuaZ609U488zo/SmtY5/jvp1af1F+pk7M5T7Jg+jZE0WldrbT7h72/wyoAQRQd1ijTzVoYGsc9
DYUzQ4pazRp+iN+e5cWRWJBx75HhFAjJmLxm8Gg5rr8wUu6Eq2OaOuJGUqvaCbhU2IyNjFG2C0wf
eOST1N/5azSmxgZtuccpOle/Ylz06ZlQiyGYwkSDbpRWuF/+QVqGdYUwfe5dFwwSQXYzTSXCGRop
iyrgJ7IGPDQG9RxXwy5AtF6shWEbHoHmI9fwuq+AGM/MQUUzCpNQO/Tj1NmMhCfQdPo1FkiOV6IZ
GQcrjEuB8KeEfwNoNcJATJw64YA6owJI0Ous34PyCnBsFHeNVkT3Cxx3ssggN4gOVePx9nhVzrxT
vtPy7Ypzt4NFKXD8ZyVhFU/W/b7zmWQ5AxqTnlZfTfcgGg129o6mLJfuyr5KfQpoUsIdPS9JWMUA
xw/9djpAPJnCl251jrvrTwd3l264qDnKMlL5/t2OLTZ39kHHrpf3j1hpj1TsSWe3j/jeXyufT/ko
6blVv4ILULhV62j9lmWjBrEp/vdEGrWWsRDipF5TKAWrBJsAav2HHWScbF0o8qsxfNH/xy6yqCqx
1haKX/k5VeJ9kXSoLLuGwIZSnBKkQyJP+3JEJWE2m8mneSdOy/JUcdA/lQqzbugSgaWDAoM4tcwe
gF9OjSO7R1lbVNmdHqvEO4VZ3soZYf6zZDwE0n/W/2SGsclRhivUQMeHsDDTuwAqvJmn9wG4f0Em
91cbjWZsVk7cYP0E+md+Pqy6MwWcxxIpIe7mavuFEaB7vatiCCB10+MnlFTQQIK0HZYX/YQiVspw
oh116U86kOZapz5rlV2VyNlA3x6Xk8JtZ7S8+/xFZ5+6u9nLTdbBvdf5mPVXxCIDHCTh3WT9lYET
XPQAUEFKoFrN1O+BQwrt9DtGRSItzuNR6n4xgR7XDCreZR2LDgLn9Pq3ChdTuYhGmep2y6Zz0epd
XR7pz+G0kMzquJpPmzTK7+91suOgsIO+rbR+vfMPL6dyLc7oWhjVX7FXHJjwVQIEbMKp6cuRUbyN
+YaBSHQpMYj/NaYhh6Cq7lZVlHgYwk2c9v9EkJA/lTAKh7f32BXLW7Rsk8OFqfM1AJfBoqFRBkBv
TWfmNRTVRVKXe96b3PwXyX6yWO8CTaA9HhCdzJD/j+Z7EMDFBI2iEeVy1hT4m72UAPNcjFDrItPh
SxYepjmxxdbpgEH08ca1hVbg6KIjuvszEZlSzVmipQ7KwTKiE0Nm25bVSsJYMC+rFD7OPD31fk0B
3ooLat6oy70MtHBj+brM32wQrI3hek9M3JumsHzZ8vU0iDVB+PVLdDVJ8JM+1cMO/JwZ2UxBLXsy
2VT/NbGY/u5I7wq6jejZZMuoqNpeLuFxQyMuaPl90iI2o1lPMwaeSvkfBHrncBNdPt/fm0LqSuQy
sJkwfBI4Ygrjop1YZt8cHwBVGxW3lPrqbBRYdJL0v7ezAvJtXE7Y6YIizUVGaswVL4/CkzfOffdn
rsEvYmOQX4aGrlyv1oIwcMku+YQctrdLnCd5cKPuESMUgMbrhmE4cFBVYF6jo4rahJMxrffjNMCE
37+LFpHRMPaRMvuIWNRPDhRKzrHUiwD1/pP8gKgsNZPshUhYYHsKuVRGrS3lMJaKcWpSr67hdkur
N8SfwdM6acAdHz8sV5EE7bvF8VdyoJXUqq/E5bUTZ7f/cMIGZvpJP6c5XdVaD5O15dwymQQ4AC15
2LG8t7ZB4b2uHLc+JVrPnrtTIpVCufGggp7Oy8iE+29aJAPb7nwUiEJDJZiJqR8Z8gvEWaQ2dKPg
rpDAbj/I+ca7BsMcm7VWWywFCbhUJrq7whuHCMbPc+ZzEiZcZi2R+q2+cx9yCz/8ZAjb+fuhIrTi
0WnHh5njC6DzrTc0D0U6srOaCMGHPVCB9ZAenaDfIM+OysA0sy9Ny0HXMkg5E4S+9L7hksYAKoC8
ViM4E5foul/PNRkM5nuyxMuZ3FJlZ/2asCwmb/XecEwfgCNOojw5JBZP9AY86NOIPLRjaVsUvfY6
qHpPcjVYAnO0NHAMLlmRTA8W2dVhl2ri9vlg0383TlrFHXMBalJn+AdVxoSiVJ8V0pxlWcnWNuh8
aNdhaYOn7IWFnxy5rqMKp/3ElmHk9e6RpHM6dDf14oHU7CPPBYFXlPGzxEEjTf2g03BD+le9sH8U
2uOS2HVSEv/WtYUYoumVLhKMzQ4dS0eG6n//RT7L9i1hkgRmoP2wGl9nxWUhzgxf9wJatMXT34hx
44bmMdzKELGoTKmYWdNwFD49JnGCmG8CgsFrBN5tavk5YyyumD0GIoDtIhkhM6VktYg9iE0zrKc+
LOuWDjP4e5G9kYFsnRfP53trH8QeFrKEi0rAhzPhZTBD6zLNDCUQGa3aJzt0ZaKEVPHVrZPnVx/x
LjgiYVwQ66OIfLyfiOaX7o++Zt4XbU3Uwv4Non/UBzLLLaRnA1R5af36h+4thPU0opHqvcow9A/J
cVxwT1ze9oD1Ll1OrsYOezhRqTtblRU6UboE2I210L3YXi9SbiLiM2hBG4g8K7g7U8gKDWZvfI5J
Szv4nF1MMolm/cCBgR8/iZ7T+jtwbwsdzuHnoo/MduqnWn2o6mkJ+Sb3ImO0xj12l9N6HQRk0zbL
F6EETgTpF79qZjtfCQ7Xrb0kZ4tWnfRngM0b11N1FJvT0BaLDyydaaCORoCYD9ZM/y9TI8BDq7xu
/sxQkXnIXohqyphBZTnmaOqLgc2WkMvmsHICeFp5TNQTtyFmCnCoUTKdz7Q7HLqlgpnVnj7TcrHB
t+tNmOqlpJnUBWSZ+Lv7upxlIF9nk0f5nyuniYZByiEogGadqoDd041lpgbV0I/MGNCBd7fGs9zS
PBkZ2DMNlXmFMtUlEThXMqhP/znuTjEJDYOA1G0f777yhZdlbarsjfzGWZGhZIdMh+B+Oxeh8bnn
Pdmnok7P8RokD0mH/eptTjMii1AX7tjzBNeA5ZBjYobXIr86b5PZBxUSOYg1Tss58cW0WGOIbRu6
XM6uzb+DeWQ+PWJbMVoXko0IWz/s0PNlT+VILE1fqD6AZdwihxFX4JSV3ZXC4UK57ls51GU6MkER
9gsNVOlapSS4UtfQ3lHiBRZtpn6O5rxuwzti8xLXDgkY8m8OWDEmeaZh/INb1nLvIQQmVDLbGfkg
xUHrpGuKANxudadtow5RnxFsf7goEL8r/R+F2LuL0MgX4OJqXMB4OaycISNG0NGQCU/F2pt5rmIH
4EtZHYRaFYvluIKOekhdgmiDNTkXdcFYMylRIXoeHFrkcRrbylXcRMrhC9QprnDrOKqSjTmMLf7E
CNgsuuIMrictAtILyPgTmBNz0Tr0GVG+0xMkMuQv0izCOdm1FLm0sJ4IWhFmB6/fGhM1eE60dNa2
hOYKe7GGI0PpfsoAZboDOFBY07JKldtQH7f/dVtaFc0M1GUahhaiYWVwzhl76Q2iOFbXzMOtX1ev
mSdWkz6Huz/OoUCn6r2/woBkILk/SGp0nEvw4nTdYMPCF8s/nTQYQijvWjJKmp128a6uVpUl8C+u
kmKT3HsbSLi0Rr6NxbKG3RAVJKynmfBJfrsizbujBt4VVDRL2FCCejUqwokBmp+UWrMXHPLBMx+N
5fkqwv9NEKxfY/dY+uQeiT/YV6fdNmsnahsXssabMT9oh2MmyG+YdR6354rraR1cfyDC0dHcyxxF
Lw5O0I2hY6Vp5Bs8FMq+Bg3LeViKhQMQSj+yTcDOFDPovqpevb0RRn9M7pULSYVxsiO8ZmYTdfsJ
Nxhrc8wbS4/9yFMxdXff5cQsE04aMV66tMjwgFbW0K64GiX2PR0Ue6Df1PKcxhjhBBH1LVcCYN+E
H0ew6UsKVcIIeKkgcafXONmJ2dopnmngFDEERntPjke8wIpJvJmHbxnf8hX1/aCIJzkjisfYg6qt
TXEdA0oWBp0ZPSU4/10FPEkzwC1dWPpRUe4Fh3ryhJJLSmfCkvf5ej1eA4HGf8TsXEdS6VFpsrkW
qJYNVR6nk4/lgaabP6ZQh9FiKG8Pvg6vO6PVHsRRqBSCaSZw2IJAfpco4WqGeOPg1ReF96fKdGsK
AHX6pjMliCBrAuYpmVTX0elKNxAWVTVQ+twpTND4yEVxNI4/nwVyVfBR12xvy0xds/b7Ib4nszhD
iBMzPfbdp56QEjoCdWls/rCdq6bJwYHgOMnGqhWVPkefbYM+1z8/XGl+nAAITY8rRs8zv9/QGWFW
qo6rqfwjkb+8+xwL4gYR1CaEFhhT4dLOTE1LJj8UEQCO1AOPna8q0OYqmm/Mkh+BYNdYFeSYrzNy
tGVNRg5KrM0p0AIQuwmeHjfeaaYmWz5+4wzT1V3PPrmZXvYnLiwsgF2OBgAO9Eqnk8Qz+euNDmf5
8JyPT+EutCNDGZ0+mOrOsXvYvkuf7S/SgNOr457HQZGc3UQ+VC06OFFE9o3sHJfD5Ox+4jG6fSNu
6tQnizPcXdF1lu+cFiOMMUpkVxH2qwgJrI7N2XknNJp+vUkq+jcQIVJF/xHlfWKySEtawiCbLVpo
QGsPWWJULcifgs8SfVLtnVptJs9+vnvSg8bLwtgQy8TnnslhrhlIvRUkwz+ovrvJAEB0HvBbfXTJ
jaX8F514blTa0sPD5nESx5FdkGJOIEAHbpvTCjbH3gtHBLckg9aLeCXybLk74iI16wOLngxYfHaN
Wy/oVhJZrJ1W6gPhHYA18klr+7tlugwlXlSHocfVA+cmq0yi1TEC0FLMD7UwAAvKT2Em8QQUOWiG
ZKf/GIo41WwpzOzdSIzMfYtTjEeF1vsV863VH9XvkQP2S7X2kATkN2U+s/HIETXkvY4kyyU4nrgR
V9qybGcNCNUfVP9eaxXkB9ERPnoOuAR38ivOmbCAW6pVZQKAuZgMtD586GXMrQNZe7Kw470gFpmV
7jF/ZjYB65h7ZaEALAf+JTXalCJxBftes8tltby8/9eKuTV1iTgui7rqzTpD57vi8IVLCIxx5qUO
1MXgzoYbYRPc95k0mArJre7A+ax/6dLez8Clz4RKq0U9nvYpNsLRMLKQmM24Ao9bebIwQgV5o7GV
zBGQCkMAQniIdhxIUgTsQ8wlKmipyzedVGB1dvrzauCcADwC10i0qJSPp7UC0Zc+K2nzpVfBD1R/
hNVoJYetFu/uMaU1QDy4rQUeIHXQdOvTjL/Rs7N1SYCGBH+dBd6zks/mDZZXffr5LPmouMepIqge
auU51mXk+wXDthiPom9XkCfCELzfRqTKzNQflUtbQBfxwE/bT8DMXKBVSAbkWKmdRgrg1cbtMcI+
NkokMerY2m6IageXDkOCq7Vw3vVa/UlDd9rLkSooQ1ynpdE2zPKm4rVk7iqNf78EJbHIxU0oJx33
GzrtuPg6zAKh5hpi8AeT1P0IzQPxKa1N3k7KfZDG/cBSV0o8f4K8dgI33dlWz9j6T5Xa6ylekhpV
OMvVdR18lzd0HiUsKYjGfZlJvZIwPyS0j7nh6nlwhdUAQrA+4x2aG7s7T7UwSfhFiiTIcAiK2rlv
kuz3/BKw5/cwg7gFx6gHNhvT8yU3Vtw0g9rs1i6FlagwyZAht021cNLesgJvQjMljyJyC15QcOiL
yVTIsPjh2+B+B0tCxypWU5KidiYTPcjonFbjSbn1OFyfRcQQylLDokbmGSeDz0JXSJ0ZqITV3eBH
UkjDs2Cn/dGP6IfQ84j+cnKXqq17EIcoou9jgdAojL0UHveuootY8I+Y6ACcf5Fw4zidTn+iUdkd
8PPddMh5zq8B4ulQnOmtSgQ2v+AE+jKWrzEdGG66NN+2dKaz+JlqOWmCN1p+e8JA1/3NbP1CT914
xOywnIWm6GeWGan0VbSEpPxqS2b2OsWKrABCHIRg9oxrcrlRaLm1eGzCwdY4bjPUM9ntiz8QvQOG
KngA6juNTj8O8aeb/faxprvwiZVgToG78aE1pTyX7E9/hpvBfEwn8wSeGjXwO2x4TwJ11hykA+nW
getunohh/dnICKFbdiuZvU5WoHZxmZzp4LgDw7TOhiQqn+xJOxqRo3WXXnzZJREe7PuKpD+DfPvv
iNpeuipen2JBGqVecpcp8Ck232W97aZkh/3PylnGrPnDbBaEaano/lv9lZ9W61XSIaJuM/WNyTN0
e4ycookPWzQCt8sUz+GHu+FYby6rAStqJ71E5E4+27GNi4ErH+I2ge8WrtRZ9pDSi+EcOkrc67N8
3CwXNMVlhTSEgm15UkqvCXOnWU8t7wCEPC3YWXLJCecXmMb3OLoRfq8Ie4jpc/NrAyJMEu7Z5I/1
8hDZpsLCPJvGnKg+fSPsCAyqpzxmQ3NNSpCGO1VPTRsPOsVNbMuKN+FlXVw2Ym6dVpEdY6H9Sxeb
NOr92Gb54PoFw8rUoDMI2sZPyHMJhAz4wKhXvc4FdY++uKvvf2gHo8plXI83sGDgLVTAQ1i5ljjV
DI4mc/1otCpm0Vi8mC5P9TuZSxNT87bU1ddKtHfQK2+5+Sl0aF9aIA6pDnOUYfJ6P7knkRNM2zBk
el0WJRl3rfizrl+bbd7bteXsJDMV3nQql3lCqbu2MOjb9j90hLK8kb4qjqVUhu1apKPfIYefVtCg
u8mk4+pQytG87PZb9oTzVvnOogrCbGvnt5zhWTngsDERIwmPnXyivWyRUk2tfY59oUZ8BFE9+dDs
YLxaCZQUWlqbLk6wC/H3CmDmYM7x77EKWo7QXR9K+MlCQSnZABBOdCRHFiDeZkY+BmUAJxclbq0r
YCxIy6F9y1X0Mx+H6lRuiIkJ6ePsm2pkkuZnlC29+vK0At0qjFHMHII+HB3wSNqLb50KFNpV6Bat
D0MEyHdMn0gvYmaAbyZI/FSRWAUAo3WeGMLvI5WRjsw8bumSc3CNOzwJw2/vm3xVHjqCXHOCF1B1
IWyFfIltLSPGdPQqrnMcrzTMXKDzDL3Ed/5//sJcB+g1U3hiGEp/LDHM+2S8HgfIQGkBWG6o0D8J
HCkSvPbqDT2LuszyIZTZHd6VffBVI4SXMYtzoUVKyHknSegZ6aa68RH/ZslHJYWE/S4MKvu01Xlh
YL6BfvEszkOeRDwRGBnGMgUVv/21+JcAW9HbYM4r2WBtONccwycNlFLAIA4hTcDQdELuDYaKtXrg
sZy9PCqUBrczqxdGM62LBsvmNceUlQ9RbP38ZcysppcHaknD7eiHjaCvSc/Dp4f2aCSniIdBOYr8
WZ+nZuvWIUtCm6WFndXBJlUc9xnwTfB3OykmRTPLoO2NxU2Clmjs+pRDRfbGmD3xuR7TFWwB4OSn
oakllNFwiFhL/sQYjXqyIuHvLcXuuleDmXs/nF4D8by2Njuc98YdU59gXCf6zAXZdeyjHAaL41Dq
6xnR05qikl1Rcr5THhJAH5VEeLkq0j1zIApg1LR+qP1iZ7CYL7hJkZXfVFAQJJD9ECxi052e1pkq
5lwNqqHoGVuwDbywYLDvk+f4OIFbAoKL95KBl7/MAS18g5pcVubJHTPMSTYiKi5qaqFzVq4ROw8Y
vGOciZEyVD+l8QSOe3lYMNJ/mFkA8+zVeO5RBShSD6P1Ga0IWcr9f7AI/SzD3IyrO0kSmmIQq9Uu
ejWMSlzlxc2KbFVvspF7DxmMxK5r6VadNC475uFwIzQjXDho5x88+hTXa30VBRNQzMhzY+WJKpD3
5kWcI2fdeXrC1LpgRPdyY87ZD9c1NOiviMtn4rmK4K+VtcFChz28Wnwq2vsdkj8Tx6cDBpMplrti
WBZpHWDkCX6fch2zXS4dKS5UKK9vLyAONqvKGUTd4GWOMwW1bdyy0XQ8+v9LR5Dgm26NGQVzzM3E
6d8OTvAfgAwExed7/mOczy++oDv0fDt7GPR5PpkbivE3Br1VPdgCQtSb6J2mjA/4+Z429lCLnzEP
FrPlp06nD/VtGpRWtAg+7BUJUdqxorWr1+H2Wz0XQLoFqQUvudMVSw4dfOfz+ou+Ibh+swD347ZF
CndNKFFwXXWsgXJaNT3qCkpUMGMbk3a9hCQT6s9WSo/VzL/wWwBS46qHrSHU0tCybmkKf6+xsUaU
wHs1Xtdbr4Ff9Qc5hNNWKSpZUtGo/thdCHYWCXBnaxYz++CKuGRppfIe6ACvgE7bjaC3EXB0pPkl
oZqRS/gz1DEnuynDYe+PqdgCfpBT94cvJwh7ZLE14o0oWr06XlnR+NRzN3NHHiCo+ffhgLWt8VuW
vrAGC5WtIiKfZivlP0+6HzkxpbpnLpZl8+r9V+poOVgzmx8msoWp9IOOXAOgDQK0ufHrGpAOnWvs
fCr8j1Ut0eBKvO5oygmzUn5BIQm7y9p7N4rv2790Bwh53GdM4+v4+cCdzIpHqhOcWiqerU0QYBtE
iDYZd8j5vdkcF9dJoY7y0wUZ4J28yu9TxWqajMBpf8qj+tj/EWIXq0jx9n4Vjh5AzyPKz6MKcBwk
zRfP7t1+qtLpRvSIgMoncCDSDHTDYJnimdPsLlLhk6bHnFJzqCmmx3AH9AYOh8NXonLNNl4/2uYu
efUNthVaHK/bpWmvLHUs5qtcOz+p5AdDBI0ekh6/qYEMsM94R2fN/2EkX9Zk0719opSZhJeCVfhR
EvfTMsdAqyY/+DMZWwvklohJ5kDBpUZ/KBSl08CuZ2Q00NGdslkhDst7ef7B6Z2gT3/H5qV2Du9f
F20Z1DYie9+URT5pxW+llbeOgRge1HLRb6f6NSiMcQkmGqu9IWHzQZwOm6Gho2zs5zJqWqbY3z2n
Eo7+IICoTEzrSYAzLVtdyHme5JG3u5PxSV+Vm9aGNBWIX0jZdtYxD5wRCTPnZJGHuXN4w/vjpuZF
B4OQpgyTvS/d9OHOp3f0OKf6QjP95B5RZmi7QRruNY46DtQjEghbA91yvUGpwJEl4+xkIneJiv4m
SU3oUqzjSUQvvhQ/kZS4YaRUDqIg+gwxXzdXnmR4/TNsV0PSIuCRgGSHGNzWGo/xxWv72c7nykmn
xFw3fI/XfOK/LDPDjVkcEbEmvbSkg46LRQq+IU9z4KLi3HI79HbYFCnVnc2DLkWUJKLmZY7Szksd
0sOPdJRT/XgJVzyAMH+ZStKcDhv6ho1dTEOc6o5CCDYxHA8NHlpbNDTSk4fGHIQ+fBN3xKI0kVDD
ap9aML2cEaK2FoCOobCgSjOo8gnQj7D/CsjtdVRWWKEHPuyt7XH2g6pLhXLP66mQ8gpX5VgGmrAR
7Pb8kmHNRTOLTUND36oPOpUmyzzVEWpcpfbqpUBhbqX/bupEoQ0t4CkRe4kzMpwPf9bAkqJ558uO
uzQAMmxEDQiCZ3z3xTTOkLoF+trrF83uxph93AVGJvxOtSRB9OnEQtozQRp3E+qnR14v7cj3gyfE
FuV2sXrvLON+TovPE7Epx/Sd+jPoqWdeVAwZsBB74KGGXX8Ifl66HC0cM3Jlh/CK4AH8IaXu8fnk
SWd4AGZR9eLxN7C0XNqAP7hLLV1zxE9l6/A2I6/usxVzQCAjYw/cHZHRDNYlcsQ0T8yBMEOO1A0u
EPfP5DzEVY4ENEGcw3UsVuuw08xjlQnzqYsYUGzDGkYDOmu4iiDwMtTt8giXA0YanxRZTsyX87gw
uDsQ5pfpVxxPsLBCIhLnuejenJ6VvG+fmNg7R2xVhgqT4hu1E+XWzH0V5oaacmVQXykhaBkhIWKQ
n9JZi90Rktz4x+n0FdjlP9u4djNz3Nxq/nuQZDFFv9al3YBgheeqnSDYNMWlg6Zr44q6xvc+4Q2o
oZx7ynQshxO2as1j/4golOYi6WWAa8/Wt1i6+FCvVxQZ4weqhluHUSefh+834MRO5GPnyrfhz5SX
eOlXwdt3JPLBvNH2vTfRB9U34keKtzdvi/ntsV7BrjuboslEQdaQao3z1jFpJcAcssy7IEsFvU+7
f3oMy+Ot32+WZBBgH6Fg3GCim4S854eeEvpWG5UVaoDDuYid7qR1fz+rGUqWVQEElbDBRrobP99C
b4vPTIL1cj6S/fZUgybu/SkF/Dpt+hiojZUtL0K/cE+f6ZsZzW5rlDI6J3tkcTpDyuACzxmiPQtT
LeD0ypjrtQtxzlYoENzz7GLso7ET2ojmM+sy/TNdwQlTHWmufS1WD0sDO4E29wVNCCqHOXCEXh+O
ljistxDWfHw7DYpt2oMt80cCF68df0CMQsmcvg93NKrchwtny/ZGqGjXeZcfRhcVCSys+gbox++2
MbErsLuywSjKFrgkjUOiHKTVhuj+HPwzMqqUvORwTOIe6gdD0N/gY5c7oTkXOOJ5KAZfGe+phOof
cvGXZWO4ImO8fumPL12FcwMFUpt0jqi3+OY8L/wX4P62Fj7uudH0igwr8cJYt1Qc4c9H7WPGfnob
l8i3iPxlFJSJKplei+u/cjFG5oocmYRvN41qnSquUSsveFWWf89Z10TiwJtiyClWLwG4DIiwjDf0
9XNHOO6GxItuS3nlJ7nhI9xhhSK87lzNl8g7fsZz8d+WVUYqnI+HzmGuJT0phqgyw1nhNqYqiY8r
CiyfS0IsKW8Hi3RQ04L/ahIK5PYilRO/y6ks+1Rfbgmm8++CisN6I1GE1eGudOJ2qP21LGqYC2Mq
YWgMHhVU+OIsuT/0WcFYU0dyiKktTu0ywV18u0aw8EVQdcIILREjHscDEl7ZbApeFnhB1o/UDsZp
XVRg8TGnLAP2PggLiegScQk0dgDlaSGIAUegKN6DikKwScl+kS0r8zxCWF5tiSsfECJg/g7nrzs0
wy1ODu/pJ2kWuU/6WUcssJL9x4M4fj2ndFrB561yxIlijBTDeVlZ8SgtNjEo3jEH79wrH22JpmRJ
oiwWr4VIoSrSirB20OksPQP/9//95s7BCSr84WhHUx1GbAPZtYztzcsQPS9CDMRtM+92C777xQPG
d+91d4nWX9oc2mbUJT9Tw+G4aYSSUk4mAoJbdz9Ujjex6OrwyePtg3T06wWJva9mzo8OZtljgnG+
kxxfzSuwgRESecFDUpVngPb9ktH17mPRHQTkDR1O3/zDeHmbID1lGTWy6UfMPdz9ZnOhB/rHu1CO
FG8vRQqCCWx9D4MFWZzDFjoOWpxhcl58toncUs73G49bAkYPf7Q+jV22khHIZRqVMGjC0A4Gz5Ro
7H0MoIKiSdYa+tiUTwTwOXwzmA9rhN6gvncrJJuc6VSt7DkQ6DB0D/WGegVTNZlychtFr7BfoOZ7
8aZRVxGM0Qy4hLBTF9uOjotear4sbKAoKaLWOBeGl/2HEbsWgNikNUo8V/vlZyQ8DtkXRBA6on6E
QFRHqLvGna8e4RCcsSe9iiU20y0N4358W5lcMBm11rQnX/IpOdvDmDHh7mSHEN+07I3QCmurZrwh
TJOljADcPke+o/CeUWUlQg6coEx2SEFgktkoc9igBCDbT9JHSG/FoTidtiRnLNOhJ6pcCLJk+a3I
GoTXxYMLF7CfYS/nOC31Pfhdgj3+O8SdsD7UounLOdyvq8X2WNbYC0ZKsgRLsl+IDd1xKmVIsxzE
PK+gpPuCo4a04a5BFy+HkyN4olJeeUHWUrQe+IMAq4s6kUODEsLSN6Cl3PPLWh13xhxKvkEdaqcm
fPnNyssAHk3G5wzXTsC9KKB3QLRgvKQBlXv2QHWnRxV7pB9KOOXnE2/3S9u2Epph1FoHDwQzzM4f
dGqMNSNogfa/6bT6c6zMBPoXXlLI8JZOpl7+RbGrQAwIP3seanWRf7mEiJFj3h7zkbDJgrdlqLwq
UAv+YUjseF5jGvL2LXfFFVHeWryvAj15BAlSM9ctjU0tcCNKlVZl4L8n9BlgIY4WGMjBl8BDGrFI
EIiGrm6bI5ML/pqyF6XQPa7spPN2hjjzHAOoFToRL8R/kB5yT4U/me5wAPAYLfoydD/ZVRiAEXmb
xR7+d9hdIfkoClOt8g0ODYGeX+y1HqoBgfgUmH0/W3NmPw9EeWiFYEA/D7kGhl+r2JI3lXWwBc+J
IDdREVzbwzBI/JVzPi6JnS2fjM3RGefe9KNzXQXhoiGBfFJpazSI1nnwCWM7ifySzXir3AjEI2Hc
YczoR1AQ5j3NQxbEm57TTgwnGoKJ3Vk4hUvo6i+aPuYrEQlSe4vX/RT/xkvFYXBHBzXq7MuhUkX5
qeV0q8efwNGv/2rk/vK+XQA2mxAYCKstwPphBZGT96/+xtPDVZfTvj3G7R96dI81OMw3IrpRH8Km
o1QQZtvIedXBkcWBOkd28BAC9Pd1YRcZGwtb24tbwVvtm2WPPV77OA67a0JEXVqrBsRTPvjoBBkU
pTlH1QIfN5YGYQSZbX6jXif7L9vI8IB3xeo+EpFB3Jhd+JQpKGLTYOSPxsxSS4+2Uo6/uOBPxwrt
YBvGa5UOwQYLTT3fBTWZAPdL0ETzSJVqrc9swRGlBUWPWX0PqhEyCZj4+1hYy74RscioageiTVWc
JX4LjQZlKEPlRHDDdzrS3fE0mcJ2ho59ln/1ds5UMEJoYKmlL5K2mXzDdDq5852mJEIK+YHJyFcT
lOtQziMXbSSa13NoBMrLFud/19/UBOK0BWpDK+6v4GUr+oDAN4hxWxZCrvtMJw+eW6UIon47UvPj
H8/3HvAKhUnpHSz6WI6Ae9rUYOLq0EHpQrbeL8MQHYJCg9ToKjLFLKZ68Z0C9CfCS89ckp3IoLvR
fK1ruY7ltbC0xvJUV9+jueUSpVqmOhuK6wpcAheWYe3qF4zV8kaNJNQ8b3z+jf4QybGuKy4URAv4
OArMD8dBkZmzZkGs8yTKodkSrLRSi+gk95B13GxpRLS7yXcgBI38RoxoCJ6IlVQp3TfXjzAVyLtM
gEKX/xdmkzbOOH7VZIHLTKxkX3QqDE+hpPwd7l5HYDseoMKG7Ux28JVcXh5qqNzm4V571GhmPRns
QFQGzKuQFtnizJxZVBTJcoUnSedtT2wrgEqvtaG+arL8WPyiiiVrViAKDXzrdHd+QwrWPJgm93dx
aULUlx/exzaFsNh7jXSwU4CAcm8uUwhxleowFu3Ns+oUOLABprlL2SIyeBvBWeE6gRS1+fi/Zk4l
o9zU0Ebwf9MpKM0A0kYze4rQNpmv86/iY/Aa2l1EVR6L1PhMUn0gJ6gqji5E5QyQZy434ryd8Dat
7dcu3jzG6veVc9WGCL8vIHHivz1YR87/9kDBtjB5vGkaDrwN5TRVM6nsetlC1d6BhIth14EeYS5r
Z8o05CBI624bzW9DHjIodirEKEcvV8eATpQ612CNS4o3M6AL1EiO4NWVF3F5k+/npo/qHHixEHfj
mbZD7+OTbuwVzWVp1UIuj3P8Bg0ilcmEsfWzkyVtnsOoPrV5SOMShXrflG0JIU7jlVJFTDWQZeIR
0Ft2Pl81O2VXsDRDlSX8RFqKSNDQkzRV65I3dkngN39bwMUXUBcn4PuMwLLcLbVWwUHm/4IpbHf7
EpVVliD9CPXI889Ogi5iPSPlO8sXNHAluTwgpLxW76tPCH96z4OLuETyL50Xz/JCRD2w1RKhQ7T3
b78KYACZLvLTzBM7P3AOSnFoBJZsjhZvP3pBjVGEErAKGM2pb0Yo9rTx+jDR5AsCiF9A6HCqt+FK
XhlEH9VIPlS+1SL7aQjtrevjCCkj+28oQ5tQt0Pp01V+dVykdnI/W//fIFmRdgMaVonsB606ZcQQ
urUgJucceODBkHYoH+NGIvP30mW4g/SzYoed+slDNhyMXdTcpRYaQTYeRyaSntiP6IKzI6z87x4P
4QCBGiPQfo28DeJtt+P/UzGOK7LFm3vEvxCx8YDP9eaH4P7142w0Za/5tfE2kAYnJ3zqhoEmJ+an
9sv19UkPjYFWj8TNM2hDJ6JIX2kzIfCghjWyrEySOnhJW4s0g+MqyIinGsethbuQ8/i+FZQPSnP4
xfF0v3BZ23cR1i/jPoZDG0J3Mh8wTrncGtAcm2M4zgXwf7lR01QEtz6UqEoUv3fM7WwMw9nowd8c
o/0TDn7Sl75vWVo7k4pKKMmHtRWS8APIckFimCbGSzJhNgN/3ZjQsvEP9/n/jaK4Y0vlEOeZ7dH2
FJ7VSYUn+ZYpnSAT26+DZl59OOw73NHjRcxQhNLsz0Q9qJTix1cpY5phIcXuIRFbMSU+JRloycXm
AhGAttFKBTQP/IwQzzpIPTA3I59QAlg1ODJn+mLiTaeUupdFIzQg65eF02Mo8gpdcy6NveG+6fhz
NyGH9eESRBzBVNDTOIGv2z/Qz3XYktjgsux0cx+/lVwMaT8Pa09Sjqrd3Rs2+Y19AmeixzkUoPmx
8XiYJUASmmI2Wq0oZQEBo74Od2ZqFMebV+rXaq7gjwomZh3DIPDQoDIw1EDcV4bUbdVCl/D2vTAK
RF+saFBLfztKkKhYyDYJyQIF+bohAfUHB9AHUbM8ay+GmkbGJUIMhcHG2KLZPWFNl9J64U6j/Hrl
jv/YWQqfZgQgCxH0IXiwr6OWpjc1ucTK8RPAUpjaGIHBwdIbEMmGNMtxRnpABg34CKjL6qOL6f8w
xpVsdny1SNtJ98RskwMgBjNnGyQ17UWR7i6BOP57tK9fj2quhsJWgOuWJBTMBmu3Vhp/ITCfxrms
aA+J5IUrAsjriBJnmCdr37r29+2NfNPD6Kw7LrZQJEX8w6wrTAI6k+MXNs5dk7VRqHqfKrcSTTo+
vh+bSXpFlqyHsvrFOnc38u4+FS4T9xC6imbsWtnd5F1Eu2YxgzwKu8dz7kSdMT/+orIZ+vlBcY0J
w3bw2B/ar4zZC9hihij6JkhD8piD6bwaihRCqJKuJ4CDixUOz32HNCz6gPygB1v2V6uYUgdp/TNG
8ChWqiYjPBmvYfGU+sRvvJY4+8xzOKrCnYVtQG2Sqayv9noiByHZ2coLoM9R54SKiUqlsmZiQgmD
+ialek1/14BAlRjgujqGXKubYFSkBRZ5B0D/PqZ/Qzi6YNXPD9jtC2ji/4FHszAA0V6SdqIMm9yW
uUsBVeqQ6tqBfZaYGb6f0yVGufvL88qazE0pQzaviVhvjua3GREUtd+p0iLlzVzIEK56QXEhVShk
9HR1NY/fC5JzwSTyvfAO1TuQMgJmCNfQTUR/9SWl3A3aijhr93oLk/zw69H2gG/CH6XFwWKWvRKK
uzouWlnwlX5qVM3md5h4Rm/HSoPzTfpEtaVm9/41j1RhBzWgIKotHTqPb6/8sUKeX+aQOxsxo+1l
MYYozZ3oS4O+ZOLdCJLmPsGyWgFskzLFtqgRmmjqjEXl1rlRvQrzjLogAbTkFuFBrKRwZhYl8Wx4
uw+5ctnId/3/zkBLfkySama6M4+68t1vsPGqio18JGTBGmWbQGI+NVKTIMB1KYa0cLpI50VDxkWu
k8Y9htdHSFImd2xIH0HGaMHjW9+ycMyq9xyk9p8ZEOTzNfgHsJjTFxTIxXrqJjUc8WfoDoHqqHDd
mpH+8qlfl8aqjjg9HNfvWlJY1mdPMZ7CfTYS7UaByh0abbMP6mUP2ibzb5U8a2wkpUwZVWDMyJep
AU7/iRNUOPLXkaW+qmwt7P8CQXadZ0Ovsygj6T4mAeS9w+Q3LJPS8NPNe7cHv1C43FPSyC318Vsg
LtMJUKOplD8C6s4mHCpuDVV2GOKfVe25Zgve4AWGPbF7DNeR55+CHRxgYo2HXPTyTs7SN/zq2G7n
Q/fk/9edgaBWLRcNKgAT5TFP4FQWbeFUpQFo7pdXbuusBV/2hTiLDdQ7lw2FM2CdG1G9mnBC3UkW
w9HYPtxuXf4cuBcEArolduBM3FGSTH1p7l43W8UsdmlZf4IlNrQqT6677gunsDn8G4EDNnvVXLd6
lRpNH7XZ2RuRG/xb5qr/zvxGwGJ94UitrUV+xjJJI4KjGJ2P3NyOCOG9+EdyNbTvTdWju618qotS
4KJf1O4X95n6oKQffRvTpaEH+KdCZmRx7LTc7aH2MOiJHNi6cwS9A/qL6CeXKaBq+jzEnyeHSJeH
flV9+p8+Io8olyHXncZrA6S8Ztn70lI6+8It0ngUtV75Qe4IYU1f+GUSDDOsYxgQkFB725FO2bLS
xUfUgI2d/50LYZESWVc6/PxV1nixW++6ziexlPvzjfXbYZGJmqmI/CTjGnALO/uoKPhI2MLjkDUQ
IH1SJiykq0/b2yosxna3mb14P5rRtTvcQd/XUBXN45OwowTZ/6qQnKvtOmyKyEOwQXOq3ayyWKwW
FBzMTDfxWFSAQb8phUPUHYQ/GCAPb1AsLjU4SXqOjpQvcCLa8ckhajnA4K8FOx4UuGyirgKAS3fG
wQ0frVFvlFXuDJKF38obL8706MBellyKs+oQy9Ei+CM9RcFEiA6CsFqou/v/BXJFF0oXSeIMQ97c
l32cfodMkTlj6TZ//xnpD8PgzPNpwnabo7/wpa0II4qU7m2w2bWSnNCse4r0Pzu0kZBX55rhEJXD
025FjAfa8JYOCXj+AV6XfVeGMVCWaC2s2ccQT1MQPsXNzSPbpH910oxfKwjbeBRHotNaubGa7qPw
J23qrMdtpQhkiuWGoDr0slXNnLejtNLslHyHMCui/1N3rg9yxvgH4ndxshksmV84cmWG4YqXC0Fm
ro+zSNo02WAoJPKCQKWTY1iVm/RZwbuvEbg7vELARSTsqRrAv5rhmI6+STEXfF6KV3jMMTdzZcqm
Fuald9dbgAWsczQodSNhTy/OTiOLS72TlY/LOU0qqSr1BBf1jnQBL9bIlqSu5S3c4FrUf2ozYY7h
19w4baIiQoCTEbeD6+amP7Gu80pbm7vapql2llfe5S+GcpmjircGflggXgtHkXXg2BcHBy+pMT1U
M74s4+Y9wL0D05Ft0aIZXLPMbcFWY9Bhk8W4XCTqV14mJazteznXd03VA1uhcLXBzT3Gh+BnfQeW
BFgy6s8ycUkbTyjVdAlijuxEyrbbFUqFtDiDbKBC4q6eAQq1m0uUUcxX4vlUdBNs/kOvGbv8gZjO
4EM69I7jHgwFrnZ+qSFO3wsHmn6LXssC4B0/bSHPDFai7+m+sAWB9o3Zfrteh1pR0B7yPp+oefp7
3NqEITObE03Ev1LHlvjX1udPXYDbz5os4XuDIIFlWllDNdO91MNr2EJDhqTZDxe6+Y44+8m6TQTW
7j6MYCpXCSN2gSlaWU8GL9ByLZDsKsKVpKs99UD/9mYU2AkMeDpLM74OmR4bV/Dy1qZ01U5zoMaw
PLCayHH54+N5YQYC6QZvyJh1Cxq4dokSDgbjRQziiBlU6GrEd963fStIFvqdecrjWpSYuncrit85
roczTNUmDIcy0TaA/n6mYlnWkJndM1ZAgMNprnpkt5D9w299Um2uefejNJPqjz82lwftr/UckMsd
0GH/1foA9qRUzfpSJdL4c9yX65prehjW4lek3nkHZtuFKDCv7HB0yI76UVMP46R996eKuV6eFaaG
rqZO3HTAw6G0V7hdIhfkm978VBYitdIJkEzCNpQfvaOLWG8w5EaPA/UGPkYw7mgnN7bqGrI5Ckv9
Iac5FE56uLkDdw52BDk8e1ujaBahZDfHqUmJgatwThqwfKny+UeNA7Y01YVhDGOXGBkstDbEQbED
HnphmMzYxqBMt9+4D3FP26LLoGUr/r4PI0fBugIMkul31Zpnjny5vNVYnVIGrXskOSHAtXQ5ZIbw
F0qLr1aQ2kXerfNtoLm8cbhqa44ENY0vR4k0EjE487PqiKY1BTP3dqtgWQyqwgzBwvgMljXWwOC4
pobY73gPgyCPZ+MFaCBBDxebTS1KPsCtXXbWtHn+HPZF7JgKyp+CFeCGS42UgZJ9OtB9AxCOZdcI
tvB5NTNeNPYaEh2zqf+I3AD2QhKnqKzCH7wnXnKWYdkXVRpMlIIVqcG2VQ3/koY9nnv3ZGGI5EHH
a/I7l/TXr5G36vfjdRNBlIt21F9fEBl/YfA6HZR6WE5xjF4mEqNhF+FsHBo7vuXivkBIhOqsTsNC
q71CdMCmnsskGHfq+hQwP3aKaQbUd8pJIrJNVGHl1PvyzMvuaXELcQgTPV7S62gVVDFj8L6o28Gk
7JYPqxhmAoHZkf8kenZkv7FSkzSrrY11CU0CgCSQ797NqYK6qPexUWutmhmMUOxbti2xRymLEIR7
c2QEs2iDUVAGm+71K8V/AEXLUAoqz/zfnZUi3JmwVIVBbvM7x0CtrUBiRq1/c6AVu3dPMu0T2DEW
fJAfmAn3rtKPQKW7So4ljfLMImowI2ZPoqR1z1lhyQ1HEHjR0vusVwyxluvQ0CyQgnw8xJjTYcrW
gQq0+eXsX6EdxCGz3pr8NZLZzwWj9XaAFrHFEC8T6JOwArjLLmb34/V7zFfH2/5rePb8NaIyqBla
mZYQNGIIFoLMbe2c0p+S7QbrTVBB1gW/gUVoj6XfNGWQ9oNAU0Y3/9orQTMoOcGKjZCTJPCXFy9p
hBc2ozNqvxY48n4rSZ8ZpE3X7DDGkvqzEcp1MBdoUntodmffBl/EHHxXcOQxnPZRSUsGIHcoC14T
9GI6d4ZSQEX1BKUxEaIjUUaKcgdrZyexHSy/tOhV7es675ReQzh7A5KQrRQPPBeou7xBbunCzwyb
7K6H7aK/CCdaP4TU1qIJSZ7Q8+BERSxqMRDBo3YAIXEyrf8LjF+0LTBGU/B/x/pldO1cP/xuHqoE
oSSICgiO3OkYkFrbaG9xmwiz7/CXYJxLmxgxFVSiAyMdYKa+/P5FLX3eFy+SaKVUcO6VqD8eGx+Q
xgahTBJbutk4aZdv3VGirLTup1ENC+WEkfb6mFWCj7l+Lk4m3sby5wqf7Qr/3ZQZIYZdVbVeUu2l
ihQPTMcaMIJlmc+nbQj+cUF4OAaEQUYD3ppF9329tBmJIdR24Skea5a8u9oDMRvbSd+7G7coN++s
TqfGvo5O6vmt84BsjroBFJf8V1peuKvSFOy4W3GIh44drRZKIv1VK9DZWTFSZ3klqjr7V22t+p68
YOPj3oE49Qyfe1KipEj+59H1tIR/O/CIVxA4fhO75oCY5WbkroWM2i7jEtJ1c9TuFRgk/mkti0oI
0Pok8lAT/pR7nYmem+rKbPYEPlz4L3XEYeOQNG3sdiA+6AqD0uxWl6nDTaF3H+XgEUeHDTW+NiPu
XNsOHGI/UFvIh2fLbbZpsS515hmTwLm/xj38NDxGLHX8IASz9WuvE638u+mDnKJCtvLqX2KcdKWt
5wVktBFWlNMQmB0B8IC/VgiILqBv2miuYFDzSnV4uR4gyfI2njGcUw5Ip1vKouQ3ZMTv3yAaatrP
aOai3NNTtba7zrZwZoFFY0whzXHruUhf7j22owVXdrjygwC7NK8Hi+X99LCbFUFyvksQ8/X8ceMW
obIjG9SkVV4FPvFSbR+3WYjo4B0Fwsjo2GhrNDbCAIgDsQJEboW8IoeQhCZHIdgk6ePxN8DpIhoZ
ovpHVl8/lrzlHIbkRZWCDD8iSyk8im7/ArvG3K2clS58LIykupRs05J8Bvoykomjj+9M2FPnIvjc
rRcx9oBcrxNMac5JlnjIj2CB5cDeEwEwbSM9lHPOxo1oJBIutwpWK9ep33ls1TZzbNn7hQZK9X2U
t7aMP7pCM8HbnMKiI7WR6P7nFs3MCkHPQ3WZV768qvcO4LroCOFts40RM3zvb50QbLINr/Ta7I2k
vwzzOE7qFqg7Di0chBL6pocDUoTjJ2UMnb62yHLJL16A7YP6Pu9pdkNYCZF08vs15k/Fxa1GzV1I
5o7kajcgR+DTP9huYNsNfbbZp2CBT+H3b12UtNlZiLceunGn5K0du/dWhozSVp+DDxWeLM9YYnNr
mFs5qgXzdwtcgYzc6YjhuSySsbpVDBHRF6CrD/VVJuAGkp4rRuNlFLe2XFZJTw29LnKZdud5WJ9m
V8V6o8En/porXv1iMUtvowu6BW9zLc4OEj3aC4u/P+8McNTUJdpWjZ9rUfJm67yZyGNqEt3qUhne
t2e+Ku4XwAeujA/8q/GS96XL8YmglqZuvN8Vw/v6JFI01YHtxkWuBHtHSo1dYEBIlTktIu3QOeIX
N9ci/Xic18WkIKukVNvyXGkJrWbvPJAK4hr7gZGcFowGw8+cpJNGDDWsuSMQkgYz6RGe5UsR8qpT
uCr8Wt8ohVO18hnWHe1Yxs9/w82WB+I2ey2IfTTvEQI1d3XrhvMrKGBK6TVz4nIxZP1jq5lCoroq
JWIw0du2Lilk0OzShZ37TRCnCpF71iQ6wbuibDpju5EgmtdiPUqp821OOSdefMoXLbz+yWqdVUvN
I2FKFHbIMCbldoF4aglB2Ha9SKRKpSyU5YUhwVzFhGZ4HGyrCctgkYP7xKo3k0YICWVxUnCN2CnY
XcIhUdxbb0f4to5n7lfJJpPMRSYYShCqYIrN2mGorCisDIQN/S3ofg8ZQYKeel+XKqVHRq+YhA2h
m0YBc+iMbK8feEzNc8AxLq6mKUdOrHIybEiaBs5+ekG8scTdgHIIWUU2ScKff7JWAfnEgb8AlSjt
SQ/LVvt5bOuBtL8bl+cKHy4KWvFioLboxQ/E2sgSto+BeUFNOSMW2/iv4y8uSpZwkkmaXeUCdyRr
1SoQXj9ZLltchUsnohbxOMBMpzQ1VnR5ChHlcJ113zEQv66tHheCMhEL/sJmki2aWfkfDE4tYwf3
/KguZjAm4s632yzqH1Dj5+GdSLIEa/1ZzxlwQsZjp/ufq+ADk0IWQOacsEW50EZ3ep+dLhRWGVZR
TC9KOnpkWO/TNYgS5xXe2w3obFZo/oMtb4PLPDTC2BzLpR3UPGYWobnE8bYBJMJHYZR2CYs9RBGS
57cBteOTZNKiKUNNmwNNXwongJW9p3osdtzQBFYeU2Go8jS6I7PaKBrdmJI4UQlIDIvqq2iBH2SF
a2a2TyXLDJyriJsGW2AyiLhjV0ErkK3CrNkFL836LL/3Iup5f9eMIdBdbwFi7ho3Dv1PcmJcmuLF
qPE4B/5C8EUuZi66lu2Ug8ppgbARl/NU+05uhlvbO+2qGhDk/dkGXMjnihUfZ0T4C73rkQOyMWnD
n8rRRlc+24IjOU76CjwnvMwp7lSr7BqEljqBzWU4o44ehVU8tWIbDxWdf5FNsQOhMzR4A+FKCbDw
9KtW47j6WrX9u+6RBrafz7+IGV0AiluyvnLbJI0/pKwK9Q4zpxypET3u4z1Ep/xOod30KKl4L7cc
vGIdQMYvmYRR2m2E8/rLnn8G5uDN/ic4VhkSbfM1r5OO+QFkQX85+VnBT65jhF5C2C09cP16+0AZ
M504tDkYZUdpJJHLzjDE/v6XFnkxzjTPwGN2py7bHNORs7A0HfUuDAwPuXy37DHCg5/+5H0MX+MB
H0R6zcRNJjgDemDWrlsWh2HKeDcDQsx6EdAjRiVhV/Lx49fHC4IBBJYSChxT6S8/FVANxc80Hxsf
/3BGnw9jiSWxPBopqgwa7DbJRBceY5ptsaNVKHvSECc/8KSyAF7q4qJegVWVYSs+NHMZZekmH7hG
gxhYcgERQytEKxcL4EO8xZ9qElYa5nKC8Kz3nvl2SNjLkvXDuZYLw43NwHt9Y1EhHKqLmAfxAu/Q
8j2cKAbgOJ2ZFESBxstT4jFFH9BopQ66FmWqiLnXpCveCDQlqu3g0k+mtzI02/yEdHbfyGf8wWfy
VDQDHZI4yZHVt19g2h4w5LjzJAUCagOEnXyYL+kBHQrFL4FDwLUTIPCJ+Zj5rdDeQ3Te8e22r+lk
k5IX2YhKeyKMdQH42wVeGAfrI2k6c0JmLn0dTwzxyeRvgRlwM5X32Y9hFnA6h0w/so4xCA0E6+Li
kQtV/GswLJ7jQPmJlt+3vqCLVTv6tgWbq/FSVjc7Od6/sKIvZDnjskZEeroLbmpxKaDj3r+ENEHe
k3yPTiJbd4mtrze+bzjkEriXhDY6q+mqz0PyHlFN+ezvVg1liZmxOgVchLuIF7CC/2F3OuKu9bop
GHCeNDc/sgtRayJb3+mX7xgRBQS/FYE2YN80D/NGeKG2AlQbEUj3uJblGU70QFer/9q1ORvcl/P1
+OURoQDzMIOIPXiJXTe0oiQZTvgcSQZ34QSf/EiYLroMMtC2ltY/Spz/Ec+oBPHuk+9+Vde2HoZs
sSDa9tdE4tLocTR8nJNRKMbF5cLqFh6RxKEc4Zbq/0Q7E3Ce+UpCb2pbKvo5IlqY3hYE9t6o9wxu
yRxRfxPIHsXb05NWKLruIs/DVzo+QZuabGd4RbDNehB384YfApFLVP5t4tSYBtdti/u1b2vWBput
U4a4rD2B6kUAZWC5iJjDbuvb5DtbVApFb1u5RIW89F1G+e7jAxPpKb1o9j9IgqZiaypUV6TkLlWN
dJKJTnz0cn8GgEf9jomd0mgOr/qv0YQfTY0J9zZA+napT62sxyY9ustOJ3VfWIMM7OvD99V6qkIw
0OVlpc7T4dzoBHXbZy7/nUx+IcKXew2kSFL3Ff7RPTAV5FALD2rfgbuO6wt714fYh89Fb3Q+DvXl
tE5JCcxYB8GXI43/LO0Lk+WjIrI0rza5yCDdefDYSJoOw1HOqm4b8urgp3AwVW4lQ/3yebYYAv2I
EPbYl2xQXoPKXpsFA8xDRP20kPscepRXjw1X6UZRkpUilbiIXhspy+GHwuMfVZiPVt+77dy0yFck
oRQsdPVYd3N2trx8cI2EJ1RMDo9Y000tF8o0lnCNDfJfSMR35qAndvCF9Vq28AdtLzXAUAA58k3l
Fq2nU1ykBvE7fCQR3i+AjVEjo6Nd49vnsanaRt7fRbnWyfF8k4Z11XrQtu19R42LbbaFW4YdGYLP
W8c4Z9D67d+9DwL6xwOJ8R4Xy6niGV6RPwc72iaPb4uMOlMceI4mX5W+YqZf5ZzxQqgzX8q/R2Xm
ACo3QAy5S9NMpu8y1XS6pOANnCXrdDtcrAbDajXjEVTbr5OdGHD91vzykjdJlGx07PFPYOzP6yGd
u80Di9sArzsEkRII/eWXlgTCYiqOkQm2FMj5IgS2Fzjbvwq8p7oE6HkruyAbyvJqY2jH9WhU52Z+
YCqkgv1PplWyw/o04/ZhDs1+YPhbEgt+IirtCuZiRV9VRA0aA3VDINmCf9KBLjKln1XLu4x8wNMY
N8HKofqMwCjbXx+ba4/J6RgBClgg2o09LAVf5W/nh2Zk0JbZ9xytAN9UndlSPKufAdcSUqG9i0Lb
FGFDV7SV3wrRCgMQwVjleOfRAkh4F9K7N2wbcvPA8/Z23tqMDDK23MvJfyF6y95ovvgzzGFmzJPJ
Lu+yDIgyPosgagAFn7AuQ5+mI7slPZF5FmHlTlJ0vNyy+0WdlB320rWP9LY2PlFHX+e0FZxI3VvC
TvYapXpTAPc0h9BRqnM8uCGonq4BE56VI1viWl/kdgeei23++4fTOKNPkUGKI4rPb+YOgXddoAUE
fFmypfw6TS4QKRC+UF7V0iS6zYo24Oz0SGU7pj3R4A5zO4xmlD7vjA8QLE6SGZ9ZqTOiXcUSpCnj
t0chm/El3jQ7X0F497nRMdbTmWCASssYI2WKhgDe8cBcuyK1qAeuy4OYuXMW4glWzrss3zqA0zvi
9VnbqWORF9cXzqCFsG/Za0O06eAPLXpsXC+jV8VsLbZP3v2AhuhM0VCuE2rcxdJ3g92ST6at9LNI
43EFRatY6KegVLfK9fEzglhGUQgoK2r1xSjLB04FWGnxxN9zWxan1NRsy2jHB3Xb3G//HaKxjJm8
swzJCNwpe08d5vJPNqzmS+s/xjx+DEQrT0loFHUCyPcGtX8KCtVg32bZHd8Kx+hMYwm4enn+Gkmg
RF4m2I5BCBkZMSDqowfzHjem1NAA/wbk5MyY6SdCBpzVvW5f++tzqK77VBPbrNesCjXpB183mGBL
LP5GsHhDZy0+2WUrP29fKHU9cMLHKkE1M50Dd2QXyleZhrB2vaVETKhU19DQUxaFq/543PvzO7me
/uzhi3+5WzZgYAf3vzVrfKvHe+M053wjF2PHfaqn0jsaAFMvHtFduoSCrGRnr1FoHz/Cn7daUnGl
tUURlB2ImMFpxz+w3EPN3bpQvKEE/kml4qlIxlGi8B7YJBr3B/P3IWnLyohBVNndOOtGZDrcFq7K
3gbmG+/8Q7/Bd/dCg4PcWLShLKR0MnbNOs0nMM/rO8jTFLUQPWEWiLfCGDoRFKUwhWAGCOaACrhe
NcAcHxEwAlAvnlUm1pKy3tDSA9SmPd1dcPj89ZOYHDtwpajQhreu3OFleKR2hQRfFlaXkYAxVA82
WwFG+ZdQy5CqTrcQt6mAovKY1/omeSjaZnQZUGwvH7lQTGD4Uw7pX6XXgT57w9hVK98DICOLYp+A
K1zY1BNSZp/VS14zUw2Nlc7QEP9lOTFealvwXgYKx4hvdvL91eIZ3IkOdf+KU4ZatiuaeANDrPPG
vKuLoxq7L0//gBZxD656X9hi/rBz1fUPCaz7Wx6CpxpGwDHgUKuELUAt3Qz1ysO+0gp7KHIh9TRx
XFzCQ7QzYAbOCmgz0GrhOHdK2wFivxpWPfb+jsY1Q03L6QP1oWocd94e9zmR1D4k18rbKGQGHFRb
NMRmJ/hWfCWVjtbypYXloAOjD/EU0MeDAHXU0V99612gPCppmFf+fbM7znF7qV8HLdLQm3i3RPci
SZyeu/kagt7RsDlPzOJZB27PXqX47FV3ZX1u90su5Ghl5EyGhIzX+LcVBeJoR4B4Xo74OAWJo3vG
pudbl2QSZNgt56YaxfghN2HYlxlvoIo2r9UG7zpDhxmB9bkqyIXU1OY9cuUdzMbHyEX39e7dpw7v
DiZ4/ViBiHgD8k1RS+LJ7bVO5DeFT8l9ofHSfEwri+zt3SZHTtqW6N05AXJfaFfTncDgveD+4IWN
uFiX/TGexyWh5PUYl3cSU0ZK5ZJ9qWQAuCL7sEHK2lFfyEMFqXr3HWpx6glRx8rNtkjGYpEU11S6
j6+INJtnV/J3GTRrh/Bf+nvkSDO3EMHDZAkb2EssFtAxIYbkhKPqbma2pfWlwjrvq0f5NSEGOzoU
kVJgOEzejkuBEWF0XYc7Vk+RvT1Wc9bNA3xOo6r78TgHFJ3TDM22DYYGQAN466OUYQsSeATdBdgi
RiwGBiXWk/1EMQcHczrrpoZe10yLIm9rpS32akABtD8Q3gq5CXm39qM7GoPGiMIPN7P5vXXHlwWv
UJgarD+ly9gvx9s2d8jJLbt5HUgwm9fSJhFlwCZfmEFuICOFi1qNiQD7J+Jv13lHHKQVBXs7cB1g
+g3cOrRGNEd1lR3IxLpLCVmbPCxHnUvEjyQ5J21eu+JmVkL56MBetKf++A+wxCtZOPNKilGuBa4+
CXJK+fnOx4pn2BuhdnPL1HIG3996/POcoOE4o5bUk5qubNwam38kMRrtFacSm0Ga3j7jmPeMKdSP
weHPMit7J8C0UxcDYDX+9J5HOZ8m76PYQmA0pKDJoHCWAH6VhPDMHP8U/tZMC0kh6/NDDsMbhFcZ
1NBA5KEKCJ182CAGau++LMKR5EGOQZyOVlWqvRtpAXcDDOXvLPWwhcYpT+JLhmPfnAoeZDnJTC4H
dkUugoKpfJnvGbWAjMt+ScBM8hpFe5x+hxuvyRtUsKktn8z9DqwCkW99mpKV0jIwAcW1GMQAQ5qR
eB3rL23tIvtJg+oMISTg6MicdlvigJTwsOPhUABXlKJwZK1dQ6ue9ROL6NdlhxSROROApdajaoym
rwhh3xfaSPgzffOumvNqOCd71ifY5DWmXbJD9yFY0TNqAT3CJd/7QBwBfFNbILpCl7wrJsRTTp0v
aVDZTSvMa8YbOTZ5JOXlmWlTXz1+Szjx7O4FtKS1U02rlM41PM5MXzTkxxoDDq+Q8lwIhgQ5xkRc
7QtiMif0J+brqRQL58XtZQ8jVgNrwVsW5/wekvR3zBzUKb2V5s6SC+sNa3Ymyvbx/g2OULVTwr6c
L/RKqxkOSyh+76robHBdOBstrZJDMILUApfBviJIEfpTv65Q7c+LZVca1u+qdc8L+AxbcwouFoSj
NO0OajL+zGYKaGmBwCLgXOYGxCCOHm0Wq8K77BhxiZdyafumMeAsDMoMPzwRE67e0npTpqCuOG1N
SJ6BGhF/wmri4eBAekUtUlpRgM28TOzGRZQc4Tsp21JTOIb9VE657KekqunoWWtM7WgnRsSxA07n
qL1CGRaw9ZuKbpMrkIQAXe48v9qVQITIFshO88FaqaUlJAHkV0ZEEh3lr9Uo/BO1k/ChED6bebSi
vU0/v8zC85SzvthOVPMpfVkwsNCcQmWlw68kkMRDAQ9ilUlzAi1XG7xMOmRN7R+Nq8EQy+B5AE5J
hdZrEK1TBwuJbAx7aROeS12dDgdBXVfoAp05hBHl9m26IfQiuBqxpqNNtI8fC3jutoC99ibvc9/b
x956vtqDa96HI8GSJwPI4gt+VuUWSWFSknZCwr9P9Q7VjQ2UpTHNm21NirH/3+M6LXIi0WakZ1Wn
E388GhzxWC5sgmn6jk5IA6V5Gjw7ain94mIgUGanAzrL9+pjX6zdxj+E1wxQm6o3FvXg7G+fJvrI
rq/Nm4d+6xADSNgtgKxXoIpaDIsz+8NFkfFu5xfC54Prrguq6pU1zGPhb0FMNlRL2BiyvKtafOgJ
8xOfpdnzZlzjh44eML4dgcOj6OO6lZNDS6TWxb18htHgWpzta9ojLlAm6iNx+cbTjC4Rybee7Vk4
nvzeDKFULrGT7wwP+5N/sub8mIEJK2jTzjJ6f6WMWgmZuyYgf3lAnOor+OM21iUzB49rwzMmai9j
nqTY8H7FfmaafvoaWXTAqb7BdaMU3//DQZnm5hiJgbHVueXdq+PLQhhc7uf+j7XXMPATVqIItzFN
PRAkbv7x5zMswNkbqQI22G6LSGtO6Fs4CKNZggpg0/5Hgoi1HDIPvJWTaCTxIHIRQ7RJVwXiAp1v
A32UM6l6GsTBJIzEXFoYo/hvv6ck//Xd6XwJva5FFAEbtzw8d8CkRiWrZYDrZug1CXf5twjMTGhx
6mC1wPrGjnXFe/etK6OJFKYCb9NTNxlMMd3s+3hbrG3/nrBaeTE7wOHjKrwQAwPxPMAFuloNwNcf
OPqOsbt4fKHlwKLOZcyRr/yavXMBfMfq0JRJr2/Fr75FNEommmd5qvcfN9uhl5zBIkW2mm/QOiJV
snG8sMIneShRqOwPbRMrUWDx4QbRkrcdrDqv9PEVdwpLRVwkSdf45+gyR+Lnx9MVBlI7grpqVIfD
HSpOmiQU+SqSDHDbVRT3K6CzEsa5viO+KplhHPzaU/B9hL0z7eNdMva+OIXGVhFIR6rMQ3Pse8cn
+WfjI/QkUnuo0zZmx8i9lWSQxzoiQL7QTucW2jYpfROBfVlrdCzNLFSui6QfrWSUKP0Gr2m+tcOt
gjuEzAEuCOwS8PElJD7rL0xrlz5bifoxsNxSUZBpuEqsr4JsJk2h7jiZSAaPhqY3OurXVNyxOYrs
oDdF3rUlyzfrkrQ3Jcz5REOExpPJJZPlYi89HMZ5EUkM2S7rYJvR3arlQE7fzcB5W+lMssxplrFb
Z7k7p3MWeGfc22xEjZR8Cci8jagLIZN8HlwglcVZvBehxKKqtKo5iSYKC8UoNZXiUk5QTtVPaMQm
ChRhRAPed+V2xeiknvNrrDlUQpSPqMiTUD8Cv+72P6Dl1+3gsyAiJ6zDIdLiWt/hZIq+WKTmiJDe
Gff9zCIzIsIBMnoNC4pg9xPRXiFCimkuLUFMMmzqXaE/ToeLBHv8EFC2Hq0sdbA2ehxpyFlx/U5W
WwrTIYkL8S84rN5gvCYA6acie2JASAwdH6FZi7S36GxVAmWwMgvMZnJTvSfIy43aWdsGngJBJreb
te20xlUERtxbSm+BMbhoo/BtOboW5idsRs5Xj7Scktx0X1AwpuwfLbcL4dGLfotAnfJFVi1bNWvC
zRM3GTWqV5y7nnDqFdkWR28SEMy6pOKp5bXR1kQxIDRxIOfVyfOLOqz0b7gMX3Yve6YGQPj0nVyv
OHhBg3C85UHLADUIf1Z5SFicnwvkM3Dp6Bk8XSloriw/GW/bSuIrZHoA+YmiDguQ/xlEUDG1Yj2s
zLrqGel1zGjRxZZL+wpGqBVhj1FcPBW0hbLbTABcMLyNRjmXE1hKpsQFZ6CYG5+y8K4yt5DzXVxe
qKoM5ybaxWqMbZgUmYTEEZmMnOZ08f9CclM/wONEAIdUO8gcr6RLHBUss4wVKQhGuR3mnZbDCjkm
fS4QA1pMCuTv+RLJCIivOTS1CqNc11CTVVFxFbkRA8d1KPhfTe+ic86ZGg/X85UHqfcIuEfO43uW
EFSx/mrzfuTYlal8oQhmeuT4AJcziPuRWhoeZYAfNRychvLIxnLD1RgblmXOO5tJkc/TQkcrN0vV
qrLKO4qQ7wDOos5DYRaNUL+USAL6rZ499ojb/rZo83pd8LVvuBBq++YCrUJuzPhMWtVaUH6JiZvi
V7//tdAZFTEqMXmgCWBt35hsgPg85ICb8/y+lpwgCUKYvXrD5rCuo5ubJuc9e8WapaVP4MeArSyp
HOLqEVat1pyyRl694lqjuO44B2C+0iZv1AfyzAOT57BulIAkDjXP1bOXoJ97h82UK5XH+ppBCnoR
CA9ZCTiCgRLIURp59D5c6mJzs566PYG4kvJC/Tbbsvb905blvipBRTzYexZGLhUFEDCjlGlhEcZr
cpgkVYRmL66kG4xARIXqYeriukTvJLQk/LuuGQfuGQP2RabwFqSdyhBoaXaa2Mr4++M1YOmsWbJn
EEckDV88EzZ4qDHtO5YbpFGHC6CgtLe37dfxEuscCzg2JgwNTmFMmihHNVl7yMgtKFeuhWH2Htcx
1eDBJMiiA22vfAzmBiytEk16J0Y5VhE4Ll7wIfHAZfcwYJ7NINs2lWUw0/r1pJ2tmZT9zGvSZxBj
a6P7QWDOsQ7o8nureNCOHzKSMgza5Mk5pSSlNehUFfVEkdMglSN4HHFp5IzmfD6Ao8rJzApLDz9v
u+xJQyJV2p/M3wg+3lC9rkAkd7xWqb+U6rnOXaaeprKj6p2Z/MupDwB7hg3MMP76tYG8jYcvF3pF
6PTiBPM0hFFrwm5DxwJYtMx0uG3yANm4IRShk2rZwDFu8axO8Wd08sR/joMB4uaFyWlDEB3njvXa
EVjZn35DYVJfPFyxMu1UnCgiULrzj1hs4OmuoSdQgEu6JOOQ6y63Q7K7maSGzeadwpoEjI/uYh9h
YZKAnmejayvSxEdPmKtBwnpheBoU2buJ5U/7a7F3Fr56aBs86z8+y+5gyW8O4ZrW9jJRhHoo3IEX
LPv1UfJ37jARCL8P9NhgE0L91oWJ7HHKBnAoAo02Nb+5Gz8986mDpzW8biGh4QoVSdiTVCaDJwaL
4Hf8m0tumN96AOVh0wtjxAWiF0pTdTUihkjqfzGHVEd5opUiL/sbOyAFgbyQh5qj5gNri01LILoG
3FSd441s9SQ0CLPiE04n+dD26U7ATlvSLQx++pQRrs6rwp2V9hA+Qfy2LR3EPOuMgUX3QTl1ijU/
T0ya5IYalgVwd0AvoBcKZKhE8UoHGIqwSbKtga1I6TSEK9/XJg8/e0X/bJqhM9y55PQTdK3gIcfM
A91dxnca91lUSwaGg3pLgvPGIpaHZEyBdDZRaJPxPyeeIiCsS5o90LY4kgcgyf9tn/oi0z5j2qSI
vb9/WekCe2Lcs9t1XhyqsFnsMX1P3/brm7g4erLUrLPKSr4bF5QzrKrNNrTcxm+b3vw8ohnZd79G
KubvE1zoegR5Mv5S3EkQ5qM/h/okN1/A60pQSMgMtKOg1oTy8TVmMa0gIHxkmmcpwGqoR1V5xedN
sQaVWAnGZVRf+AZkjwYZJ1TT6RI2ghOaePRkqYPxuUhj2TVxsjVasAWSNYDAouUYrQfUWYOqHVge
KPEL4Gkq4dMY4/2XOPGd+qJepMvJNiurjHyWKd652wIRxXLbMc3Ipqu2zzc8LAyxJpm4/OVtPOGE
EjcgSchLcWWHmogNext/w2Cr8kLz3rdcMaGB83X/A1gEBgWb3865RqRhtfGS2DaaT1kwj+1aNr/z
VNpU7svjVkWAN1m2kvmnUjALXJd/8OXf91fyjGE41E1aH5Ipre/RBvPboS2s4QeJa2lSuWAnIVi8
oFRxm3lptkSWvSWQ+xFyN50rfpIsMj1sHw5K80O1xIchIihaYDOGFykjyg1WmNhnjMn4ILSHP+83
juXFqN33FbpCUgFs109SzcUdyUfA1zVupi6/khaHn9gV9Ak6yiVVEXuQD848RCZyLE+eN3UEGwCU
HNXnT0j0hdNGsLXRzpQ5kirX1vFV1Q+/0P4kHjRdvl22RPmqiw/t/iqxI2xFhNHk4EtNhWsP9CuP
uXrNn9/jIq/8R16vjgrjmEnFmp9RX8YgZhyyUaXfA6sGZwsnLBIJoWS0oJY/PBACQAr7t0fgub31
YouMu354qYcSKpznvRX039qNqSEJDq18NHk0Ir0MY8+ixwAVtkd/LAQnonGyd4Qm5BzjHgDceCnP
1zCvdRNGFRkS0o/4uzOnTFd/bLkz0oGJ9Ts+YCNFqoBwE0/aky8W6tOIo8frEVs9CaNBnrMpaVH/
ahZAT1FLgRESoEqAN2kqikoDIxPmvRAesh9e0ckOEbDr4kXMMzAcV+IHQ1MeICrgS3TTozO9lAmw
Iar+3H4ScBeFe+9lc3Y7+Lrb572dqwx5sozzHjo8qhYvqWGaF4/FLxMQB7zeACE2xzmeTL+QqdPa
Ld688JvwgXc5cMb6/hMkqY/8XftedwbrESeTrG6JmdFicGa74vhjElky5xiC+/09O/zdEktHHMyz
Rxj0jM45n+czyZAncqe/05SmCvobQcfJLMGwiNqzTdmpe7TuEjE0p10Sz52kNzsraO/q8Bdg82D8
rBBc/+AJNl4wCzoAYogB0mVp1HLWOQv8val5bn2I5cXBf4UiMgMRqFxkNie+cDPOfoHbLi0V1cmw
BdOMk6CCeFy7EyzjNEZNOLUXRp508vRmKhyxf+RoWDt1r4G4nDgNbAPCY+eGU4wkQ/GGSM0Hga3J
yJdXsGdMSj3odVLz4yAcLsoqnU8bjVxzmNereR1OKsgiF1aJsmdn+LxIkqZF9waY9kEk2tg6ZmUy
4qudWGZQxpDgYCgH8kwkHXVajX7jnpy4O3QS5HGlWiYqwFO7Z8Vyhy4aBYoKRDs7PfKcc51rTUtU
sYtW3L4twaagYVAMWk2679w7L9KSazLps8UzymD75TDP3ujYCf8943LSowB6I5e7ahy8ihMZil9B
XomueRhBiu0+byyELs327ETmxgMEM8/ZCAx5ofKt6Uk4sPj1BGLOByHPlLUT+2kd98tGrStI4ru0
GeXynY/ppru2cRde46SjRnkf44nBiw6eaelW9f7eoxFjniwkkv1nWlAJJfgM8QC+bbf857ykaQOV
TRa9Eq8k9jXmxH6N8FPZcRRzCWPRIZIxYMc+MI74Y+WVlUC/5eU03ICzjZ04o1geBGIH0E8rYwfv
tV/fOmkKqWVMkZYnrgUBvgl+ftpyeLO3zaDh8K3PDCD1c/Z3aDX9DHDqbWVHIUElnV4WljveTQT2
fT5i1sWLixXBtli7lQUYM4bN5s2JyKnFv3eB1IFkvsc8NfXRLShlET212FBZw6uamzZZSYSR1//t
jT8iZGjnA3CYFXkot0Q26pAbg3FG7t0fN3zOfFSfLqy85FC2+8Us4z/IB0acTMT8SR4i3yEgrve8
GyiZuFdHFUGgxFXny7356CWzvDSdosfgsxCkcvB3mEjxubFsIH3yvmeeptIJE6Jd8s4FKq74xaBB
7sgHDkgTbwI72C9ytPo3uOnCHhhFTjYxkocYHQxvTmCec5XUzuGexX4i8sFrYEObGc08QGS3rUje
1kBB9IdNmONwJ3DAFhtakoP5lDBJS899VeA78166Yub4aQncl9OHvBtw7MXkhzek/I4+vcyWaab3
ADscGLlMZDdno3qWSA+4fsgkpmaUQuZi+ZWeeazs1HN7U1b4fCz9CGlnkhoNddls0Df13/hkdDcd
WAYOOxfV6ytCuFXGk/n/cRhde6zvFiiO8LsPCnLlK9QiakxiSaqbkn2QYomRHpbdGK19TG4r3xc3
hume3ps6JIVCSvzszBsGbQ7eoQpxtRqVlGa/CNtUVVu4fpe3RVGKwzrQ6eH19XHy0R0R4u1CgkkG
m4N4siAr5aOVPCEQj9Xcygwz/IacCkqnxU21ONnQiIqObU40FgjR4pNa3JivMevBuywBFzymnq1j
df1ma9+OYXb2YouakPM8KyJyjJDAPvhivVMDMzBZi3nhtvktClpHsSZkfTw0JLKpCwJ303y4JSzp
9qsQMtfqBR19CY4TnW1CM2qSK1EmvI4pyoZZQyCsp34YOxu5GFjDH/B5EYINTvJUwyVc1+fkm1wN
kZ4Z2fkAomZEwteyzZ7LYvUX5N3pzbZHDg4zm2am9vPCHSjUYqI71NpOJUNoDCpoSRMqbBzAWojj
IqyG5looAc8NfDoZ6hQk7kO6stU1W2/3Zss1hPmQ8Y0MIwP3LAH9jxJ27qFtXaW4b+fImSoZHJMp
lNCQ5FC9OQSWdvXorgkD1XAF0o0j1uFgOjcRO26upgtgqklJ33hIbahP6w6rRGfq1onLJgjYAaRg
Ds46/V9REKZNqEiFyfg8NgqXFiG2Ra8KR/95ggR7Z5RyeOMkBes1n4nfNcJECuSSaPBIwK2FGiH1
FlH3G1uVeHXgi7P9y+ExfAEgu/4EufW9xMvB/ba79cv2/3V0E0QInP6MKeZtz77bQWw81qOMqIl/
U7VsUjC2KaTf3P3nh3+dToORg0GHlYYUX2D+Zf2CJM4/8f7wDe0DZG7fbpS7DUBrF7jS913zcxMc
9abPk832SfN4JLITCmi0GVTR7ZNKlCTs1sthI8IbA0N4ue8Cve9PJVmO3lxoATTtAB4kRUJLit3B
4HzQ0hTYHITnArzYPF4vWE56k0h2aeS0ihb+urfRTrROWAsfCwOR0VZ42C3ZORW12M4q4GUxbJz3
mXGmR1MvdjCccXt+vKYAVnPK8oNB9kH5yMd2cLczyDgaa3MTPhGZIp/RnmNEqmNEeWZzorWfoxYW
9GGrdEmEhK+PlN9IgVT2nFut7gnJMfoMiNqCswYPxzS1CO3QsUADUmibUohi5HAF/1MnFv/gHdeG
1SinXSItBIDOH0Z7+P53+UHp0spdlJyILFBF+35XHCk6pA+ETxCsESC3d2k0Od4j8kxwhkgus7fM
VCDr1tzpaBoxLUA8py81t9yxwbsf5xt5vcVPrv6++Z2zN9YB0QI7yuzkeQCio3y7Veqqc7CR5jfd
zlrhQ36sZBn9zE5Wjy8AG4+h/EliykMeTvmlA7sBllIplpI7GVrNkKrNX6zJiH6BP5WwTPq7CO3/
F26LdLE8zu80GhrBtdt6lIvM3FfWKzr2U4H+XvKBQsVWZ+k0w05wsjtxc4mfhiEVE1vojw7Pb+u+
A1WTCIgcy5g/BXAUyqoBZVa5h8eVfAAxlpoRoQnNpFehtVvm8LC+7k+/qfFGp0zVf22b5hsKswj2
exSSmoZr+/U4wMpWIHz7ffeWhJhG4rbzQ5voJ2j+kWAOk/llNZc0DvO+Bb0sbZ36z7D+MbjzOtkW
UqDx+K+tJ5iOV00VEh0PetKOo3qGNDs8iNdvg57cCYCCKT/QAszN8hxI4fXTKWabPD6jhPXbqmCf
2a58PWfwBE0uGnHWZJINGAqmETH15ORXBkwVtvYBtJDquxlc6j9nGCCddo6rgolOnMJYSsc6x5A6
cLNKMgSHwpnlezsd/69nCfAu1DsvOUEbpcWsIv4FJp79q2KbJhrQ7+8vyr5hxoLd4/c5fHG/6c2T
tkSmTJ/ZgNsNdhAupelDlC+Jc63Dg/nTt9CaB/Ww1ZB3L6+xoWm7CC0hfj5d+HYWMP9RjiD/Zycz
lQbr7cpFlbVlASFrjigLKmPrmiwbauvyegUZSsWyXjRU/vY14VuBa/a4NLBBTTDKm66Dm1YShNYk
4R0ub+Q729nODQmqTuEvOZEJA4YK1fPqT3jNoGfBwcE2jGBlzNgYGBm04SIKeI849LbUANgLq8qw
SPf06LVaEkI627yytYvaBoFFJ0m/RereYMSRPXhnwAm+RVwH2tGwgCLsCrZlL9EzTHWZCJGUSZls
AYSPVlk87BA4BKofGyfvpOFNvGGiypAwn9X5r7UkhfYulhC3hIkMPnUO9Gcf440foV5KTPab+ein
kgyA+UiTkn4CmSYrfslOQeRRrwamvKLIVihUcJN+2UA2oNa2LuI8uTllPPaT0vOJSy2eNCs6VWPB
zs+xy++ZfKUzAiuSXniuvhp3684DpKgnOpIb6EYzhqYa3ogD9N20RdlOMF1CcrJbf2+Ybhe0lxyc
ghb2BH/n96Ojobf5J1LI4x+2JG4GnZt3lvupb16moJ/ZBBSQVLQ3gscy0BhVsW53cl58TGGk124W
7dHsbAipJfhf4qOOSMhd+s6PKZraNT6RZbSWPTmUmtdOmxSd1dXo++yOPCYi9gheOS8EMXzw/4IP
eMcT/7ItqiByhb3GtThy0mi5tTAkySvACT03rDXS30Uw3wQC9U1q2zYKenWN0ohfrdZ92SsA7rEj
f8moQtJUJOagJIq2/OrH3d2MCHVBGwHlAgvFLsudIU22wC52rYktIedSKEy5a258IXWoXlc4fW8t
JmuLNV64AmxPuBiZvhD7fgSep99TDCNundSSju/L8w3BPLXazaWrtvsEaKdiZYR3c861NSb2Shsl
HJOkGftk3XwTWgRlX0k2f59wiehJwt4Oa1haWrynK2sBzb8ODd/LxIo/EGYk4BvOQzE9+uV8M7l2
hDjZcu7ohNUZIP14hnY3wvmMHW4CjayF80U/crjRimr3Y6FJKWyXl3Xa6YhIetOTkIe1M4VDw1fC
xEwFViVFMGJdq5nF9+NqTOG20xKB/p0kHwxbr4Li4P4k+cOmM67M3iJvquIGSCr0EfPz/AcFlZPD
XrqDRIg9g3YtfT5S00iqPJAj7KiVO8F5qa6G3FrRDT39brXrDFOGKyodJUW1pmM9I4+PTZFsv3v4
PrHpxdccJQE74EAmZdAG1Ij1KJtWayPWZuPq/pQag3nmd69pjQ0bhYXKA/J846OlfxXMaL6ZzHUP
Xl6O+8HdXoCUuYCpEJFsIV5JWfge5NioNsDCQtZuStPLIxvjxadJf/E2FsReGaoniNjn941Sn0kD
oXTseN1w+VvPN88cMjSgZoPOtiw/iO2ovFDd55pS3hxiZrG2n/fD2sbfYUcGGc6VHVdWmkd6EbCx
TuIJrrTsYOgHYcFfS6QbY+ducLz6CiDo+9dlzcynoFk7vyu46gLtCAlcTctOfClUPSo/jV465299
j+Q+MKPPRN+9TwzHphqHptyuboZ7Lw8Js89117PS8O8mQ6SZtLTLV4xz+SjIQQvpzlvP0WFptJUD
6ZqqsnUmKeNchqoIvMjf/XkOoC5NW7eLVe/cGXkm2PZTeuUYcZ3MwJXqxxlWaKtpMgqFfIjQ4L93
8O/JROtyGR+eDaHXWcvCukmGP5vLesyjtpj75JBMD94lX81FguYNEF8Z555u4EsuIyprB07HOwpT
5dxsJKuVQP3nufj0UmzHOfklE2HN5JokA10Ddx0sTqMvD2NAWm4Ih0thAS+2a8GiDinKiC5ba+D9
yROV4aM1SyjNmAmgQIcN5Otff05zaN++3vd6j4td605YvQQg8/GmSsGHNEjcap0a2B4F31O3Agxi
vf9QHpYTjLXQZh6uJoldQijEPnfyTBH3SzPgWWNCg9AWF7fG52M8K46gsaTzuKcpRVDIrSTyWzom
l+EEmf0Z7FgEYuj3EO4pbzBZ3oFZN0rrLqhfppc3omXiPh1sK/PhKRHdpY1oulGVqqDz8iMszFVw
vuHqespLgaug+jZ4g6MT6oPnJw28v4M5YC4/zA+xSEM3cIEjTG7dseFh414MlbK4w+yGxeIQcyla
rCy7j5dG1QsJXLRMs2WwjqXwnR2HgHeZ4TPMZ380xvWNB8XcKoLuwRgcsUBdSIuUoU5PwPeXR9Bj
pSDwK1zpo6O7KPZI+Tb121XBOMotruFplZyq7VwKB7qicEo1PJiLZrZcNebWyzEhA29nle04pELZ
Mz+z6nHixFCcJ56uMmP9skGjm/mBn8lu9J1d4hPfeEpUR/5ZTSyAYWLn6+rbLh0hhyDW5TjitgyL
IGAY7oKrI1AIhoQUGRGo5VjGnS2iDue6bAKIyxeEJBE/41TgpsLqvd6O2lu1cPrYOiqilQtHUt/L
KQh6kWZOfQv6CymB0+RB88eOD893KRlUjMWKchOCszKSjIoqU6sse3ST34sBro8tbJ714vvz4zJp
TAXPer59zMliq/FnekxoqgcwF/TKyAFbtdyzKpwdKk8yprZvriMOnyTizlT1KtFncFEGLC8NRBHQ
DzEEQNW/U672PjQ7XEyACIfy4IHSck1U1boCRAvt15zMDu5k+BmZv16Rc9z+PwyUjRnjaH0kH9zD
3pR5CJqL9V7juSBdHIxMot2xU2ZcX/gQQfaxj1H30dTj8efNHfX1JOvk1DeqUpWXgvh4ZRvHmCz+
7W/3mtCxHx39rHKi5one+Hpu2PYy1pmTUzA9YaH3WOFnZ8OD5BPgIhqy6zjuTRMwwD0nxBMd1TFy
RoigHw79Ep5zOVGU/HIgefCplwAyDjajFpNL3C0ZFikhZSOiqHt2ESBsNJgQzVSHd5SSQJyQTSb/
e2mtWTcj3ippMSUtDyjRkXLh3l9yeHK7XmTSzTWCZUklvYjGMLJJeRSaE0n7jseGeZ9Bk12SNIBq
cEqHgDCOMnH5OL90R88XJLTHpXHSfAuwPmn5DonsV62WMOzLoPEJKaOuo/eAuETiuJbvGbnceW2i
U82lWGtvvZgUu9JXgqklZpyo8XUq1nGrbegHH+LWOd1NABOKwtMsfEs2EckquaRla3Hv7XR2rWtl
C8lDCYeRXTUDUfdS1APPOimLxz0ptDsqyi03euLJhpf6yz9MUrXJSHuE8ROscPvc3UsDsz4WzKwQ
PllGSxbrL1qCSXqq+UDaSaMfQZre+MzhbVb+yDDgzrJtrml9rd3LPyWpoIWFzocOrOZyLVOuuuo1
5VMbMV6kXy1jPQKAOXle45mPbXGtHNm9h2kb3jVG4CNLqt86KEOSszS/QVfo0AUYELShCHDdMyen
Ie6+QKO1jljpYsiW6xX0ORJIFh1U/Y8drSd0LZKzj9XnSqn1e0y6RjOCBFH6ER6RMsufGXA33TwB
5/EZs5CMs5ibcBmU/K1zkIb0DwXrjBv9Fu/brb76YkWYRanHn4F6Eyf5he3VQqoCjQxZw74HGEzM
O67Jb4XLfzyB1Q0UFvoPpB6kB0yqcFHw39AHgoFQC1gYhWI9UkbsSlxSNvlg0voybogEA++6eHWG
Cs16q8mJwr1GHGpx2O8Ewz7sRo+m1ix6Mhc/mOWGOANL6+9294BwfhQ8rdbYSF5F/8geWmrZzfmZ
TnofnVh2VNZ2Q7CnDj0WCQS89jqr+77Lp3iYxbQXbiBsv5X8WgiMcQy2CJ6GnaZ/9ud2I8pjWuWx
IlfNYKYa0gb+uOfvz2g3ky4/JchOd8onNw3RCJTcWzY+mBeamFCFI8qC+I+xughl5ppKHErWP4pH
67rEb0hWw2kKDDKAfB3RQOXKhXjGkT0avahmf8tKk/JiTVyu7GVTKUpAxro4Hn+pVjkQVSUOiUuK
Cz3rzPlOo2THIGBgWQYV4KOj9vZsowOG+OALtbZqjr9sMRSuOIwMEZv4+aMpvCW1ruV3wqln+Va4
fx6zEFduCx39MbZxLxS7pNv/PbbZRfLLaGDNQzx7CipIQo1zb25869Y8nEtxFTAUNqSTB9CNTawb
PVQ381weeb2sEYZI23TzsvZllyP/G9aB3xYsXSXluWoMYmDYSRoRspyoi1wEDfNy9SS7uPB3pjl9
djnSiYpVLrIHgBQzXfgdQGmzVXtCnVilJZ+dZEUdYC544WCVQPURmD26B9/d1f8zqCw/UVic9/jI
E6xVK7a3JO0VeVVa8m2lbcEgOp6FQ8hfPcF5I2VEl0IBHCnLGdyStk6+i3WZDUhZJdiQLG7KGD3I
Cx+hUGkQ5+78C5LOOqBYHlrqDdhsJjnWLGEjYivDddAVsfEzBNTT8eKWVfBMMY0TaL05xPXfzwsj
Z/pc04GdukalXBXOOibZxJZkDyQx4OMX7557ClPtpBqFo2uDDVKiVKUp0aLEn+OebrgcGuUXqfus
lUOZDjbteBYnyVbGRTENQ26hFHZKpHyH27tROlEzhlMTLKCOtZbGO4Fj/w/4t5c6kaQBYd7f2eIX
RW3faDzwix8eBBg7GqiyfF7wqEm2Dixz2qzazgme/M7vfGVi67vxoEyx4iYBekVhGqf8zPEaiPW5
K1ESlxkQqrWm5YRaPF8fYwMKVz3Cxjf5tgvLrImBmb/wkyt+cElpx7dEhmtxSAuJgIUChI3Udl3B
CLEfhLzAhAF+WJoU/3bx17Y1rFKpnImFy5SQqF5IopE671kx+Qev3n6WDU13XtaUhh8CkhRh463v
c6R9UWu86HNF78gCWre8hucqNa77MYy6Ac+X//6DdGvME4PY+zUdj7gbsnV2QRynUbZMw/vat3/L
KnX+9wsxYuvq67URKZ5rYKrqd+j99LTQkJ1UfdxO+m8NHSTote7qwy3qQtGVg42CLFY8T4vhnzc/
TLzjePy3leIxleUZRlutc15KDPWvUrubURvezsqajhySbD7mTybC62JMarSJk0Rmm4ofch9wNxeE
BT7fFcWHVBCL5mX9m0bgBmHAFlS0lFw4s0n8fFfiGNpw8wOAsVBxAYCISbkUGGrEb9cDXMOPURCb
+8MubW+KwoO29lh962COGUq6DVYIy3vbSlidATNcGxDTwfytEtTObqy5BKwoD3btK42QzGSYiVfC
OBEIKBKJ+dPDLqGdDG+QDJgWeytnOXGD/3o17VNyNhzJ2mPnHwdxrQtb/Y4kGzbP80+xy4delKHa
H196pVopRKUBnIT/lL1RfrPzNxKalPSdFlqEhdwU6flSA4ZQ88OH6TTYgbK/hgHMNkn3fFKz88YI
jz6AV2e2TcCjMvETg9A8yZKG6AbtzuW1NgGjH8IoNK+P7igq4KtfqnBdTsBgw5eCUSBj8V+HQaTO
JyUPmQAggG06rI/UZLSZnXpVTPfMjxObVnKiCL4DtqrQNpt1zo8L/q52EyWwnACjsaxiAtwJqDKo
qZ/J/A+A+Vl7F/ly3i5XFMFtV6sKkv+bJY61Fw2qfA5yFN6ee+w6m3pjbf12OA853PPchX9yW6MW
l541Xng7aQBhla41vwNv66LMZ9TdFen/hGKGm2RARMNbY4cPa5BhpAI2TpTCucOMq0YYBn568XAc
+9OK/Am0dgGPXtOYl/tDhtmrVhEDZgjUanZ2elhu5PPTIw8X/F8jdllYktVFTfQtpRz3Kv5zn/d0
7fG2JF/zo9Lc7wG3j9F+CLO7GJbgPZlTZQ9dGCTrR1UrrQ24yevFEPsyHdSmWX/+wGwfJ2Ez6dju
TkiIPnJFlwDghDnCSHfcK5E+aC5WWoki2Y86OPfArAuUs7MVWhVmp1Bnm0lGrHfHlQSOYqjG5u+G
pKRLjthrtvddKxHrdSN9JgC9fIQP79YYTprguF+jKpKPPH04TFhpn1DDiRAWVgZvQWGbDsyFfkGD
/c81okYBGxmVo5IvMu8jaTT2E+6rGTb0qtpxZ/Mox/tayvhb/gtceG1qI0Y5xDJSc5+/boKUKmIf
K5KvguSOgbqH8b8vkoGN43LZC8G8BvSJ7xesqxmApBDD0vYBaV8MZdyOGQpDW6poEyWooN2UNfbV
rSFkVcLrSuX55qeXc2VFdo6sZTdZvL6brfNL+caJi51LvVBnXH6CaVgTRo04gp060+7mF+2zvCmy
qF++/YIXyo7VBicvjkxiyC0qtNHW1jqX19bj5yokIGnlthe+R9rrhsTxnDN54FeepqTqtdZK2WmO
gJmRwo7aZDG2OS8B/vAYdHlS+6qpHLY+pXWKN6uJSwZszmsLqFqObcHNdBhGUkw8KwmvNjgNpID9
QbJoEDCRWHwdUPySbo//rPiCnkvO04JihgDNmsxmncUX/VCs3KYKESALkY3Z444EUXslVNC+bBx4
9TIBKjyg3pP52OIIBomWIyouBDp9RBpr8xk9Xa77ebd33fY3fq8Rqs+dRaaSxWREJTpcL3G4FGv0
tEdltPOMhKc2Cc4jdr7LyUxRLXBffnmofxAxxwy4m0M0k/GCKOjl2EPX5yiKa1EHRfsdwgKcFDzR
+9JGAR5rEjCXGuQ+VDBmcEc/gG9k7VZbJtuoQozBni316xv2/RHV1frWZOvc5CmgiP1P8ma8zLUW
LpqmDm6io0G27PSel7PlFlJ8APyvnj716gI3KTfjd8RB37e5B3fJq5kGIRs4OLXlja8cbI7YceHr
WLULxvIpc2tNeXNrSajMzFqGHuVs2Ncwa78VmM0VZTIKGbV6cmEs7x10gZlRRBqvy3eqtP5+8/jh
UZ21ExMhAq16gRxgekZ0qLMjf0th/HJb17zqJFmvitsupoL/azPw/oiIPknw6MClb0TW57ZF0ICz
pavXQEK0F088cUTF5el4Y4V/HPDV3eOp9YOsDww6fNs89Uw9jslfhaTtI0Vmk58Ta1O+L+p8LT6+
gU6mojVCdy3Ic78bPJYyNrM4/UhS1OfvXYh4lNX3rlcYh2Lka/H/4JVvW64CHhIMqc87sbAP7L2t
hX9mmiJH6uiv+kkFeo4zBf5e7Fa9OOe+AeQaaSjum8/4y/f4uCZU98sUbgHAuGcz+H/xrvzNIScV
WWTK72R6raj5V6qwLiPpBFtfob0D+bUVEQgnjl0K7tX8eJtal03RVbNb352rXg5oUHI/wO12tn8+
K+5RH1KXIg8TK7S+ehg+nPAmU7Cp1N9tNOOQ3wNsAD5YZ/j9SnhYPGl1AIHNZWAhQeVpu18M8K8j
6BIdwehnwhmLx8npzqan2GMLIf7ACO6o9rkOmeOxnS7PifBzKO9/U1iGCICe9CRt6T9bqu76qr2W
m5FT3RL4UlGjFFXJFdDHZyRqSl50551qbi7Pk7hcwUxilxXBo0zF76+Sp+vysRPlB743BeTbYW/p
tLuRXbeGgTQim8EJMMf4Z0Pih4OWHiaACKyMQcDOwSbYZ3MkgpBemDZuy6+VdsS8E57UjEPxlWdl
Cp6Gswjly0tFxW9h2xg3SLHBCMqePxKOBLFiiFceQd1rA3YTqv3xwF7N7ZvQc3xC10rGA47hOwZA
shMEMb8kz/FjAcuedZ32oO5ZP4/OPDGHAT4zImuViV+XC0cJ5AyVh7Pu/ieLl+kidVlmYLuiNOLv
X6x7dcqJFLyUJb7Vkye3ftV25ygLOyYu5W1xoUeTG3zNZJDKJM2Uc7QummA5pm//FA81JK9SCg12
O3IHSEdpYKVAal/zb/ra+8eXMyCJM7BRSfX6n/kQY7YP8k6sr4nEyMuOdW7coFhlx9lZ++VwYeRj
ATaxay0NAN25j80hbvWrW36aQhNGqS5zl7rhS4d+qEw+h1HmW8GUhtpWNNzWFDo/J2NKe9WWyU1c
yrVp+iTRoajwB4JG/PxgS9AQx30oRwrYz1e7S1aQ1/1P4ledkIWW2KCj5h1pPP4M5DD0NS/Nbr2H
sPX4lOtU36iK7+RrgNYLF03/XXUjnWkC7qIuaAD/Tp+ULfHvxjx8EEs0bppsuITyhzwTlQDcrMlX
ShU/9g4m2zIswQizPj8QHRxSk54gu1KfJn1s4FNQ/4DTAflpPFke2hKCI1GP5TM2MgLTml9FbG9G
I7lDVZMKGHj8DmGdX743WLavocPhWFTTZYd7uYNF1bXi+WBtke4nc5mr8XCRdXg4nx+B7mDrG09l
N0qbNdtmu5MCU6lXQTfCjhX/AzSAU3dGKMqP6v+5xoRcbg8jTQiVF1XOJao2GkZS4Ebx3rMiqreh
vy1QMaBw9qVpMqzRVrK6MW4S1VBhHoLD17uEy7XHHnqVYJozBHz7DsrQar4WJE3utHN0Pbu51QAI
0WBixkr/Xqjrdc5bOe0C6qWkLPPUR7MeItNXsms9Q2Fn+mkWhmaNlQX/ni++rKO/WgNrU3EDgUw2
gFt/qvKcNTxGDDXtn6Sr67DGH19u/WSQZk4yLrXzaYDGHbiGsXyrZ9zxFFNWjpJCChVUgQ+ftqrM
wQ21I53juHLLpaOlSKmw0+w5c2R1kSNyyvOvo+tmzmc/GXEDlEpOQaQjpJWPqlBPqU+8s/hFqt9d
anRQK2eqPis6rE45TDDOt4cWHeUgYXNFDRoW/lyuRzJdLFsWkjoShhK9jQZMP2gdIYhPeVdB4G6i
b6nUyDBFux5VLIm1cIfP3pA3J5HfVn73EvBeOJnqoCAr5rvSio64AUpgQ45kOBABkASr48cBDFZp
2iJgxm3RFsQeVCbVMhwbW+o1w8iyCXnujVWGu1TYUt5h9dxwtgQK1Ig0/y8xaLVzm3BbtRD9Vium
Pq00TjmpzWH94Sbdmw6ddfm3EqljCONg/jEwFjWzQKm/E8V3v8y+HU2a87KtqSRzZj3nbuPCBCRO
cy5cI55/duscBd5c2BUL1yEOIXNmZziFORxMjoPL7sOda3WjEyy4ZI1qXV7TaF6gxNWURuaJMfEf
JKFKeiTKA3wkX8bTOPZtjyGwARJB+KjsGh2VJbxOLdgboQ7tVyOufEh3A3kFYn7s6Rda+M3GFd+9
aSXObVK310TVOGC3Z5dK3LToz0DH7FYeAbainrrDu9whhaPiRPYIRVLxN4inFzaohguO/2zLhNDy
uP+Om8cnm1q536NySjRvO8tn1MWvnvohASZM6HsR2w768kPlNcgkPtOs+lfVPSp2qYFJGoZ3wEdd
KsHv6FpVbVvT0CKGe5EL9x8/xNY75w6H656TCaUQFdY1sw2o6sJvnOaR2VFPvnnrK35gMvjAtlzi
zLIcvs4ZcwtQbkKES4KpOfMdJ3YW4qdKfBHne98Lbp9LUtCcJX7cNqnaDVJVxaSU6fZxfhZmKhXA
RT93V6KOkIDiUf0bI2Aixi8jl5rvo2nKeiasmds0xenj7FSKpBUKVUh68I+arf4yy2/LX8Dyyajf
QgkottU1KkKoer403241hCSJbK254kMySdm2PT96oXWkBbVk/WJ6WxZNmAibcQc7E7K2fydbjf32
Uze8iAs9sQWqsO30CIJPzDwrgqYJsGPUJQSCLgk3EI/UiC8B+SWa3UEu063EFchrGKOTJz48xsGp
cCu6yI7uUHnpBIhj78IR1KpoLYOd9mTz4ZlZkv357qH0k5TIEbEuVTR6Q1xRCdj6jO1V/fiCiV+x
VlcbsqSS7GbqNDXtAwBEcc3rWcsOpk+c2v8C9hF0DRAK2ZhROy/P4y7VkK61WEvf+qTMO2axEHtP
Ku5bIeylhdbIlP6NE+lzLATOFXQ4nZnuxCqnckirg6S+LYnwsJeV3ueBhG9ztj9b5ojUHM0WGAJ6
GBEYB+qo0kw0Q0xD/sub+QTuBY5+IzLYfeqR1Tn2tubuK7W7ABnjpFwB5jD7woOkchOj34tGJzqo
kXNaKi8PMA5g5WMd5WY59fRR1ABTbsiH9Z0cmyYrSxL9AsIDHLhr4mYgYSPIE2vQipIBplsNUWVY
PNUOmSNfPL8LjV3AUujO4Xj6+c/x34DfJfqw19rF4P6iOAW1yMTlmHmrn2nu1o1x69Td0MGyxEH4
wg8cUW5628wm72Lclg6P7INtl3GwwmVQJ6QSLxeiwpz3I1i8EqP63KM8pnYkyDtGNEQ85FAa6IGD
uvjVyXEC0DWt/4yccO5TZ6Q662Og4wYJMMWEsm7PH+lIwv8hpfeKhRQ7uxkZ80iCVhHep3XOQOIX
rJOCQdoshoKrLie5F4tWJGa5Vbpc7aBAWHekwIsVbMB45N9JJAUwnQvUPQNJJFwORXaiYLVJ7K5R
O/mw6SxOpzajd4FvqK6R4XVY7XbKOVDo2TB9Dg0XT7PaDgK0OSej1sCNwnkUextfkmtPUcAJamad
t4cO1h1aJ4ZHsH462x6xVABXjsYIijLiUenNxPdamgtWBdxBx3P22Hp7KhsTpzJVaMkmGhgV+6+V
q6CqU+phsKTKXSkguO8e/3GVqXOjS6CmU8Y7S+ZeaEihzfylOgliTIpK0AwfmkQyI+aA0CP4PAN0
0AHScTAEpvG3xVB5WDHlZjL+aJTa/8cekeGCo4hvTWI8DT2xHOZDmr3tYvJp19TVv8IUwYuGt1ZX
5PfGLRWdG38u3Rp6O3P8Cv/bdd3jEVHNhmMuSPxePYA2r8Xu6+NqtShanBRP3ERJCOxYQQQTdCoB
JnSvxgnMAUwWQ51ju7ehF/LOnU97EWK/pHg0zf8kM87okYltMbMsPrIhVewJyhrc/DaHwkMDYxfr
9BGzq2ANm+jAJ9BAaLlaaz8pja/6vUvdA3UJINfd9wNlOShvJmbCJ76/u5Ivf0BNcDqMZ+9mj7HL
M7Z5zywAdaMXVDFg2kmW7AHJnMCGx4ZCs116omou1teuLhfEkyD7yA9f7VRefoML5uZ1zix7VWFO
C7tdaWVB1Q6MG6gyjBq/Kf1ez2iEzqcx3CaNnH0942t0CIMW27vFoFhiA3FAVjRxPDIydFa2SBVW
11TQolMuch+2odJXA0HrRg8OhWtrGKqqsEozyf/fzGvvx1PDcURMm2/4xITm1+Xn6jz7PfPi6Wh+
Px/aJGxU3RHd16WApd6odZ8kygMQfc7KL1ik/PA9/nN2xbH2gx/WZxOjR0QUZtwZqyd0fVXfyBPi
S9FhngXRldm3Lc76NxPN8hGV9Kh4//oDRfez1UWK0HdQTMuW9L/ycHtwiHnXoLQPw4tYw5PDlE4X
tXd+j8nvDTIIhnume/RjkW0vhTPQqrMB4nwW7bndM0qpYZXJf3ns27qb5AajuiaJMhBAaOpDfd64
1I4PzvJfkMsjUWxoZfak+YuvNoscHCpQu/cyoojbXdIw4hYpE9PwnAvf71bYlhWUN7TphQDvEGkQ
Z6B9PJBifpi+GAEVlH8VQI9prjCQ0Eqr1iZIJ3KSsCeOz7Q1eg2vg84DkMWV15xtTydr09yX2hqM
4uOrxqYwM606JeNcw07N5EqnvzsAScY04JlXFvWb85lcwGgVLjV2oX0OY5tllGisFzdpJokdnhKb
AL0pVXxvgCvL32gpUSRjkFEy3kU3DIumPwCQgFqoM430mtx7SIAZbUVZR+McH4jWsPryFvpAB467
2r2zxESBGapHm619yD7LU7r7Dzs7Od1ALCD6Nkxvy6vQQ0Vfr98L7dGoLkbv2TjLQtf+ZBKIDQ8v
bJ34GtlnW44IEdUHLSAhcyClb2K8jn+HVERwAxwwgrggAKgw+nrApWbocnyIVDhuSIkloaAlhakU
bRR5Rdr2d0X35dHUiJi2qEvzw3ECNaVSHTq66obCsEzYVUIHw0PME4/5dzg7yMVr+MOq/rhFHwbh
o/tmMr7V2DbbBTtJ7ayK5Csge91Hl+0B2ALOXDwpyE5FFSInXlS8RKUGyPJemXTd2nqHUr8z2X6I
/7SFVMlttOnlOHOWTWEp6pG1PvJMLgrjHBczcy3Qegbfq/VOmDFeszvsHocscbyZdfdMtOZB5rWV
Na8ZllbgE0AxkuXPQaGxvnxO5G0sefbDfB4w5a/ponLq67B4unTVNBRRC4EIx4BwVxg3faL2rNWR
kYTaFjq+F9yRVrTtT68gQIKTpMxXRD6Ks1QIwoAN5WO44dcjvs12eNKpeAD/9zxYBgSHkW2npDek
r0fEmpQp0mTEPpaOh1Bkp3nMr8o93hdRnQhP3sFlxzVZb8mbr+hJEcEsB4ytCoe96ZSaXu6Dq188
xC7/78jhxEOcgJMX0bKAziHDusVWY4M4lUptlLX+5wx3oJLvkc/Sc8aqlb0w/0pCtt5ove5Y6BnK
x5uEa6WInVTCQZsJAryzOysFfgWItaOF/JJPZlvfq8vpI7RBSCEvc4BII8lcUhtDQofvTgkz5+oi
6FGw3t4V5VEmiRVmTygSKCy6ku3WqfQq1Wss81rFJWj3O/dbvWzCRB3aaKh2yesYpK2i18wd224I
DWCHW4ZYO97bbP6LesrQ1WFZd5xGcIpiqqaKlwlEWcDtVkV6kbHog8HnK59gepEcsFDVhxxmpa6B
WCONVLJJWGWBd02Qrh74CEdBZ8ZuPgi7BT2hSSijzdfIAWD1TLqJW0EWBPPxqvyHzKXXMiU7Wm/D
tPaDlnZqYLCZNQ2w51ASNBi8pkl8j2AQz0qFB2mjZxwJYME68TFJYtK6QldlFY4BECvGbMyNYqtx
FJ9iwT+PyzPpbRsSOKgBsXXOeURb+qHSMzRP5XTiF4Il9lX0Yb6nBBOYofS6p5F587acsOmjAQuo
7wOEHGSYSzk/5I40SMuuHNMsLeGCaVZORcqcKbAen2ihtt56LLJEr5PPMsvcndbeQgfZDbuMvJRs
aIbT0ty9kIlei55s5Zi+rVDfTdyLESHOqm4VKKp2d//DgXjLK00SHAOI2BWt3G33YZW2OvrRgtJe
AXYJUWamlrQIKEStsY24Fnq/lo3Ir1apT50mpLv2JRscuGY52aO11SfBmbvKw6sY3wZke397+U9i
L4aElBX5Si7jhD5v6YmC+D2zViKy0O33j0UbJzQMwdjz2jbbL4UgbOAIghixbatzxJbvHri5OSzH
3BZRJ8/t8HrNTool3viZvA3tZfXq2jfb2kwzU+VYIzn9Dv3zOHAeJivsQA5xE4l6sKezejhMCVLa
qlNaoSLUv7loi0yKPbVGJ0x/r+55zRJacNgVI8mEPJIBsh4zl0hHIU8xkZH1dJFCd+shCuXsztlC
5I7PxM7iV85yA2YLQ7umkHcyRk+y7elBEYscuG9qwwpJWuIQMVB+vllrYLn1dpxNhdsJgFcsTItZ
BHp6bn9FsCCVQOh+YLFuAeCP85qIzDMEiXwEkVSyb/xtFf4jd/XsssAYecQ697YRrC8OJcPaIIaG
ZfbE3ExtezuSMwIklNPOqBwh6Bi5NiYzPk9j+EFDoCW8ol1S7LpEnSgSvfMTx0aF3d5K0+BxOgSS
og99p5uRyhvuST+AExLKP7wjps2+E8KWen8zE/MuvP0IPsmIRkFQyymKa1GQapoymBtE3nbjIedU
BLAItFceBolPngTdmC/1Nogzpg4w93O3BtN84d/59rSCOsYPosV5CSIlOKorXsb+IEeXGY2Btl6V
ckvsfr50gox0XIGsL9fKDT+nSIROEHuZoKGLImooXZ33aeJpA8bLSgZpzpK8CAVqvmWZTcUzoN7c
pnjbHsuIJfKLYiMdc6G+Dw8MKoT/KGHcnF5jTAnu72aVCtP0Z+1UDsC35wz8jBCdFIDqVS2FykY8
Vxu7B68XbfEQXa3SC5EcGLHxvrSlnB2lyl89Z0oGDOxBTrabss2bSXsgmjZw/vfJ1a8l54h6Kj0h
Wzw7wq7arA2G8Rza6U4sj/1GfjmTLdOvQAzCkIQJCj4+uZcUSKzuujM7pitXyg5DdS5P7Gjnj+p1
rMYSa3likG3P4e3s9QkwSXYT+kO6SUEXQTdL55gKIl6JwGco2VuA4+bQVyaiXiKT3U5VJkGDDEv0
bFOrIXA4cNmukOeuTnzG6OovUNsF6XsZPBaHFK0ETKrK7b+FWGIKnp+qVvXCUCMzxEPozVcZnVua
5/Fct10vYqiKKbTfesnc4ouNr440jAzSq8RQ6Asv4TsAvceH1zWOQB8PgkwXuUY5ZI06tAJMRGTO
DtzBLQErPDIVavITKOESsFnSX4FMJJfqkoJnrR04Kk6CX5amFjRH6Xoi/d0tgLVgbggG4Mcr8LSV
yza4bWNq/eATmWbGzbK+gxuNxPhJcGQJSgaaSIpMGKKxbo2SXroxwdtOSrjsUDU4ihEQzMT85U3W
UKnWQNmS9K+RnlSW9Fz9pCNK6KMRe8U+Nga8uq0aTf06sX5NuMiK3s3jALwCzweCt7KSPdHb2Npc
nww3JrPZK4cxHizNpzh7k7ydCzhUF8C0SwHk5wT3hE+GovTqHbc+vxsQ0hK63u+88Y2kI6V/mvaU
9JCqaAdgDietRJ3tqpas6inyITLnDyFHuLE5vFGU1rqLwjHySEP4ZO1u/bfsP0p5N8md4mcj+o+R
3fLhF5ZlSnYwZL10LnMfBT4CtwrTgxX4fnfjBA3zBQ/7lF3XdfgSFlaJ1DK1/XuHyv8GGHS7Tvcg
xHcH4zIJMsJg1DORwRwIwcdZTm4n35SyUplhn2eBPFqPVFqVZcJPowJ+c38WJw9fy2vmQSXPquVm
Bj0jDj07mj8HkHyRjUE6GfbgwbgP3kg5zMEw8Q5eTCYoID6ofb6ClYKocdW1E/xjJLWsCCZFq3ii
Mis36Z98VqhIvUwVkIAkVNTWlr222D1e+WgN8+arVDXMksOdS4i34Iwb+hjaQRqhIqPMn8D1pVOi
JFOYA8zjbRyNXwS5zbIxlKjHEt2uHJhCrEaeNV0D+vmMoxLS4AYIPWNrDgP2O1paFjihdWdtCQuU
gp6R7pZOEj3P7TAJ4uiDA756OtUbZUt5ejLHp9tQr0+6VJSEO06vdiR0lIh1aDEPlk+S/28XGDZo
hk3a5bOHJBCkE0KtdDLvhgxICViJlg9f6tyc4nge4vDmHocA9fQMkIxYQFi005VRhEQI1283O5Yi
6bavJgqljaWtU3Hm+aYUflKJozBtIgjbqd4+pQYVt6nXHWpNdpwzOlRm8fybu0rZeH7eDz3l6u9k
axme+o3DN1Xtkji/fj3VBdK/nDLBRtdDQEnQ57MF9/xm9T6XprFCNMuPrvcG1UvWcWD1XAvuOaVU
KiW++E4yix/bxjz3DEHfcrOxc4Sd0o7L0j7G9Vr+k9/4cVcvY5//4RNrVP8kA85Ak1RdkJTblQzT
Y9LGfHtL9PvVji6j30htO892dki1cgyuX6x0sT1qGgEwej7sEQq+i6CuFV5YQjnJSgNbG3hR+ACj
NukSzrWwjsMC3kxtrIU5edqtvPXhgAXIF22wDTfMtq0vi/d/PD0fiFGCvcqYXeZUYcoBkLOqO+AN
C3gJfBKOkmMgXxCD7q+XNkeP01XhhHt5xAbLRK3gqaQ1H8FE1kBSX5p3USiALB+0QgR+zsCAhQya
L6ph2kphdw+KnxYf4e9lM+ZXwIPmCotIZ3oNmV6Y7+ANgc7JSPqwRqKZ4VJFwkMPFOpew1dzSpRd
0benvlppEaDKQK45vWyBu8H/7654w22fJn3TzTIv7Akw/nEiTqN8BqQLpZ3eHr7tBsBiJGUGc2f7
idU22ejdkL/KHauDX3SyBSwroUnscXUylGqRsEa84UMNVNjFPZCtoI9/IDIq5/tiu8GJ1jqZA7Jw
9PqEJciy2+G2gJ9fxsZ/u7q3NuVCy7gHpVRYN2KNpMF/pYFcVdi9pJa1jAKM64TDb0lCDnZ+jmmz
cVjMOB9NVLoPp+sb/o5F3vj1PUhVmWNu+U1zF1ci/BIbo9lvGrBjAVvzFgsvUwFodb221xN+Lp+J
q+n1Nl5vY+1BBDOB1fGjrWzT3us2x1pYEySIcp1oRuHmF4kEp10s8Ts3pFaYZQ6je4WeFaU+6l60
fIRMki/er/bptmwfAdzYuH2UiLZoJxYOKnaPS0gjUXC663G7PGNuuX57YAHgfKmmRgaUwDhkUQJA
yQh7aaXKrA4X4weq0/JpO2qUexodhxocUfrtGKEsa3IOlMWYKqh/6gMZbEErB+JOD5uePNdIc80Q
OgH90sKgj0RpALZVE4FHMU3o3ux9r07OmlbC579rYQPFSVxnAeOq94pOSF3bxViCahNgLsoO7x2L
bdla3HNpnInpC+vnuKL6a28uZttrmWlUCeqCLWjEtQ2Uvr/OgsvZOLJCKB4Y9a9cruM+nmzantRA
68L2eHZ+h4cbqY7Z9F8hXSMqlB44WLQ1V952Z75c6vtdmGs2qAtqh3eV+XoLH9lr7B1wKvVEs8xM
U33k8/PQMebbI03xgQy6DlINJK+ES+2UVQ3CmxbPg0RJSuTXEx0MWr+q7Ho+l+sI4rVvNL3ZvLpX
WD2UdTeB9nZs0WJaF3EQKceCWOjfx6uJ/d3I2031zlXFOaxqmVte5ghqI3EXsGskeVYj7/EE5ncW
eWHdCJ1p11Hy8uFuQQRv2vtd2IRdivJw2E16oAGIzfsxdKnvtBNn58T7RV67rwmJdtS4AEFH9vde
omYxnARlrt/qPoa175oTbz6SyGQqNsVotTj0yTOx0ZOy0teE4exfp/GoFN/qFpXh8kMhj9mrk6j0
u7GMSUOAu2TcHqnbmkePs5TpHWbQyTA1WIaxQXuRtuR23yNhq2PdPRw8tE4vQZmpYS3Ry2p7SDAF
MFDlHIb7RYT0nNUNYTnpCgyPpISsqhd7Ez/tuVWxx4sY2iJwuqe0DP9DGtVrbjOn9LlUlEKLLuoh
NzpEe9UhGNG+Ls+Wb6rqfyLJoxbk8C8E2vG7NSX9XpF/7I5o9nVT0U6tyPV5GY+S6VheljVJanNV
atKRP43ZrIeHf3vCL9/qT44SV7Ygfh8tXVT6OSpPwgjIjM7BEBGGAsYAF6e1GFAsR1mGlX5bS48x
+No1t2VbJPt/fJiNcNsEqmA0qEcNVeVPOeIN+9atMedZXuR/3WODcZQRBKwFoRuGAuAqv7JdPCVM
H3zRCtUMydBJ1qax44mCVVxZOdtHr0zt6E7hXbFPtMczntGGzdpoODxmduaIXEBzgGTbe1fRzW2K
GTOIwG5/LRknEJS1bNRx6s5fGRM+2u9gXbZ8PVq9NE07sorr2VQioWxG4w8KYXmetyrNkKFJyDe0
iZN5rFgu+WBIRuU743f2UM2mM/3k8BWDxwLhin3Rby5+OThJo3yoEatkTb6k8FXRpxp6QC6uMyhl
J6zMHiDMsVLkrWsmNZ1wAHeoHQV5fEy0xEb1osglE54/uwNMPAXCacTHekS+eCa2Swvm1rqBGE1Z
PiLgNykdWHdptwsXPo1DykN3luJNNA9i3UYXsYcqnwdagwBSFNe7Ll9rQoVgyi5jdDcVts9uFBfn
ypk4oV3ueR61JZEwqeQ2kmgoAQO56CvkjBwMLWMVulp1I5ZREH8sleJjovDdcIf3J/9toHPZaTMa
GUqYBVdWSYXGv7f+ZG3h/b1oqV19Mtpz44nlVQegqQWYvyZMSkjhvQcGgReujHiKLUoTtt5seRos
EtNZr3sOneiLEXcOTecz7jHJuKHsjVGXuZsDpHQPwULsLsKuMZf2bTZMQ5if9lR9zB31z7x6Kt47
RV1Ol6p6OEXY9yRLyABdAGnIuWybB7+R3Ol5KdcbHttIIVKLCiJbtnlOULJGnqkSA3ZbGSH6Jvi9
3uEDG9Xv5bMxAAjfseQw0zHYUt+3zKWJpOa5R6RoLb788sHh5qdZ+D5Mr1Xin7IF2mRbjVxODJus
wtzT0nsJbzlC2eZeVS2UhWIzeTgA9TsGVSup33tfDUb0hUsF36xmWt065ONJnSG1EZIif+RkiHv5
GUft+LwhYFRI5HxknVIBHxPqz1vZwGDk9YPcMkEfjkrLZ2HjI9BBRvJXAR+t5ruNIMMRA1cJ+bZx
gKlPhoPweAaZTWd7iRxr8eJg0r41PwaMW+YfSTM+p7DROhvWJ50KtKbWR6NweXKQ3nwCmuJU91aU
q6s/ChXcGZmiAzYN3gBL37CLNHvYSH0yfQjGICSKEWK95MRk5sSbz7QaUV1DTy6mSr10t0yJFmxq
FSL3YzrekJrA8+XzTzbimma5t6SsRzFg00qmhiYVflYwVZ+iLaHnIfzunAqZnkICOkMlz4VizNpo
P4xeKf2gB2EYqvoPORKfpl7qbZ6Bd+zlcTpBvlb/E3HKlVKdF/eaKdhDEupULeMFRglT+VhloIaT
LWapbMuXJju8yqgAeZNR6o7vgKGEprcO8ZLGV9s3aBeln0F5xzRsGGnX+EyMddhtmij301u+VTQS
Ij6C3DtqKXbnu2p1EaQrYO7C/nHoadj245wa8CpY/NTYrM7OfVsme6DngSe7O5eg0/wjqlVZDo62
ru1B26TYaXOWp26eN+LVw7/3VIJn5WAzLdBRKYBbaHKD2LSUyV4wmMA5GpWWD4RMqOtl4uw4W1fz
JRtIKdxgRG9ip/CF5J94DuEVHkLFEKg5GRsiT4nPC99MKdUwqznvHr9zQ74Rz/1AGSntYNHMB56J
COt9/DDLs78t+Uuiol2StHThJMo+N91yptsSLvv/po8VIv99rYPmoM7VCmFrLnfdMOVMIUdQcwr3
Is+KQQK7ix/hGqad/L+d2G4Kq8+AmFUJDixz3e5f1a/zb8dnpRKtxEB9zX0nGFYCgITG1wXgPwB3
T+Ob4Rpyrpx6fiVn9zswaiaoPLgEONU89mwUzEAYgiXYgnRAKJlKhcsBY3A9TkiuVD4lj/ghEzHq
wNnIEQsLdAH57TJi/KNp5ztMpd9hwLJMygyFMR24UzubulfcNKyB9f9i5ctHR25njAIM/t94KWWQ
SkV0lQdt4TQUhoI7XsVpQml0kyoamCSP3O5w+98I4ZST7yWP6Rx22v3wzSTmt2kfk9iXn0+iZkfs
4zGycJ2S5McinRrs61KnRRolCIur0TdWSsVS+pquLbflAPunXQ8JYF0osV2ZDxXbCeAs4YHutB37
Pxovp/zcSKU5HJ2c0AEIwlRwTi+J8to+H40GPZd7myrFHwvGoBqnIEyh4ft3t1+CqNfufq5HHNBb
LIxpRcxe1SFIATFM5EzLq3voMdhj2YFzCU1H7l/esiiZtdMvEFko9pGc9PJVOShQLEjSMIpRIeuV
JoKLVB1x/Z6kfOOzABukV2gtyqHtyDLOyfqGZFXNIIUONdeH16JkzwlXUP3fj9XcFBIJTznXPbrD
IAYMgsOffPsBCVplSrIbfCVs53YFnvYywI3z8U4Sa2ZLQD5WWVUn/iBlVo2/wtAlrilbUUBJ60Fz
hGbtiBkzbFZWwgRcRz+kuMSomJn6aF2VPb3ravxA1b9QBvowGJ8sAD1mKfCT6sNaV01YI08vEGal
PiAwWZbt3b1el4Ry9niw/BPKm8Hqxsk6ss/2NsQ2TXKclPDbtmudR7y172SoM6Kn5sHzF+yrmf8g
qOCgISAJLbQvlzQgzWMeyrSbN9WZULM6j2bc1bLm7Fv6Z5DLGhkJYrSUlk/1Ds/MF1gekZQzjzKO
no5p1twH01SJtkw/K1uiEiZWRofQbE59elsDkNz+mrTiE2BJpRp2T+KlKcpySYER7G+bIsfAvJcB
vbDyQ/+4ZhhbVB1Bnb3mUihK1MBFmQbNFmW/hIXbVxrPKH564vJZpKsNH6ftn5uE76IwNIYAg+ck
hP4JiQlOw2PsCfoVW1n1cjKFYqhEu+5E3PKyvnWKdhqC/hoGZzAFiEOJKH1z/yuTkylAIoP+g7Ch
4qayty2N0ckwh5xST49UlDz6u3APBb3u+1gmSlQcGcwG8WkEF9g5JbqxBLxL3XS4uPorNSHZDfMO
nTdASybEJ86rKPASop7MBVxlGXGgtJ3kAHajP7MRpUahPL4d5bO+yAtXSQzGJj7rxw5x+u/8NdVl
e9DWcfSgO+jQgNMCLsvAO9ZRj0mG3/3Dc4M5Z7SQ8dcmwwiD3sHZLpXLWFUplrf6emkpwOvgzSjy
JsCAXDCOY5k9lxUsmn0kbBM/8dTNZ36cc9Ot69HIAaOCSyZkylz8VpZ/wKLKaW9SzstOCk5a/oPt
0x4zdO+kgX/N8wpooLLEiK8K1EW3lCcT/gr/bCWQP4sA436JIE1eSOeLIIjMQw4xEMx+aFSRXPVE
2o5SHWs+UM7Ah40GiGBKcL5C2hsiM4cVpBvfaBrD+CyCHvVAxWW89+Rgq727IjieIDGaal8cyp57
1SyjCGxpxUbu1UyCIiiYfFXCGO3v7haUL4yQaQJuqqLGiqsqBqKTM7SsrFNIJj20SxxLtFwfk6bB
hQfIqpNMzzvdvMSyi6zkGjRs0k685fIWJYN7mrVJmGi1jDS/xnkmZyYo2mUT9lsNM40vvZlys+S2
Zn6OT2DXbIGHtFvDBgxTPhqdC5OxQBGhA2l+9par0TlqiM6uhn7LQMt1nV6191K9lgH3L/gaUTAi
aedOm3Jv4IzZX62fK6daU9b1j1VlTm7CeZPOmgoWegeUklhflTVA8xw0vnxpvOGDzKbkokKJYFp4
d9BCtwT7WQDaxq6zokWN++tAsXzZrfDZWikPll6UYvccPROxG91593txgUFF4RsqLF/rt2plpD2+
KSj4Lblj/EDK2bnUR4N9sD3dkpvTgL0/bftwi+4Y6gNZ4+7lb/T68bpAVo1tj9WhTeNHYLMHq9CI
MkMUUddwAp2ggE5VQ828ZdRkIcvo+cFJwqEAp8hXxXgbCn7jLyerm2ByiJITOBcoW+mvsG7H2alx
2a5VqyRfPyPnkK3dpHgH4cmujRAAJkFJQTLiY69O0JoXz6/CfffaIkpwjSnotAbw4Q8LTtafoz+K
IizmoWOj8bmcVlpii8OK5nFY99YJvuNNLToYPSv+48m5PzzfjEAEdBEk3OMgVFr1Ghs11N9xNcPQ
6rKsJdpzcIFE+2Ul4tZk3J3LsweR6jtu8A4kBndIR4Q2cXs6m2xuV/whuhT2NwRHW7GiYNNfgFaI
p1Xg3/XNVQT093LqoXBzii2m4aNUYzbgG+IeF1Oeece0asoE+SrARhYIsG8RzhJxvuXbeu0qhwUZ
U+cDN9BlEPxzl9xSEe9pHayHsP9sBBesZpR5AUNRhgx84hi0GffKDeUTmR1ziiZ6/EolntT6Hurx
GQxuMLHyetZIjF3fSoWc2BP9NHNW23bItU5kF3MiegZlL/KYKiDsR5QjkyntwNPmkEYWeUyMITsF
1fNR2U28dlVe+lPxjZIMb5pEjp405osIeEhZIqB889YT1ahZPGh6I3v9LMw4owTFremQl1cgFti0
DWe17qL69kcVJCNVbDH1iOh/jlcJ+tWsf1PkthXuGm0+tUzu7oT9AYZmL0IRGXxMlmSVdd7jEDC7
THtvzjlItvznTcvnl6U6KNodNUhHzogZtaq3WAcTadgM8/yW5rE2RmTJc6QMk6QO9AxuKY28xtA2
SCIK43aA7go1l/IJYrjmkvKEDE6/G8eyMbPrNxderaJEwz1jIQskhyUJdagyJesFsRLCwcKa2yVU
bXPbY0pCc1s3/J/tvlPMe2OQrHpn3KTBFoQnksJZSvuFtR0Aj1gGZW4w5vhZcHVJIOgmaxPMG1x6
b485SukoXqrJMY1W6z8BIWTALntarAWj0w8MGXqi2SJA4ubvwa5BfWs6joKyHhlHp6wT+UP0TgzQ
B1f96ytgtn16+F7wWUf5GgdIK930SchG+46Rv2eKEHq7jhwgRCGKMeqSrSsag0yiq13uiwDSjvMY
r0ToBRWFbktnckzkgGY1TrOWrV+dLV7iYUdd6CaLa8sJXxSLcJ6PLlVWfs5QBO7SdqyUX0T4JSU5
q3CnC5Q9ilNF7yURXqwXX8s8i8Sy5H1cQxyOFOm1LIFy2v0Zj9sTfSFgqn2bEMLwm4uYPXXKdIrH
/s6YUNqxrmKTa3WKmF4IKEWid8oWVGO24SMkTJhEuUQhy7ZCifpOuCD6O2XSZDuh5Khx15SlP2d1
zW63FefIE7OUetCanuk4wkSVtukuKjag6O3zAy5q83RI3hDjNrgGejc68k56NiPD3V0l1AgOZOtK
rtSSr6v3dCTk6/6jY33n28vz5qab/P18rk9RmF9E29mHpfEaT85CUmscqxpLSPVu/UW6HWlD8Cvd
ZMj7dV6HAo5ox4EeIGShiz1YSzZJVav0lUaTnjsubaNHj2jZ4zltvvVTK4Ylo3dZWxpdbmkYe0HK
IBlCuHmddlrtoQ9S03LifAV7vVL7+nvWpWdZq9B5LQx4ZjDxheXqqxhXiYw4iJlwgrueaHoziDuu
HkwGjNOeQ01KNt4zEH6HM+4M9y6P4wVY3rKkMzAujSHrv25HVl9pBawRAIuXZhstCqjAeJJ0WOYa
ot87F3gG1SYgerjpZ3t0LdjwH5N2ZMfyiwaunPqn+51+UMCoKjlM5Ol2FKTuYmRRx4xKdmwcCAZ/
eObQ+VJyNoQ6Dsg/PifIy8XYvX2n86LBcRA5PgjOD9wacnAqMlxM6XspA70k37OwbcNAOH+UGPSJ
l+ikFB5u5jHz+cBB6JYi5vZQ7OsXHbcwBOQUZs9CFjbjos7uRgkr6I9XrfLaU6T7N55UrjfpoKaZ
I7f/jOnhivG2eiYE2O2ICJuLcKQZ90iM+twI2B5VSfcU8GZX4xUenKqV/ePF1PregQGxI5yYX3IQ
nKVIQ/hS7Orrp5p8B7E5LP4HqzJyCqF+dzm+rRUP+rCew2+3mpLgn6MwsfKN1dfKpkX4M7v+LgQi
wgpB6Az+blSqekSrOfkwAstwa/IBpggJqjI1GmiIJQpc46zB057J2iWLOA8m55gDwBNnL5Q2Va7l
Qsr3oYclv5DhupU8r8Og9OVxz+/l5KaqX7e9BOgmDx1XH8b3BdgqA0PgizP8isFOwyJdyIxnxFlb
rk4VGvhHCDoxp86Cp5mTHRfN7DloemRcuN3QiCmkOFEHrmnVjG98LMQ8hYAxhlFRvSYyVLwub6Ug
mBPU3kV3DnCm27yDrR1+v7FuFpWeGPsumgAHnS/ztNXS2cRzjYX5V4ScgOfVWxkdDTDbRv1L5Yc4
Iy4UJHW/y0RnGdh2epDk5X1o3zjcefh+AqRSQmYdsHZ56beDFuzbgVwwpbn5czd2MNCkYhpHMdmU
fTO/J9O9HUz3NK9NBYaaKaz5stNkJSq1eKWAM8ZufDAiUHUc+1ubjI+0eZGMFZYAfz8HRkuVzsJY
5EnkzoPtze6oy9bVuE94XR/5WKOzZmdGbhXh5LQhGqsg0Sav/g0AiBlseACaC1D+xNH0xY3M5kux
+3KcFeCxZUwBNIwD468WJIfs3l5fQ62rz9IAo3JURcz817EPdLXsWcwh3bVdZ5M7k891yOO2b8fy
zF4cLpo+2W/Q2PUN1Lj6kC5zUQgbECUCnADEHTr5DtyvvwCGSUdHJotuifUNvgtmdVTlJUwA0BcP
ROAv+lDs5BOwiUhlJdLPn3TA/qimlENgn9yRBMc8Npzwzndxn9jERMN+jFruBAyFRHZwu4KZxF7z
zp2eMD+9ClmNuewqZ4pfPbrA8c0gNQ26wo0W3uDbI7ZJms0FWlHRoBPavC3yzlz4jTEPVh5qCb5A
03A1ysc7C/BhFGcdxor62lR+ywyuoTgGCGTSDmPCb8/uoqaYfaViAH3FZtZjdiUZHIYSxfnwYde4
u+A+OaFfite+bjkMhKUEew/wX3vepxhlEhfU09yVFzwiR9zMq1lQy1Wbgb6ZJ1Emaq2UMKCe6kdQ
4ZsakkH85bku1Za2C740fwTm60m2/Zrc3fKOzN2FlFj2YOxMa3gTKR7qAE7sgPUbpsV/0urkfYJw
y/0qBoB24myUQ4F6iYEXfj3R1rMlZUW+NZMtY46e5Hq2EsfLeClD4SbdYeenxqB03VsRTsQaX2pA
ESdcuWEFoTnSojHbcDk/aTT8OGof2A78HwXDUzsBiGYYHNUzrERDsbHmSSjzHY+Eh09TJTtIFmZO
jLvUgwK1jJ4W9QTkP010zMwi1mAcNwvCtIdyoX/Uvfl06MHHMZz4gSbP84khlxzUkBOhFWHGzo8Z
Q73142q0DytVjbDlyj1gtI8d/KYIMHEtmIjvRSRuu3xasLYapjdjL60XBEvdPvMA7Ywhl3UiPdOm
ykSUbMfcBuK117ZWbqVi1Rc83+OAC+pWjmjHiuV07YY0P9RJN4tkNkRSwzvikZSVB2lpHNREY9kX
SY67xVZexpJONfXXV/k5IIr6lMKB3a7tKhQD90t9tbQ7eT5AZtI8pAyO1gdKXHSNFzykbkmegA6+
KXDiKXzcCwTU3x6lW8w+Pn6VLy2ZO7NQAOP1IqpDdbHym4IGdCquVzTQFVrEtBuKNrmfEUVJAcyv
fB/ePXQc2L4gSTyeKnx495I2csggEHol1K0BqPXx+v+BxdobDFZ9ZTB0BUplcrEpHCqpH2RM7EGd
ZszZFBiOAo3hvtUFwEYYArsU/RwpMm3th+yyP35/uaxx51uaObHlsg9kZv9VBx8dFobQmFYlEAn8
TfeQBqgGTOqQQahoQjni9B2252viItqKwf3MzUodDXfJT3Xxozabc5AI59ZURFB0E8B3VQ14/TLs
Mw9+F1RMk/aPlpl1W9TO8WyXIHKZ5wJMuQEcqJP6rPrH5mKmpIwh8ZmSY5Tf+JBGLNSysJ8qyhCR
MCXbeUjmdu7MHZb9ZXZ6SxM03jDbTWb9KnU7RClPWZaoIgILqf8RCpRPXDlwk8nZTFADds/tuYsB
Siq2NrLVCWJJy2qlDtViinrGNpwNnTkIWueHooTbC6MeOEHI8dFY7dSXaYR43TTZ23vAAVspZd41
mNT59WF6PDn2Qs3W8E+A9cSGPhmBENnDX9gRYD7c0lnDh6ZAu5MIXY9AQNMJyj8Dj1GjvlF1B+lh
bCOhY008z2IH5diZ4kUlY2mvekdZzzgivD+hpoRguksVTNrh61kJXr85WmFskjrze4q5Mdwuf8y6
tVVaYQztD0bt/u1ai0AiEwmwW0THKIxdFwZaaeiPGNejRfkTXDiAXxyU4wNf9TtlQMHpWcZiCMi8
oDhTMSbcGV/Z6oc8cqAHd/GmkP40HzLLTN3cbOHRmhf6DW0v+TsJvkvucJV3PBLwvRlIt+f4afWJ
PRCP7Qd8mGluzmaN0VQWomVQeqbSUNaRPEgpODAxkoNU4WxR/4glk7bE/vQVIR/kcok238HRHeY+
/svoEFBGlnXhzLbPmA90HbfvPtrl7cFyvHP993ousojgrZlgL8avbwFo0igFMjqTtTNzakvdRW8v
h8r2rtHg8/1b1AhUd4yIL+OFjSxt1/6/xfsUKLdxK9qoL77rVnQt6u3YiqlfRaBqx3oCvDK9/vkg
mZjBD9lIT0Is7h2LU7v5BstCRe65ftUlzG6PMK1wPhZS/0fbw93v0ytyDTSv/bu2LfXzAX1egcs9
ogPBQafQtd+ZTj03/ToNBEN1moqVanWAixKR1caKj4rQHhm4DA6YVlwUN/bn7tbByWVc4ye9o65N
be99/ABQS7qgfnRZcevuyf6Xh8A/K3cL1BmMwdydYNNnvYeHMh/ruMvtQjvApCXCREubfaEGReRM
pHCx+u+W7igXqKTDCQd1tuWh9nTgoqjDLpRY5GukZdzCQpPsAbYQ45wGxOBDfrRXCkkD9+FM0MCj
4My2+NTGN9J4eV2sosTh0y3zYFFeJCN4flE2HElGOeojltEYBiiY+Tco6WvVqdwCS9T6bb531KMe
jH36GBt4VWr+zt1hxa5zaGWTZQxO9l7HIFBkE0Zdvii4UKD/z56bMjI3+4VhCczFahn6rwHTdnNR
flwJDEVbCf1asTZ4Sr1HFltLYzGpk1IuBXBx9G2IYXTkLQxmNW81u4gWExJOJ8FeE8GfdYjWOTPx
PyXyrFqotce8K/KZbMcQBJaQcvr+WHRzfcApDVsWOU/AzUjkzKZvVeG6hOFudZ26MOhjz6bhPY10
T5g8WcT+gdAWWXEcnRcrSlHY9ibefouKBJXrL0cpTcV+Pz0wE9FKy4L27gIZ6z3LDOPFOLgLG6BP
V/IBvhn9lW/Wh/ybaCWCrYWm2/Ayu7qa2LrYEjJLpMUlEhvggjAw0pDvwXu7mFSQuJEWdRo10ghj
HeAHkKKvJq86l0WcwmJllwNAbSWbvHFq8tz1oQmk7kh7i4I/wtLIhvnlNSxxwV9Ce9ECbuP5FLdh
4LqIlx8ZeaVv1DSQWANqV/4SW5uR2irTTasVW3RDsVj189yk8tHxhyMGrWyImRhHSHlQcdgFXxaw
AcuWketYXFb2YvuKhuU3GIfI3RYBsJ6lo8lDsI8fjjSo6u8xxaLRYosXGomR/jvahaFZWhXo4J5w
X54tGmqWUYe+Yv+LTvZUkVWS/ZlT6DmfjhEhGwxBuh1njZPVkAvYPFs9eLfRmBUb/vjIeOPSo5vX
YwBYxnAcYffLkVONBqixr4SdLLdp5+6qEP1WL/9huxVVm/C/LqqO2lb1tj8cwfZNnQ2XcLoCWv/J
XN1LbctSxfo9D2RhyGaN76YTnCHjiqsM2ug53xPf49LvNWAA2yjRect1iUVCfoB/SuOrfqjRy5qw
ReMsXp0M2Q49r228pqZBtXzukIaUWXpIS1fJVCKsbs9KsfzEOi80y+7tDcx44pYgBVEoV3G1xxMW
/qGNPTHvWOtyoarrcxPVNP8UjV4c6y7GvJK1C6lnoc9PiWMYUF5opUx3FPFl1jU5S+nFJBG94jHb
rTDiV9fA9IcUuyris6pEEqp//OltGpy9ou8m09hIRsBi3eqbvvUcrh5yUMETcKPDf0oOE+Yz+N2L
bm7eIEPvaXelP71cmL5FphV8hhBWuV4B5yN66HfOIlLESgFkjdb7O3s5jfWm4UifnsBBuvGfLmKs
MYmNmJp8BHZFaTwhS6bOzXQHmXvDxJii1vS4q2SwzB4osCPTLO24f+t8lT6wnykL/Dwy9/k457Gh
9+VvWPPjbF9v3j0ePqT6EBv3QWGFZljFjEuBgNJr7da374P2LpfCHGgoUO0lZjC9GpJt5tzcu5JZ
wpwlJN8+QIHxi4TbUYeCQd/uGsjsmOxhJPh7jtHGd/ZdnsWzizIHrHOjrhFtuEdmZCtdzVPWcL/o
IU5Xr1CLiEo4kISTckZsgh+6lY1NIjrSGIBuzeD9HsfATTLKlTlaT1T+XiLCSBqMKoR6fUcSvT8O
GoebUNK7855lMc2N0G5XPgjgCn4CHaquulA3Scv2SZQj/EXOVXPkEn0F+SVPRzYqbpptn3PNWOGc
euAGiOeFgRejxS9zsHCH2WpSIbJxXSUHktama7tojDphzA3Y/d61bC+P7/7sHUJseWmC0djyOne2
l9eeRDPhNMDHvWXzqoBjGyeh6hcuJwrX7nuQAv8UBxws272WqaWJOnrPae44buyVtzuiTcqSd89i
sonaqLoN/wBdEYZTh9io4RsU5fti9NFw0gvh83iJVAe6bK/MOKhvjtG1ExY0U+cZfUPRCnpp9awE
h1OI7LHwylBNxiZ6IZTLnKiUIWC5b92ZT2xmJqxaGM+rbh9nUSzWdGo7KoVX03X69BZx0IuIHM/n
/Jm0F8VbjNXVJtR/knxROZoD/gIcmhCxd/LuWDHXQUTbqxX7OywAYUA5X5s6zwbs7b3+XagKj/aw
3rUA+K3QHnd0QWk0qjb05CuS0BX9uq5wJzxMI6W47tg6KWgoTLFQ7VmjF/uyaCigRGIFkUgo5/hX
TgUNAVKDjm7iyVfXZgctQGCSfczGLDA+HIMIzeXith7eg4c03p9qLeEwgNR0d9fA/pQUwjvFRTdb
xXy734Bq0jWwrAWde7Rf5w6eTLF5xAnfw4SxQL2ESl6H4CVT7oagu8SqJ5UGr2CljXv4vY1LkfZS
ZzmWF81udWPSNYQj7tzFKBWNdyzXRycj5Vnbwi1Vd9Q49WFzFd4DPQOTH5TozqFmCK7Ve99BCCwi
k3KNN60uF4BCi2Yf5/GuS+tFIJCBg24QOdBDlxdTXWD9YVrLVEW+qF0w5Q2ht138Me5DYjIT469R
eZOObEWkCaP5vksGtMytkTD5jyXqRBSVq8VIjDCL6mHyBPVAr5c0R4m1WfxMK7OoVwm5UaQa2hgu
W+xvQhpQclEdGNeVfrJQsHMkYqNUyWJ+vbOobJF2lHhrTfDOjsZPILm5nxS4cG/N7+BjhMu4hM2F
diYymwBynwDimXTs0bbU/RA9Eqf0ttnS1h7sClhWx9zZLgKCnmJMnO+dmmLYTBZPNi255c+iMHFp
ZXMrkqbfMh7GmZ/tpoAbLSMWZUwKnGQjEuNJlZDuG0yy2LWdsjpBg3rJWe4f3c9n00CUYiflDQEM
8X6JpHvq8M7CrQqoZNwlhmGzPr6QPyCi6DosIhjGqC6rsxgEqzK5RewwC1gsXdyNeI/dAh1fNjDK
ldaqpszYSAn9SZoukzf4WzRrBhBPh2gCJVfXHpRnU14hPirNiVQqOmzvvDIhWqOgiIE0WwGY/OBB
qcz0ciCpTawzD7fLtaDmQEYi9rRbtoV724RXTKttGMtVOs/hQBXCTuwigOH4QZnkRjA4A43i3MSj
SeeMz+2jyuJoTXR2jqQMPBCFqpy8V7HWp4MU03CEvRVflbpEGq/t7pbT7bWXn09MEKSLk8da/FaZ
BgYbIZ+7a2Pj1R6fg1EilXZ3+35WjRdIG6f79v1AhfnQK4CzL/toRzqudU9hE6wIpUz3vMTpaPGa
znK+dWorPCck4dZJlbbv/eJOyDCcz+un3BIQg8+tAWBAaNg0ojQtqLP+G0it3d5rCaXt3kO0tMQR
0nORPVSzBC1MfSNg1GZfe3KfxoS+1F2soCHIwRlU4VDg1q/ZmoqKA4J3/Zi0rpktUyWt+dy5/Wmp
3x1PcwKlEZvDlhL+/aPv/IwfU8LKvfV1aimdYZus5+c6dtnEHyzTqIp/HgJOgXF2M0Mgu2LFQ5IH
MT63+Ecnt0BQouw6FB7k0fyvFDe8cs3AP0QO/4rAOCkiSKNffm3XDnem9lwevQlZvYSj7h84BwLD
flmjHS6caaI+9E8jUVzEC0Q3cP9querjSeh/HP09aKmo7k2PHG0xLdVV++XzlN73xb7S95mb/ZZ8
PWz15ej+VhhmgOfkH48jHpB8XPUqk5p80D8QDzOaJIDrNgEZon1itV8GQiLGN6Om5x9tA5+ShmTZ
5C48ngLlbQOHL5PA8R/G06+Ypbkpd/ZAazY1gKZ95ToeD2KH3uksV8YF5OktlJxyHrA59czel2HR
VarKV+hjd5IpaIOjDW4GlC8fv6cnvqOpRqpesv87pF/SxILld6t6pO0jkpn3XUuW1aUsy1kGW1nH
+sBae6p1c1l3bPwCT1SgInxf7EKq8+HdOk11gee5NL/FzDAewDsUDgTJlBiHNi04Ne8rIaLZbnI3
9XLJlD2Gg3ClHVqLgzVOZ1jcYp5zFgXxoC2Nos8pgt3IEMTiwPuoctlfEi0EvxpLmo4vb7e4tjAS
dpXWiy2L/8IwkF/F27kEEL0zCpThG7b6LGXLFgHSxI109sG9jXrbYUL5rjVLpjnorxzE2c8hXY50
yjngJ94dPB/L/aaJZNv83KWH9TJLioxCJvv5avd6io9SgiHtuOnTIG2qi1Ag5cn2R5yN0gcQbLF1
3unyqQsZejVV8tAYAoyMyL9YONHYAQRFcAXjdTI2rMPn4HFjZThmLe9R0id/61Y1Ettsww/1atLd
cQOLW2kXolmV3qSDYqrCVm9YjZdW2+Yof2q17gsDYAhO/iwSwcM0CUJ0YxtCacG61scVFMLrayGF
7hWbbke5vBirwSBT4+OmAiLVruqpImuGIegNb7mg2WiAeNscm6LqQAZYylIZDBM+bQrueUW/uwz3
zoEBneiIDXAM+JVcbGcwjQ2upBzUXjhkRF+bHRkQnyKkmm379CP9O212qM2ik4G6GOuO1CZgtcMV
qLnixX31/Dmu41G8LhhjBywOBKeTHVZPQk+DtZlbWc8TaSDwJufgr22OmQ29uqVuTrzJpr/y5LF/
GXKP3t79hXpjn8vB/VaXYZtXJq1A364TdE1Mdmt73nAx/SivPfCSkwHT55l6JYcacajCcD/gofvt
E+7G2Zvc3kw/xte+UOAwuDBs6GAemFSccxSxhj6wTuJynwXaCPXYMBa0yjZ8k8aTjOdJzjTK52c5
vMS+3O2ryDE+cPUmyGQkoJqF9FL2xoAHPDySq3t19ZzCqtFyHuS6GQGwFkBzmYzV8YfQ4neH5rQs
KG55CgwzwQGbtxtdT0A3FMlSA397+FbfLEWwrKVTGWmn5Dg7YXYaaDDH7amDW/V7w3Tl++CE8tmA
5Vnl57uAhHhpAmqTh8YUQPdwH0KzUKLd0lBD10tX+qZw41hfgfLLmErvlyJXENZwpHhLOLRDTOw/
aXv5y0M2Qwf6Sa57wos1vLYwfzb4l2eK1r5ovkZJVTC6en7UFetR5EdQIU6R59vue9PkGLiGuSPJ
vlFmPeuIWbbhfQfQSsZk23j/clUsLFtpHUXfd+fnytZNMwN2u3YL8EUI8wylNfL4EM5PvYMgiiia
1qatYEaMJyCiirmLuA26ZW93vL4T6faxlKBrg8DBeti+dwVlmMnoxhvMdb6b7uknIIBVNk+KatSv
THG8sdNlrNtplKXnJ0HDqhHLwQwpfwmWQFt02ll15bRfRNA53YqWX5ZFIxg5+HJfBKYue2jw3/Ja
RaYvKlGGxke8aAfY7TdHTHjpcmZ9IGD+wiSc3TSDiZiiobAwvzMt6/DSjGVdcEsEHGq3I5Wo0vDA
0Ez2oCvxEHt38wmCdiSic6H5Cq4MYPdjjC89RZF2Hn8dPo20jpyOjA7vYrhGU2DxcLfMxasrPCHP
qDsFuqVoXHDtbaEIDGq1dru82XjuH7/goIBvFhQVqiX31ana8rQsr+DQebkQQZ5tbTJAnk5dM1+8
aeXH4SeVi8si56DDeOr7UveToy+bjmAgkQZwXx5+Ky/rS77+lGS/N2Fqfe0FDKckN5vzHyWimlfg
QC9Bi4UUoUyJOYrNErmRmgtRwzGUoOEwc07SL9N7cdKs1lA+jbxKr8xHvZA6QDHVfKyuRjKQDkSg
djHIMBU/0B+j4RFoRKm9+xClZU9nOZGdvvpRBf13uoqnIdTy9Nr2H2OrN2sfXIDyyOY/+OcFhFU4
zXKEI3buMn4RU5vsD5b2QKTEzctpUKpVHw63g1doQr+/4uuHVzRSMh819TZtvL1o0s4reEPG2IDi
/imHeQ25S5PJ8xewtyY1+uKQcl9qTlwUxbVWCGp+TJuze7fOi+JiwnDqIT8bMyXmRgfInY+tftMi
V1glb//Xho6VAT6zKCtkAmOVK4QEiATc4FJjvLwjQ6nXAisu6PRHtNj2soe8cNSc8/vuuCkajLby
bH7Ssagu11h9kgRnQG2Acm2JRDjD3+oQZ9NuJOxpOJDNu8wylU2UIP/ISSRCw6IYyWA/FUoiflUM
bBNn3v7guj3xhs/nFpvKnHY0PDAgdidOwhP2Xep9b49yaYkXiKiVJDtpR7Aach01rpU2kdbzIAkn
R/ccMPivfYSTrLorYC0csSY4mdkXlsyzi6GIDsQlap34/qNl0D4jZPqDL4fModcTr2sSyXR0nAUn
p81ce/q/KV0H6OyVduUZopxTtDUTwpligfIoiDOp4tB1I/jeNKsQgOjAHNqbM0b8G7+qRj9KMzli
zC6Uni2t+IztrKSRlFulVYvktcg5FqM7RXORzZ713SKvo3nJfhWaqx/eYpT4VVF9K3c+oqaifJPK
I2DQKQTs4gKJOjth9svwyBwjzupfC95rxismWSErktyTHL0QtevTe4aW5uJrxc3vC2WOetGPMqj1
D2+i7yVJl5fr6qMsJuPsDUh1oadD7k5zmjZzAdcY21r8/J9D8RiXVIQZR1amL/A+fF9qRop7Icu3
c41fLA5SvNob372ESs/hdyIQtUyvZ+k43zGxR/+5CK91vaVq5uisE+u+wW+jc/MtXJXvpMhzTLLf
zI/2a/7Ernz05+640yVHOSxCFRbwlZ7CmwS0slb9r6QDfLAxLz4m9INuKE/lOmpQgx7Z+8AjrKgZ
LXVwaSB3RriqFUg0x8HRalk+D8gyLLtDToiPuQxgHsm0RtCgfCzzpT8xprHlG7ImounTktJcJYQb
mBU3AvSrm6zrcoaOOL8IgKy2eaT9Jr3UUG3RVhcFs6OsWrwMzaI65k4t3xNkPXmvvYRtcskbq7oa
/5IwvVuy9UN5OzezzFOBMVZr7gmHOhgOKyfhtY3/x4negV+NDdhHCGjmBrLujKuUTgvG6LpfUYmz
G5bj5fKPdwvThpnF8yYnSlCcT/XJAbnwuQrNV2TkospudRisHGXwrAl5imFH/TRXKVK+XsFLHmJe
apq7XMyodojsZwHSn/YY8lnfwdpwyPJVgZijbYCi1ICB7YK/QMs6oLKtQ0du2drh5QdWk3STOPiJ
ohFubBU0Nd4UEzdeqMC7neLfwCLt/CzxIfYPPvMon/HTDIKbKN9tvHfbZSD9shVVdp6mCHhtKtIK
BAaxsjmT2y3ILpvRfYSLHkvgMHfLv748xBp4QeaGPRzNG+UqE+R77ak5hUr1hTBNT9vVkUDAo8jS
AsIsrXiTM9k0tdnRCQrKbTtF2TvfjshlIzb2Zg2pY8znhbMiQ32bhevLKTtXbMDqggpDzg0gCepG
wLGTGx7hd5mdYHkTJXapLe8ezRmB5aJM4fY0UKRylg4CYK7Nnb/HD405m9eLeJnQoJvk40eJh+U/
t4tmhdzS57rdS6UxIYcJn3JzGiljucuz2lQ4XNogUCsX0BZvhWHO3ZQ6Bb2Ry/15dK7NIimIZd6m
IsQPoFYnASoAaJ3+rDJRtCUB8UmIhgiYuvPQmGV5R29q0NCTx+6ONutWSRRkge81ljXQ5jPlQVkQ
CxE8EK1CH+qtQAXJN20fPc1p32UHoZM3CIBpqVvl0meWAGPvbA93auTaM6sQaU16VLAi9RVL0tf1
Pm3IMbpArjle+7bW+Trv3X0FAWbRlaRbdvKGVCru9GyipImc+UtSbcujj/VZNvMxlpbkhU/abOJA
s++X0zwzXDCxJYyY46i4BUufCn7oe4Vm+17nTtG0OrPx7C7c8V6D/w1K4NP+7NMMzKdsV7jw7Lpx
cEt+0d1yP9G0pglzXYHmft2sJ9Af5qNMhRcEiEfGICiH4QqIEgynJ66znzGEKHsRtRT/ScZwAVFZ
W0+EtrDuNlIGADyleNJZCHhJpEIRYU1ubprKoAEtTUx9sfkm5E9YV0fbeBpna7Y91Yj/Nbwv5Fb+
vutMnzOb9bxyt2OBb97/zHrD/lK86GWxvuaOiQAo5Pd+CS0bMSNRRVZg4S+g+fUFnFdEKCRUrL5t
PKs4cQURHCOEse0kd+zbkRO+6x6WnfF4udLrQdp4bBpUk+8WRZT1qXZXGwWNstD0UXRjlU8p7S75
MulMAODc6iF7KaYVIg0lafo9yZjVY5REOcJe7AIVHQo3mIF8KHrG2buRKyyRd2npsOPdw03uPo6C
NVp1mAfOdS3i+ow1jNfrFJRA6MO1CkbiEndd9EmXvIUvbtSkbi19b2BL55ShO/fICFXgyXOAnnh8
9awVcGl0OyC5Z8o+aXTaRoGH40rHj8bhcv5EQKDalBOKO9VRtqv4ASY/Pqv+QuEMD+XKx5hEcQGk
JSM8RuFLAtJi+Mcsr1asfAZxjk/SzcPSgoV4hjKkuOHeU39siUC902MA0+R8YvfwFOnvl7BQa6dP
DebRX+hzdcId69kRhrUEhoZyWYdu3n1zmTX1taBOJx2/dDllFVbJPEpx7TdIbTWFJbpXg2ktYUaL
jyQFCq/4zLbi1FhAi7Qr1Fxk1MbslTEE9+QJUBISdrR5QK0oMk50uH1q3dhRvh3Jn/ITgXPYEKs5
Bo29Yr2FZQtex62eFDpJCAUwcG1EudDONnSTvNiIMCb/DqkUefMrAs06icMr2+9XRHdQebtnD52L
BlzegC5JI+bNSYYgobHAJd3AdB5DEPNKpfmqtD0YUXza05GTLwDc0hCtp+o8jbhwQVdp1XNqROYn
dBs+LD+If2MfZRyqd8hxGaIDvOYDkkibDQCIUiP/EXn/rf3RHATRBox0kyiuV9Iqg4ds+j3qFCY1
hEpLu0qWxPG+PKAFJPt0FnMfv/xf97c7DyinsJDZHZLwBQuUDK/NoXLjAL/QqXT8FeH6FVeDUVVn
nDAt4jg+QIteonuGf70ao8r18/idMS6otlVEKw8o1A8r3dqqjXT7IgiQBEzDKTu6TQsCw/OENfbz
8b/lPqKs7uKugwG62G8vt62cy03PWWEd6ktKKNQ2AdLIfSwiIkkIdXKhrcPhLF9abLQ86D52tm71
BgkGPfOL37TsYAIJhEMC4V3psnEKoKHbuVpt2vvcoF4XQhHDG4lon4/Mo4xcjXkI4dqEYwCYFQ3g
cM4ia0Woe8DgNqrFjF9JSflXfUFaAPYLSxNiUdmfiMBt7HnSB1rLRKWih0KNsRgMY+lQITgDInrs
3gJ6y5BTayoVMSkx6m6A04OG1f+r7p+P0qOEDNV9e131GJTYTBLSBXgE2IVPziejHmqGom+TBXR7
fWg5E4C8uS46ohuyem7yhUxwXesR/VHgs4pQdHgxIdQMnu4jHEg4YKBCWXFtuJEwNV+osZs9T2to
PadpXurNfY3PT9xvcxP/n8J3IY3KZSL3SxeAZ9m1a0Gu/OgSA17pmRXPp3/pDjOvaTb8BmTnuqQa
KPmQAKlC80N8b9cvP+z8IhqmR0uKZVHk32BOxlnWWCIhn3lENrIp1irZKM+RUynb6o7X66kR5GEn
r3h2LdhWVEL9LxY51oUo8DHaQNyUlDnMcibgi+0TW3iRngZyI6M68fJpelrYjbbZCc8g1rvodTUt
CjICzSoBYHewJGrWr13cI+T3OkQrh9+BxhRB11tSI3B173erA/nAatjWOs09ZGc/fPs7WSx/uCgT
ZwiOfEz1gMyyxGUDzxn62OhJ47rXU0hIE84rg2jSZUJsDTDgcYchWK/t3IIgWoU/nH8/4v8wDLrD
egZe+u3P1ZkvUhArG1QSDufedAn14damgS3TiRiIYaO0SgFX+Tqd2RUiXOODvaNT9s+9GD0KgWAn
lJ4XzRjtLNeEKAL5KfqSdjaQxKDe9OPvBXGVlo5yVdnN376EC0CRwIKhZv4Rl+Psg1QXztOXK2bH
2fW3u8a1riNt+VPKJ2VKAEEzUHmFmchTWEHdGoNE90om+ET5Itflb4tN2jvVKymcMau2dI0xnZaH
8h3YcAf8SYkX4EO/UaCIFToJHCM8d76UPwPkYR61gktGBSI1fM4FwPz4IbvoDhLl8Kew6fwe18IE
SwDpvg/YttqNua93o4nYLYhA9cjwpAvA3HPC2Dn2oS6XRUQafkNUTUNAzWcOugRyV6w97h9ED/J8
YeZZWqXNJ0hI0SMqjnjBcWenOrTuxfHvaZso4OLHOuhBssOV3ByecTB2z/w4FaI2LPNGX67GUswS
v0MTIqrxRqplaunnwgeFadnEmdoaqaCGVrzV4yf15TTu8zpEwoxeECT+nG17jz0eQAVTnG4WKnXc
odhISgbiF8qhH1VFbjkGFlZaCz4jwiKRmfm8h4ZZ2nTZ5OkR/ALU8aJQaPqb3Aj/s1549fdHoVnD
V84qJfYwZ7IuxTUFUdG9/dOyTU/Qfrg9qkd7ZK+4zKf16F3AtlRhLZuNd+VilqYFVZj5FSnTzDz5
cKJs1HE5lh7m5G7LDRjR7Tt1miAA2KHeN3P+WVmqGNmelqUacW3xdt3M+oxSwwjhEeppamtq7DkO
/O+6gvSHM7nCre/FwAHEJNWf1S65uciUEmXTAf2fjGL2pJBinu+gWhsSv9cE8kfPMYFiCo8Ih4KV
64NZScq7q8cdldXhrhW4rwLcaR6Wl9uoT9X4UnqmHlzuMUt5aIrc2gIKayRBsjM+VehCL62IJHmT
FUTH1miXkvooY+RhAO1ZDZuxph/zxCZ3LiNTRGwqreuTIaFwE8ZtZwyA6PhTdcyhKTd5DSt5jqWT
7cd/y6WDFOYvrqvxIDVEWItePYtAmJtRBtRbwdLfW/MYEj3kpmmLq9TewsyYmRBqbtbwIRNioL/Y
r1+CUTbPi/JNvOQwbgtlHxOorqhWw85oV3kffrqaz2zXBeYB80sUzD9y3WPU5I2Wj4vOVKT93vyy
Elkc691V1tarcuLXjC65sDmWjm1klcXYpz8eBYtxGipt6BCZWfaJ6PhsQ7nNiz+gnlbdzz/6o6Df
+4rYzaBpuDOQ0QOd5nbgUTP/KwWsd1bKYWmVHuHEZByHnpy2Jm9fc/5BHPLrZs+M723o6fo8ZuxR
/lSIvVpBYK+z/audKI1oxHHlwh6Jy5QClKvEVnZW5sjMT9KrKLfAOW+aPlZGLi6WIftVOOwFJuuC
m+twTPeJlKy1HQ0D3vZbE/P8dX2cNTmNR8dZnZ9m2WrMIqBIkz1Rt5Zk/UEIIv3V38hKyEqiEIHV
ia3IfjGlRtS7Mn/1x/zV254f8cnvSVDQFHhii6x2pf4UWKiFTaV6sPucV71isu3ownXm6Oowfvle
bMg2pmo4J2u2n7C6T466p+eJY7zwJ8qze/jbABrSNyDGmUh1yiiJrMXbhxmGbAGxVukvdyaMvAmg
jpfJj01o/TEZ/LMHz3yB+dOsSTsbNL74vIHc2BwNTa4sIsHJcPePHPVNn6n4b5s2NBe2GOVG/RxT
+jCNRmOIOD5v3A0S4rD/wSkoKsUszkm8kavsJEz2+N4VxHITwg20vriSxiEyRgZ3SAxBtof6Pn+T
rlIc4YP+nDfZbdHPoHa1KAzaNbUMvInUNcr7qYh4F9po6mkGAnmFzqyOc8FTU887LMibnpjgV6dS
iOCRcvvUQJ7rLkF31Ndb6vzUg245rIIkRK/VmFwpaNbU474IeZ+ymTOgi9traNGqov6smiil7545
A7lB9Ro6dsy5PdEpRvPyplKntsfhy6o4+neuCeuc0lx7dXA/aUj/a5lqFDuqM1vC8Hh/SvibLeoT
Wcmm3WozOLBvjgOQK2u6vKLpnHiHE8OI17NeaxwdYzGR1S7ps0vURRevFokcngrMnMsXuTNrROt9
dKme2GmyTmFyo7Z0yM6TxB8K22Pwsa4QU2NJBulTVQL8sS3qnFMjj4CqVB8tgy1ZQWc8cwaGxcB4
C+x2lSCgyYmBjEB1ofyPjGOkUf5hIMZVjKql0g6TJ1iT0Gv25XJ7R29qRo8rS4mpWCI1QNVL02bR
YQcja8XfRW/gtHyLtlvbDwLEiRTZID1rDd/7zvVfH0s0Imt32FBPHcJ+6gnxa6sI0R0KPu6hufwY
Sszjmu4x7mAeXonwyfLl58Yn+LF7n/R8B3hVA8ke3ol5asV/jjrZEamw9HF8iEsOG6+WNkQHCmkI
pvedAj1At6DvbY6Jj1yffjCM6T21ToflbA/K6USxzUSp3Nj44BRDMptdZDHTvHyO/rZxDe9rO1oF
Ybuitfl3QzWKIP4aHkMJ/Sjy15KRt4JUmO8qFBcXtGC9ekzGWDoKRqdx7CCZJ8vfb1Kegtn4oZxp
2q9QOULXhGhntHvjKWiMrP7ApQQnuif/kPaVGtX3q/4PEvP2RFThFgTLnOrmbyua6sc+ptKF5mXE
6Tph/RWmkx2urm5BV5Tvn6ADdmJbY2VvM3YdhRJjNKz8FeK4M1xOp36s0Xkmxezle7We7GVTJ/k1
XPDk5XFMGE6AZYrSQXKE7fwfoElxrZSZqebexvXSLnpiMQqkmT5tRPM5sizl2aTzg/1ClJE4Pb7p
9pey6Mu0WYBZZntIuogiA83pQWN+2fitTLHdXuzBtlg4lMgygs5rRn4S+lk3urx/cI5Woxc+Tr+V
kQ6o1LM5jJELiwPALC20mUCyVe7nnqRcGU3axap4pNgKkAWfqKceHPkPROTcaUAU/+CP3dkAM/we
13iWNwtXl3/RZ5VBKuEuX0JxeN2SWeE6d8M/kL/RMeWEpIx9blmyrntAlXh4o7VRMHBM0214CbxR
jzq69rUldW+VLn1mxtWJNUAUKyxT8jqAaL0ba5ZIW2DffRa7DJ4pYGLK8eI2MVeDrig2ONVQHcgB
H5736E4RP/0XvhNTMF6v/l2lIgWUebrOqbhKqHlL1D92XfZ0IPtlyVVB8NV3BFViuT6Y+ZBz2y9Z
bUnV5xiPkZPC2IG8hRvG7DKZY9Zvfz/+S7Vpe3lkD8Fxa7BlHwtzffoPlew/Y/2BPZd9R8rYlOcx
A/eVw6kdo6YTE2mXlsyvysWHEiK13P54OnjrR+cQrYOmypj391Rxrb+cnHOmuHUjSG8sQNIjhTd0
/CyXUyJ1KbmtUsdfdzbvpiSsesxuWymXaaeaW0V3Cyhfvz2NT+VfO05NPY+NT5LT38tiP7hwNETl
uz7BY+us14kpjHEgUDTWD7uw27B2/Td60bAbHGBSKTiLFiIFG2rILFRs+TLsnfqMb7eNvHHGNsy1
LX8hp5kI/uJx5Xh17Y0hZXSkpXok01UVdQRshgQZj8AKicVpGt4G9Zkk94ZEfF+I8IN+JOfoDjU8
PNWQ+0pnr0Boyd1hrHqrQ73p1adcowlC0Cfq3WjVezC5dPDwZCYJHBv+l70bWXZHoelylo7eXQcS
qFoQ44YfR2QLa1kKOuneYfWi2/zVYhfQ/uNH9hF2mtiL/Ph8Icvm5eMUrylDmfkLeYAFGpV/gowW
/0kfjKrkq5DMIGQMLaaWunpPPpCD49AkWVDjbhBvjvlfEmbdUfiQkp5Oo+oYs47WukG0fqyq63f8
Pao9YaDBe5v69MDKeIIze4irr6mipmA3nhSrdrwop9GnuNwS4pRIWDXrL7IGMHkY7d2HFlz2nZTW
Z2MquwJ9ax44OX0N4sffIHJIqNzYCSM5fF+GGG5/1U1aFbzJvlCi4Lkd9t11RxdeJ4s2msDN28Ea
aifwD7XxhkJD8ReGYdA3hLYeKPGU9wfo08JKpnXecsHqehohOTsZ3TKrmWHnJGLZlf43AjlX/1Vi
R39E5PTk5nK3XnASs4sezHnn0IvThJXCMR99ieYplJ9zE48o51YKP1pFCLC44eEp0cAjv/2IOIHu
KS3XA24HeD+Aolpul3gLq5kGgdhPlA51AyXAbepun8c+w3zxgbgqMK0RF3uE2IDJ7cjHsVcYPdYM
2WvjOyX7aI6N98cL42Jt5R7Hn4bwJpy0AkPQA5ZnSTmY8y3lKhwQJew6nCkgujq+xG4S98Ak+QgQ
KTAlBuPAfiTe7j21Me/UTvWAZL2RTperH+ul2TfTHGXGre9D5fGLGfrUf7lVZpLyZinr4qvwJSqD
teYcZhrcTAnlLzqpaLjbmwHSjDUcPaGx3GXQTMCWCWLw+Bcp1TOScVTKuZSLifiDKXvrMqo/LPHG
Fn5o5JfeoUsd56qEr4TSh/DJkFPcsM85yznz5MyyPZINq+LxP7XP6ebEudoKBEx1IfgPSpvIFpoK
1FB7ozskWEbq//ZiEcFL1WMw8PfyicAedy33aR3UUQPAwdmvOTE4pz99aDBWLdiouW7YCFTV4aYu
sC3SSAykQySK7bwXt8NH4F+D1M+17d0pHUu/Jm53rkII/V0GI4nC0bAFc2ZBc/2wIOKSCaOq5yrR
Hwkpr4i8htwHkP8uMBCLVmOr2PudB1itGKU1FVkAXEJ9JBjUSIJ5nv0gT0ENxaFks+4lfeC2i9YZ
bPh6wskTS83J1IqFaJ+TdlHsgInBz9UVxXomUHRMPzmbh8DMwhLf2HoQcY/wm7uJcwt95UHhY+HG
Ck6hpbEV+T2rBNGWi+MVJnTXNYmujqThWT0E+qt4TRCqHGYesDlx/eYxgUbgLX7evEVWfcTP9ivo
Bxf1SQBFMeooTpgAN+bYh5opDVIuYz9KV73y1UMFFWoD2s3MymVGXwA93Gh8fKLDI5s6esFBN0mL
5PM4PxapWwi6guc0jqYfSrI/CZyQXk83jsjNsedI6rZrtX2i0iSsqIOIn58sTrVNAhCOYJZ+c7TZ
bJZGQwvajzpzXRYV8IDvVqR0AwzZX6FaQi87OZSSVfrBSCR+xFDVwCl6NNdw27RGTJ/qShx45B0S
ch8NKp54Hx8fVE5WKicXpe7xZ9ELfZdhsit47XZq44Q1akQC8OKfMi9sGx5raJOCOtzfdxI5nKVa
mu+NWScVSmEnQVxYNhYGVoQPhslXLbdtTw9TLsINIx7qLqJo6xL88aipd1WXw4MWsAPYcrW/iR6h
hasPYQKsXL8EtcsGFv2QFJFdPtteU/hayTyFC7ZC1jlvbyM3+bwvzZ9entHOcJlmcNuBNV6P12/0
t8VHU7JrFhmpsm5h6vGbjFANQGHaGV9AWBu18Cv1yRfssYg0cnUOVa9oYLlHqa9KLUvKhb8r3r2A
f5IJJXPxDxcQjXnVlKHsGS+9E3h3L+DVd8b5VddilTofpcl08SyPErpdV8ccJ1AKQRh8bPGdZnGW
aLS52zhsWRNu0U98MPkmzvbzozvqyRqAA78VblrFbuJBHkDIMZsV03IwGirkQx48TJmukgzddvCS
3huElGc4X165t6bfvh2C8PonPoS5MHZKVyoXf8USGGFYd9MvurLXa3552a1dbDNx4A4mjWSDh5Ks
jPstIJAGRsUnSPZ7GZ4w+84cDEyc1Zh0/ekK3W9kaDobYZLXjFJPwnIR/YOX/MwQI7PgGAxQCs+r
OmDjXE1fvf+txLi0cNAf7GlvDtIheNVUzKLhE+KxZF+vYSjYdG8qedjlSPBaA5Rij6jpy/LJHcTi
xhLV/Hzs66a2jJHhkzX1C5OXAmbxB+j2MHhFXUOFseY+GJSWINvydVbMib/Ytm7bdCVtX23BTLSH
W5XoLhF2owoB4FrpWawyCzubcAK8hRqlhm0Sb96MzdTyRTL7cAsm+ka8kDV50B0mZZ93oAbmi/fm
1ygJ5vS1m49U0YVD10wnpqLF3XL/sihdPM4k65ZCItEwDp4vQq4/rmeJTA23DE4Fv4Oepux6fdNG
96b1OWgiRvnnQjld28Fj79vZdn/odJImpTV2R2rlYNIz2CfEn4qw0dqTSs5aJTOUwTyrBZOPq50W
WcqOPaYxp0N0uQ/q317qePRgdFnCsacoT6MGtDsMPB/fDPuYRyRuUQJt/wBqKqL13lCMzUTWna7g
R4Ggl5DMhvIXt8EpnfF3SuI61xXIVEhWSmxaQfDXChzabYEmA/ioYlNb0cLGz46GE6oKQ6zIKSj5
Ho6jT6iPErUGYKLolyF0HMMgwg2n6EFD3McOOwbXmqzh6EzKyjrmCLHl4s8xRnxWDMKKmXcjFUrc
zE4NK6xEJuKin90j7oWCyAJmMX7Wp9WR/f9H7d0HbgsX4S9PoU0kcXYfni81yhAtPT/5AOVdQx8b
C6FNFVCKmZxk0yEAGEjrccF9paq5Sgcb6v3Z/FxTkB1ks8GmvQclr4D+n3AnZkXGh/Vb8LaKh7VN
MS8u+R5WeOUnMEhISqbj3ta6qo2RkFEezSqkYcGpIzk7JTxQrPF8yUIujxuKcDfYN+aLI0Y9dz6Q
RgVuK9AH4MFQfOsSGvQGvJsqtlU6Tqnzc6FYRfw556/XA6n8X0x/Kqkbro4HoZI1OE7yZtS0UNhd
mDWKRyTAmDF11q4n+MXKzK4DRLL6CSroN8tzR9kc0HuaO2I2Y0faXo7biyNCxDqB3i4Fb84yRB5b
bnjjNGrIWubEwEU72NiQifSamcz8ugfBNohQGd3MDwzhvc88B13kuTd7j/3Jd0gsvLwWRa0kdAID
DfKkRHx7Oespx2CG8i0zqbHr8rOsgTdDYw3SFBOeMn5zHawjMljnhC0DAHWceJiLV/IX5xE+AsB8
1z7VHjtwn8IaBVMFc42serBO4Zk2rHomRpZpRO71sKYJb5hA7WYbk0ZTb2xHPaTGFBnXF6pbgTBz
dMYYoiy4XVe1bFU6NUvY9+5vRzJN2mmjbCC59qFVTJJxgA9Ebiw+QzpW0Z3YTGqypb4O+tFenwkO
WHSTWO+2iqLyRwMuXVBRTY7meBg71PrTrxwUH1SvAV/impK9mg6KkHicrbq1jSs6V4gxaJkdJGhH
jlWZUV1B2J+eILetTXn1URnhEcgfcI3+n6uBXN4un/93+jWfJ0m7Ru+GpCGP8YQHv2KpYsSwX39k
bD50f07+ppBLPgG1ZhaSmH8XRexCqOItugWD+ZSNFHZEn/mAe7XRIlWGRunco9ndfQXCT6KQiSQj
VYzO19YhOHJOi2ZSxVRb/T+uEHKoAsVyOdGwulxm03Ab0MKbzeE7oWcX9DBZ0QjSrnYZCo9KRU+Y
UvkEXpGcX7Hx/ieBxqhiy4LWacOM08q6aJSB8AgXgV0ylldwMpX9OjZup+fe+psrqz4OmaoBQnTH
H6eKvbIHe1EnWmwGefCj9tEvLjBRX9U7PsWAP01Fo91M1wPiUMCB0zUBKmumpEW4o1RPecH4oVPi
mW+03fFlCKReTqcasLIwY+FLxIf6Oh0bR0QzX21xCpLy4242U1cOhDmWOKnMPNjKwgCNTPqcqKhE
XiKozmgYRopQCaI5LUkSQikGDh5QLoLUyjqWTM5b8SCa42VFZyHRLPD/6hq4lU8gHBYKNFlKlbeo
lgcn18qq/l/7DFYNAD2PdHLdMSMeFdT8exUpYWQXRvvSUWjMpTL+x83iXWs5mauAtGwHCDpqkDcp
e+J3dbUJtaXvxrAQiTIIhm+O7NDNiZfvb5ckUFmvTMQvX3dBVjdHHbJibrdDWhcRSx1EXB2Jt88k
AkbY+rSamEjfw38l75UFeHQ7sgT1Wha7iDxLKnW5/VNUHvIpQSQIh9BypSf03xI98rOZpjrAc0/C
gidINn7WdRagED2wNSPjQ1ysbe1oU1R+PnlPEnyLSUeDvemlktkY7oU27CF9nCunn1/qdq0m7o/m
YR40oQMLuUa4epyqwpJWgDLSkJeQrY+wn2l0NW6qDPkRu6jjTCS+gx3kw0I2lADQdIaKbdMstcPi
4v8AXrjzr3YaBo2glhBIDVIq6b517vkrPppwnqlCoiQHLQMmHszYFn7bY+DoooUN5HEsIP87k45c
Gnk+A23VtiX3VPlB/1cjPGU743O782CNO7nS/ZCx9ZsXyERSFbOw7bjTwurrUz2E5ZA2OUERgl7I
AB87YNamIs5nALngAeUeu1wf1DOKaUC1T4tiz1g+t8/aPHONutNqg1w2wuznK04UQ3AF0rlWIL4B
dxEWmaWVopWIfOuoMYxrn1Yy/bF4rsgHqPtJEWQfHwqs4OYi7CmR4c2AKqzKEBfj6LXUTlyf7iWR
TQ3j9Utd0PoaWoUIzcreVLvz9sgtsIR9sDsm96krGYVYFERbxB9ymQZ3Iz7gAoTF+O169zmuKghD
/MzUJQZ6t2msFz53oiBEq2XoSA/Ut5jDdukKRx3CHtEMyMK3LiITq8jsF6TEpaYyP0qJq5O275Yr
ftX0TpjoQ8S2TuBVrFmC/YnBx87VbkAOyCP0P6NHmVYRysg94Y3BtOAysoionnJMwy5HxGfSg9j9
6yoCz7SIVUIjRLX4KGu2aIkw7F6Fhdb+kS3tMdVMiBs1kkhM5OOHHxq/ioXCUHRc3RXgZRMQcX51
aadg+1EXCxyCu80nplnk1dpuisvntLJMVTQkd0+EbJywtOoL8pq1F+7EhYpynZQVJ0OwR2Bz7JFk
l391SbMUpZx5ozcvo7VcN6rzXOcpNeln80/WjMLs8Pnegu7btG1biSq06o1z7dXAIFQix8QD0Vun
pYz8LafLLYzxvftz5ouQ/+ep57Ilbp7jG+BxQ/VJAxVk9rmRCCoaIZZrOPqG7bxrbwQEQ0+h9C2c
p9+MwShGWJBPKZPfWU+TkcAsK1l1PHRfCM22GV2XaxBny7IGrR3dWmYa5fcgyi+Xf0TIFXwRLn0J
sRmsjmRN239IbDtgnBIW5n18RmFFWnhkzaORDIOgaAqcHyRY9WjQ0asY01Ikr6Akuw+ZYiKz88mU
ypJ9L7vvVj4c23EWTZA48+XAVVnnWQr1KRxJJGN25Ls6tgwJ/L8QAgxTodUaACuVmKCbISmGFl7M
+fk3G2tEKVb+WfgZV5JoW6HZvONDAxWfTVpiVOU38EVi3WUVy+zY3XgiHwc9Btcl++XVFRhoJuUx
+SWJiSm8xi4kdOyUKF/Xd9eiV6v9WZp+7NKmBRXbALxoFBHsvUbCIxqi9GmA8x6x2HtKvc+YDJ0G
F8HrFWSlSrwYIA3NIBGFQ2TaBpjCS1GJe7ogu+R/Eon0qKVhVvW7a91sDkpWA4HQSi50I65Q5xdc
FDXl8cVCki+AJKJpNqJr8LosMSNC7BMZ5PAFX8jRcbiC4EV+BpOMkXcGpX3+13hrphrwaRbGMD8X
v7aXCKy1eHX7LKKtg+DulKFnCUJO38lcaoP+EJEaTqQU2efk0nANWPEPFJ8Ym4YXybPIETlrSlf6
BdHNyv3ncZSktuy7drrIF3Iip1VEc74upiE24wnqg9zjAN4OUDRog+lC/w27F5TSW1k0vNPVt5SQ
auZz6SLMuiTYNytskwDGyX/7YiFw5ZenrsjchF6sATyEdnzc/OKW+SxjG3wsyXmREgrFQV2eDSKm
gYjc9xYnVbGZ2R7jkvwme2l7c4IOhI+1ggegLFJrwT2X+sCWIYQV3+Zuagc8mhHTuiT0GJsrryZ2
46U0zjSSm0zq0FLoJQ3HfyV3dYdBQPEbc6XZGOS2HzvnGDNYdPX4Y4Kk+DINip/URd5MVreg8XpT
btoClcfIWTXiUBhZcDsFE/+mOmUyXX5CQZDNdJOr8y3StzAKXN9M7HIx1H6SZj8C27kUL2QyJ20U
f5gryUb6iRn/1+QC6dI3OI2RVNhHp3qwn8HggTD3ac73hbKi+wogEvDC3XluOTTKyX3NnDhBbCY2
SURkWi3N/Lba4XA495I9DvECZ11i46Whp/pX+CEcQFw6xbv9uaEcatLkbsWnQq6k5Adk/nE2L/vE
zdQh8OByojqdbM+n95TWHI0CUjI9rU1zjA+8qpWyWarFk9DDzQZihB3wdpjysxk9Sj3JIRYi6tXP
PEYy1a/4FkbfdUtWj8PiFYZnLP7IX9rimVoBOn4tE8sDWjt1nX9YEP4S2r3/VsZbCvq3ZDWF7IDa
CEWrxRqV6MksyfAxKZncpCYS1T2FcF49XnU94pg6dfMTeP5viOn+9Lq+2zNsMqFRZwklkka79RJ/
/LZNb8Krp2kwSjgBHHvlx0yTQCVGnHdo6wwXrGr4T7dhA/6O4teMTC/PzBF9EBgt89yL92qe+5KD
X0QoRX5i/cr0rmHqmc9NKRPZUlhH2kuuKcsh+lSvjbE1+D6+WlfmFc+1Bn83azy5DQCZUaWDSjST
cBE8yM1K4vqdz47Xs2TDMrRH1X9jGfXxk1Jr5LlLgRzq+wsoCJZ/f9gQWBVAqrgaProT1Wr7DucM
Q9tXmJ4FpWRgsAWIzp4G3WiNDMaZLJK+oHQNRcD9kZZK1HKWLSo1r8Yzmt51h3FPqB6gjLky39J2
s8Ppce5UiUpgTFTXeQXRjR8PW4OgJYgamx0B+NynqCfehIKF3D9oNBmKJQcEEyavNftvnHGeFr3l
wdo17B5Wjrz/E6xku6lD5WB7PYPI6SWjjkN3iJaQk8/775WZAQtafps15axwdQqOim2fsn25+B90
AUR/+6nONeUkXl7eD+Hffv/ToIBkI66NPDCWLjhHV13yA/qJ+a/Hb7Ep7/fA7WetOjNEIT2x8dIh
Jb1JsP26vqvniT/Um+dEzyuFbpc2F4k0sFzk9RaFNfI6vLmLhGp5cjjcY3xP1kVJSofNIonOlGmP
xsdJxMlgB9lmk5/0z3JsIWTwZmbOhHyeB+w18D8V70rCzzWiEjg7SKfxtBQOeWKdv9pg6l4lLWlM
nX+wi283pDcEpBULM7mIcX8oxbSq5jQN+3EdcWDxKMVDPspbkMOL2SAl6YPP7VkMqaqsFOG/2zyw
BIv6lfNfUPIbbtucA9fIa7l8eSDIVgpiQq0CxkcxhML7SlHlcfXdArTw3fYCjXTS/rXtyTAPqAyZ
kXqSXrb/Tciu8eDEhDyWdqz3MdscuyH9UmMTD8sa5zRHchbTBIkF8vmatwM0roXldxLj4aUIqtlw
s64qAt3NSw9xtHhWPlT7bmVaa5tij21Pj4Vssc6BDuPQwlKoMt7L1L8d2+TzKrfxLBFczHvetkhD
Pk5W2Zic+ZKgQobR03Fmq3YjW/YbBOuhMDsLupmLCuo61ITojwkBasO0srounblNiS2KZAN5PGWH
PIWgMZCUdxWNPVO0Z3P4pkqQZjj1w/B8UHl59hqbb01X45hkrX2OaCEljN0d8TPKgENclm1pndLI
cjR1G6u1RT2t8pHP4VH5mTXLiSA0OoXqRkjpOvz/3OanomQ+i50cX5H3+SQsRfb0pGb5em5ILSqv
oBwDQlEmj5+9+eV7ly8xvHUp93XMcmMeRykvFuWsdBnnT0CxZ4hf6+IQX6ojmfRszQ4r1+iiapzn
p7Bt5jMHvGiGKW/gvgu7cBv3ZwA8bBbVXRdSZqYnhtxfez6mptYdboYk62rYOpbYRFF4Z2BqFlbQ
6rXT9yNHBZeFM20sFfsIuQE+0QbfE42bqwnqWhFqFnDk9ATfjBmbj0jljUEE88CznU0GEsYF9Xo5
dyJ1+r6nK+Br7sgZImQ6+Z7USjWwqfC2fTiLnQfpAM/A+oJdQv5E4/RL/lCAcNGneF0D+Lzjqm/6
I1taJxh7pRDaiGoIF+EwX9B6mpr55rhhRyYpwxUAi4MlM0upuP6Y7rJr+cq5FA5rGjfZLVh9cjss
7TyeslBoTLPj9ohooKn0jBJau92ylou+/I02sxLGtvDYLFsqsgqVTuLP371v7CDPCKl7LLgZ4gm9
icmUBZ7z51Tq7SKCM0d6OF2avRGWQdg2PvBNQW5rRJINAdKVw5T24f4zENMEUPxI9sLhIi1ZbOWI
ixOVj2GCR/QeopVq40xzkPKEhojYMwFXlUyFlx7dTlvYgVsPbeA8Ii8uCvBm7f1wCtn1gTXZSd0p
xKuAiVhs7qtP5VU50SCjYlezQKZegz3PC0qmpJbEdtNe4XEafSvYiC+Ogn3X0mOb5L4H5YMPLBLe
LweQCEFOj4SXSahd/9wKhK98fDXXVjQyR98vyiYl7UIXEPUf08BdYTQqTBCYjxT5pTQ2+i+tvH8/
2es4ZgidOGrlZktwlBRVbVza0QJ/t7Fby44LRmLN/QPNlplVPpMpCR2hdMBWPSySYvOlbdCkGZMm
LETmITM4AjhHq3/LBp5dUujsTUTLxcrH/0YlQHV6z/xlQ71iHMi9LXLR0kfkAnfPbOvc3mxH1n/6
Bsk36rDWJwELdEPURdzPNd7gX0N+/UI4qwrdAtKhymWkFF8WW75d9kly8Rag0YY5DRsI+E3aUO1j
4jGhsJarV64BJMCAmBhI7Q8tilfNgnsxQqJfRkNm43yFYdrv5nT5vhEXr4iYyqWR+mzDV1umwsNM
sO1Y/aaVAsV1obcuW+rTTcMcJ+xE6cQ8e6CXfKF0Y5rchFN2dbzf1GbP7vjZHl5AmYuAgza4KDM8
sQJfDI22GjqarkTUHTgEglVcp5cIUthgNlxMWh7aSE5zGMlkJjZVT8rUWzSM321QIRVr49ACk+Kb
+CItzjznUG+rKtoOciVyfqokL8pxILxowq9kL5+sLlO2jQNHImg9C+Z2OkyEmnEvRaTuyolvj4Hy
Yzdo2+FBJ7mXG+oXN3tBR0RogCY/lgqmi2dzVR0gmuqU+BsvmsdY6nLg19QYb47jBKRJmaHp10Lt
u1YQLr+tlf8CkXXDA7Kkq1cqPhQdLc9F8IDbOFvoVrYb8zQs6TBUINZ7Jl2Syant3SVhpQ+u1Ga3
12+YK6S7dnHKpHEY6SJfepTV7d79rSChPRnOxIXkiGodeNN5eHGaUEqw5kc+f/RSYLWtOyi8IJHP
rOE+t+dktQttOO9lVUT9O2/tfPWXCCzZrRUtOb8UX2LBBwRzUeR+fOLxwg8sQqVAklUZkiMJuz8n
NXZbJoLKjwVtI/Wvu6p6s5bAjvR8efLDh5oitz93Zr5iOFLNj+eS1xz+qDBWRX7t51kwyEb4c/dS
65Vd+9ZeA+tU3zF+cvcOqEuoioUAXyb4s0/lLBb1cqIhdqwlsf35eYmttl9yDMgLaGMNDvVKMIhR
ndMMPo/emSo1zwFiVSpZKg/BGPUivSxQVJ5ilQfS1K16RjYRLj9wymBlL1gtY3+nsv/ExyrfB5N5
/fVtTt7joVpculUuBRNmJYbZSbb/06aDBTFkqdQx0MwvkRvQljoWDF6aQM4fKee0Z0RK/bQQyj2W
ZJ5rv8dN6U3PofPYHLuMSqDcQFgcexskmx77jw4FdINTRSRBvMcufObo+Av3K8UnvI63ZNk/xo9Y
WiybSDYfFCslmKwUcYi503l9B2j6dEVRn/EAx6lPkY7nGsLW6AbEh5rsl9x97O48IZ9yLh3eXAJQ
otomWCJRMp9hS/GDnNv1LFDYjWuNHYDPQKY8xtlJd3V4egZPEanpNC/3BqA1UmpHM0zr+LQ1V0wL
K2nw4BWvkRPvN9sNImKL/gKR0WWlvFKQs3B62l9YOOhISVGu/tgPklGAjiX3ZunNJPv8AVtYI348
PZWCQoymDaQh31kn19RX9b6rwzUfdoyt3ZMlrEyPlm/scH46+v3qyj4oVtOxdLU3LjB8I2JJss6F
XpVVEUK8mmKprqDIn7yl5d3pWvDa7r0nfbq4Wlj3bffwc3Zpx74eC39ncdCUVle+Yvffs1oEv9N1
YZtU/huCqED25M/BRNo8uM39qTgWQy78Zk6NXRjXJnxFKTJ2MD5TUXkNsnWdB07356taa/NsRAe0
RLv0qhsxTEFjOjDPS90WnKpPBgu2pShX9jrqNhAAsk8o3U5sJxdDucwp8Rd10iRa8By+JfRgFmyR
0FWrpob+vGgB+jxv1r6AUFzd4dybbkXqx7uliE5NALwcA5wyJJgVFi1wB6gsHsLiWoYzlq8nD8Vv
7no3CwNImVFVju0OfKbOOqcZqTqZUXbikqq0WgPxEByqmdhd8r2+Y2Asrq0IdYrL9c3j78fLqgph
8i6/6lz62SnGudbgnraJfT/c9rss3HP3HIEYyXRu8WewZl85t3Pi+q8JPwZw7q+rPBj0J4Bp1flz
lgmQxNIIMLp8v+y4vuQxR/w3GZLM0AxOXZZvAgZHSdjGzsVNv1RW3KbGR4vF1Ohl/sg8uD3KT8si
+LUAJMfkQula/1MpwuzXEJrYxk1hxx0Q3UDg0llb4QO0LVkmpHWZXFPXfsPOEp7byTKrVDU5O96w
jFhN6WFkuziWFcBipjgqOLvEufHOVDJheXX/y3XEflGLc8SENr2bSz6iGBmfCNjoZ2qoxUgASKkT
EY28+Tl9aop4creMPJncNQRtU6wKkxdsLzmBprb4wKcknw+pnMuctgpHKC/R+9LUO0fZhBN1aoG/
oJQ7JCm5iAhvNKziFGG5XMz0ahTpLOZhMH397p5pOMRLemiSAYb3fUZ6MUeopIKDKbMH61TiEZQ3
t0Ek4jQdDPLHxkLSjkIwYU23swRcXHX8xlkNqNE6DxdXBi9YeDKZ7i2erkKRrRFBY38U7edBm/0g
P77ZCCPHqy7W5WNbNjKmacZ1x5ZcFB9oSeiaRjSx9IfJgp5Ng/K6/A1v2NXJR7f0AYFLVqUpKlPd
bjXFyPfLUF9Wj2RsSS1Z2HaxkyPfglHnV6/obCJZtUlAPbxhxKwrR6vNR3jmG53o/GFwtHZ67WiI
67NCDWVFdsGTdVFKVrBceXmBLJh96aib0vyGJ+doFoPcICjxgTExNMyVx2TavqfEK8kpb9fmrYiB
lKukqmUt6zVn5qQrQTdq9E+GeWIjvVthw5I0h21kzP70wHAI28XFV+NTqg/S9vpVGSYvNv0qk5B+
PreeooePZECs8GZEVzlWpM8O7URvfon4iGVoc2dX8gU8vcMAjJ6WIjRXBg0ffndV57XzRxeExoHD
/BTKKfMksqiNLd1l875tPc7VdJUgKVGMLzOH4Vvs4nPeHVQlsHVks9upb3ZFR2TyaCikXFKiXg4m
YhwYTfM0BZWl/lmZYt6f/AT2TYPuldXloMem9j1UHmJlkxs5mFlIFRWBgW8BWU/RglnxaiTT1B05
oAn24v2NDz1AeM3UtetT9POe1c+CXZXViRWqU+/TdT13SlOxPMn7+gTTWOHwUSN+i8DA4EE5v++O
J2EBF4mVJwKWuiJFAPS5DshJ+zsX0dz0eOsN7mnsfrtzk1iAZZfB4JKpXLo5hHx0RVKmDEy7jQkY
CHeiWncMfRItBg6M601H9vYyJJJnohwbNPCy/MLTMC/gA4XPk1jzRVDSOaqHCwM0pXT6JcQxu030
Vdt196uicUQlbHdf8smAsD+TvMT4g40k7FZKcli41fXIkQGkTymPoGlwl7oROTyO4ecVxrWDmXgp
SfSuF1g05Be4ct2RI/q/2WqFzmjxnmAAP5AeAGUjeCzEvS7mvyVPgBWP4dF7pcU4M122S1Bw8mIW
hNkS6/+jYorEfoCkWP4JUZCXAHPfqOgOP4UqRGpDHf5TfB2/TeMOTfGcwI/oomor7xQC/+pxdqOD
ylVlB7zcSGwTdR7+fumfKW2JVCfz9Ng0fksJgGukuVHGsaFQrDzRyL9ziT179hSebJIJJjZZhLyJ
WR/2tL5EgRYxhKbeYCBFXAfdLdM9opAuhXdJ1bNk8gh+gpnPkqsr08doN9XPY6IG4yzaODcKKTz9
M/N/bh9JCrYgDxb/dRx9UQ1KlCfgWUeZgi49HpP2XhFgvbx4xVik7to4uh8h62NMuTnCV2ddfaJy
RAoTDFvJ/6FDgNc+HI1o9W8etqD5wZxsI2LAZVTfZtRUjF+3+ykvBWPHUP1RGsoQ2iHHZgX4bSPu
hlrgsa6fjkM17WAj2KOBbQlIeult+8p1va4ll7G+qKnf+iK4kFYaBaBhKRhnwqqmHent+EUm6byW
5f7xtTTKgMdVe2YURkIdUI1UfsYCukKgsSPPtLlZ7gNZ/iYSpy2IVf5OUuhicTJCNwNEtsHgSZFT
W3HFzBmxVg7vi4aoiX9eYiab/xxt6tFr51pQnt8vgQC7EUvdafSgWUWt1MVUzyL3EnREKzWM7v7V
1h89TKvXkWu/jleyrhE6Qx5uFZ9BSAlePJRFHVdSDZS/K1lHU+zzdUnpBiQ/PO5+i+ywt2beusx/
GbXw7H5WBtfTqs8t84JXipigD5pohG4CIxbd9YMhVimNblDNm2dmc6z0j1d90qlbYgPtu/SLUhbx
I7fvLRmQH+uZmQiGxXQnOxXLqc6I2UrBCq7HuXNUbL0oBwgBYHauJSRF4qsBD5CsC9STbGGoJa6X
Aw/aNGXyitdRe5GHklhF9cb+VtY5gf2/yciLaVIDGh9z6jrs1nR0lsQHgon91ipCYlnjaU742z87
tsu7JY5D0s2I/VwSWOCLkNZDmenEOmWNqGBvlQ59dNYL/77Aaeyx6swyGhRH63xM9/p3wP6oZMrY
3U2lwjUgLcQ/lkE/thvH8t6T2vKvmONFH8Gq83/A+fwVQkwTWA4L4HRST/vH4X2GOHC9hFykalNG
5i8q0MfvoA42oCuG7+hlKFfQybB2vTd6itbYSD1CLKbHAa3ZZRTQ0pndrpNue1mQJ3XC0ptQL+J1
jRSp1MUqn2Ebnuu5NZCJwAZ3pZ8AYUnXx/Seei5kKxKuVG8MzEWShh0W0qd7LEmrcF+3hM6PH2ba
THuiH6ETrSSU6lecoNWhqG5+UpMoMGVOZC/HsE4/R0Q3OaYIrgJQ6JdWmxP8PT3LsYTLhXCpALoa
9kS9YtUKLI8BYOxdeC2JVMBAb5wvx5YboQSs+MHCSoYnBpHsdSEycL72AB80oZtSA5AK2CiwWyep
uv2/dilxy8pbYPSAvixbNG59HFF7ww+pw36gIA7izotOev5OC5NgI4xjLim7/JEMBpit+1f1gm1T
x9ceg8HysPCf7NCU/43ZYDHxxb72RspE1lrSpTNjlw/nyDQ1iYoyGsw8WIiY8Tzfqc0Jl64ZWX4v
1R/0vIfAIpoa5AKXIKFRUauroHkPIxT9x/EASCYLAOY0O/pAt3NSPc+YvwFt7YY2Ko9h7NYMh+fl
gleJ/iRxHNYCm2uqT6cqnDNpr1lNhNwr2pfMPVVNhnmwVMtQ3+JR2gE02E16KvpPlyEhy9ymCuBb
VnHDJekqV9/t1BNmjDJ2E5O3i7JGWTNU9LnAvra/wEr5a9mwNBXHxRS7h94ohJ4zwdoAeMk37KJ0
IfhMzEDERPexUzupymvyv3sLFezI8NGDmmp0RUoH5DWS9fnEiYGGC+BIRTh/QvCguyqTr4wRVT+u
x8kYxC5MN9bHCR/7FIElFrAJcEtgaJQFIrVLEu0iOWyH8Vy9L61fwqYS1VlAENaFM/hWQGyIX0eW
fFCSl4xF0ZOXIOru6ZuyVS1AV4cPH1xC6+DzAwyeqb0Jazm6L9VmT0T0D+c279xABMGSmnxztud5
vx7cev65+FNRQ3ulpSJGZkuwfF3q8m1EU29PMxqs28Pjg7h5kTs1wWccpKahmdBDS6+y67GpT8Yy
2KeI6tXawDFxICGZMmXLMTwdM2VV76dSX083+g9KqmeyGePPpMGKxIV/eHTumHP4vEqX4BB7g0iS
sGXZGYwRh0c9uz2xCSWsCBvsvlvGeesrPkNW9V02rZzw50yiqgqlQyKgxrLSkaw3EjgEYC7206Lb
k5q87ufNOQdFBx96Bs3Q2r7ygh30GZ2sWJoiC4a6m4vQPD599+ks+rlsJ/yPl3dgrogDiJ2G9eS0
wSeZMIggvl7XmXAEJoNJQHmkj/9ezztdkRUZzcqph4btmMyIYQlXVaOpXyuVL8zVDiZscJFuzYDf
GlvSGNHWK6zp2u3EhYSRGfUSKaoahrLl2FgUvHYZ51gUpVBEeB9wMX6GRi3jC7fNVUXRCDsQp47M
ULjxWWW1jTQyiCEFaazdM4/fILu6+Y0A52Fg2FBCjgIdjxjbUk4haEE/1pXQmeems9Sk96oLTlrK
S+SQKafa00cAtdOAVnh3iFFoS2ewLUhl2s454rY/TSz3qDYm3bJRmp5VbZ3iZ17GYN04jyVhsC9j
siU8pITxQlL/0C0CJNJUu4vuL+cep0z/ve+VMTZ+QsASf5ZikcaXAs/Pn3njWrJL9CTNJ1LYVOui
xxiT76FefxR/wgqyVfCjYcsyoWTCySFflc0zxHajgnNxZ6ACGZ4PQMnEUuifNeMeN+3mLHSgAw5q
ylRr0SIlNdY7LqL4FA7bAFJrSgCjRftVG6CGxMMtpBzZwzajsJgESqLYrJTbHezAhsLqV6FCT5S9
1/M7J2SAOQx+lDJgZe6qd3LXntiFMAlF3dF0TaigPpumhKJu4sCsbkd5aoLxIFNfxJ8G8THfiHWJ
9+GcDK2tz/ApkhMSjwA+ZES9nGp5PHQexROj3juJTG1nx/Y4O52PBU1TIK7wR0SGOvd+qMCQUJFH
1c7Iobl/wa4knA+ZZB9NOqEmWh51KoqcP+pEYbBfk8f+PO33dyqR0pbOYmv0LGGGcVpRhGtJHGBm
xQOpfqpqKDk8XcHnnxpPgtkaTidBZCmZ4vHX/ZPHX5LSg0xj1RkyKC7MA0PYbYw6/wman603No/n
qJCqwf7/YUEUd+6oSPteoKnBOVYp/aQcVvclWWxTDjJ1g8moJHF9i/Ur1N+1tPk8LmjDzkoAtDZL
yqseBdxh3hqKiKC4xQDe2cebybI7tvpd2yMB0JjVblYpn4ZFZytbS0gaWiofjjV4+TpZy7wPl/OA
tuHwvtV4cwm8Hk6xs//ws6iTervqNULTlNrdaEBvbv738tzmtvqLkZlPfyF033tvOpK8L9qZx5gg
MWSwrCLSbC1nHMkJgMO1CQQ5QDASq79zWD8qwIEIGOpGFpQnY5yOgB04U1QKnAbumNZkzY1vIxLc
YFHamt4HMR4+OvocqkUagkCJ6thDKDWd3JLyYp84DB+ytlloKJSAOKVwoN3r6O45z2+Ph1s3uW4R
X8xcTU/TguE8k6V5kmvefrL/zd3ETrzwVG3g6ts/zihdO8k3vW8wt9tasGVVGGlU/RtPG1QCvjG7
PXzXtXyd926/YewnpW/wfbU/q6xh5NfpaUp1A1IGHpDMHIfPNYP11lXdYk/37JNHBKM0gLYagYHZ
hLMk7N+Ib1omjtPtqxEU6dj1qKosGJtA3V6dvR7o64ctjwGrUQ1U6jlsyWy7PPCgfKNEyyyWY6Nb
86Rm85MCyjVjV28a+io/8ap3p+wsK+d9yc7P/8ri5Wr3m3uNyihNyYSsCaJDOB8zeih2T2Z9Pi4k
fghpH+st/StJKObU3gAZ1fqzHocU3n5mJdDDmpYt5Hwg6GAMDzktM9BR5FcX02ZhV1HonPa91PJ4
NEpZb+S/QK9StA6J50+OM8AXweKJvHr7zSTkX7lkIh5oNpbWgmqCEN4U9RmTMTJ3PD5naqm7BcOy
sVLL4I2GxQJ94XKoCWQHWQtVg4plEWcEbXHx6A/mXk0W/15sbYfni2DUzXrSrN9iMrbjdsd9Mtrj
agLyRXdETzX7AnzfUYYTG3AXdvgitGJJZi9h6dsc2IZ685h4P/60PuUtVsgL+lzLvFYNJ+7r9Hv9
c1KO7jHqukMh9oZmgcM2LdrKvz+L3zb9IJZZ4/SSO71WxAoiFMjjgZwXPsJoyMHq1A9kJVlH5rbf
XGMTxgjbtZCMB/BZHtM+CHP76LBIGlb2W7RZkLbUdZMps6aOkmW3Qx9CQ4Ly09fTqwPRZYT6u2Hm
fhk1ysc9yfpnYC/iY47AU/JJjOUpGS/Fw0w7ADI5KLihNXPFIE4ZmZI/ARdh50DG19OlO8Ef9EGo
9gRFKJx4tU3K2tgh9MKossMwUE6qbU9oNaYDa/6g4E8TeWgmM2vGlhZn5ILXeohhHi5Es9Mr+rxt
HoJ+La59A/4/ru+EoDyt9/Dsoki2ct0ruX5Zy5DkMTORIvEp5xzzO38L9UsQ44fnnIgw960pzoxr
ktkq5NP/Fz3r/6fXYtTamGANsBaGHWFA7MgG/GqOaHAiUiPlAuNrLcvr1Re2z9CRQopKUaGwAWp2
EaAgo7gAAKwEwpHoCO45aONBX9rY+P6tJBwkEMUly79wx+RXySkb4GNEKZ0Gegz/w/vfJL9awz1Q
EVHKwYWO0ONEG+H0Y7tJfmhYsKiTp+p86UK7jZrd6bxNy9fIQ5YM+w0iv7Cj7SZUsST8ZAX3Vlao
O8Dt8pC38TChwn5SQhfvOCW5ZWojMItCLCkqS69uiZ3llOXfakNsBGajN55OyX6Gb3wkvhTPpSPC
Pj6wS/Za439NPPpatoCq7I7SQT8ryEQE/b24qeiE58uFabMoBOgb73zVrPsWjwkZ29dxngn+jM5E
7jxA8LPaZIX+fXDZSK2HLe7t/BSkzwiiSLzpUNMkGPde1EkUg2V+QVIShoHiQpLpCrnbSvghrdlS
K2yAncGsB1v7+9A6+V4R/A7jSy6FynhqgJuPEiGnKaZJIOP5OZwyJMvMqOx6FM1+03x9rBlm7R1W
esbQELwEUmQcBsOlWfaSCHLN8TOnigt8ixS7qxs/U34Mojs9CQV8dYygikRmf+H1/KEaRsi21vZM
NGyNXm5qREILQQTv8ho2pMu+m8C0PFJ9AQ1F6p1P0juxnOYmgnWWAcNd2eJ7tCHT/RmvZRPP7QNC
kYM17q8OyzqJ3rt9E7GL2dEhqg6GxiK93UqMCBRm/PqYynnaNTMvHnMigJqS0Hl5L5YVyVxLoRQ5
AiMlCltRqoic6idAhcw8upNhZaCD7N2WU+FJG4tfCDYGrg1NqEvATrA/aWDlJYviyLbEja0LAgTp
QlPTkd+zBFCVgisKaz2vWF0jCj4dG4Fp/Z0g7vzUtikUAGfNKBuSK9HHmBzdR5TlZqCdrB5JeJHI
lKgv4fo+QA+VlPZnjiEZTS5UIX7opUgrcsE4N/1WIjOv1yhpFy2V70CcIZt8bdhGUResBuCTpr35
4+fMEu/b7mncJ97GHhfekCAPdVKoE0UyExTKX/3JIAfgRY06JeMy66RAe+LLrtxysT/ERMoCrEFq
AZMnAMndZ/UZPnqTuK1QGv3mT96h2Q12gWAjLBYODrRo+T0i+3IE9YJWj+AVNRA9DG0jtpGRdb9d
0FNcahCaewknrHkbkib5Mx5qeNUW/66zof5CF+DAOwsibPPnTeTJctQYQLkfXE8VdzqtIOP6cLqv
lNKJ7DY5zZLp9Ux5tArX7Ka2ekPVLRVsRscd9bmUjd9wQ1RYvUUpNHnyAlmQ8+I+Tq617w2W6mK/
lffaoTcfYOnGhcqXNLhPMVArEzjkIE4Tp1LyRG3NaCP526vof+uskfmKIXffUfaUCYfptKHeaj+a
WiC3tJR+CThVYG4PKoIwM0hUalaqwn82hRzEXw/SDIesEPUvBrIGi90Q5vJyz1ewt0C8vdb0MiYZ
fvodgSN/1Nk6UajCMkZ7zLH2pTCanfhb0DcFDZefzjvoXzhg4PSwCwIwJGoKnMdddiMXtzc1FHUy
69g+8/Ob9U1HMliWwOQHQUwmNrkm9X3IUufhZruRnj77EbN/gK9uwHt9RgYXh8nk7LzGEA1m7RZP
g1fzGwUFEfanupIoZeU6GxZbfbn1nf4G9HN8PtD6Fl7Ajc1d7p1zJWsqGT3P/SOXX90+wL60dooe
YrVDkOMHwQPybSO/eifqYb2QuES9Vav5PguapqWiq5LR9VOSDm4ZVHwO/GE4wax4TIF77P65pHLC
TxdKrBn7lqxVQakGNS4eYz0sZHRhFAS6s+BaRodx5qS9iPCx9gtwpazCLW2Vi7E1AJ4WYDsfiMPQ
xfFORrOxhj/c5xEmV7EVp+zdTUoaDQcy83TFebw5lP5voIy8DjCTvM+z0P7Pg+4/cNO06niySYRH
porPKQLiXu/pf7n031QWHXLp0O+AAP2Ha8Rl7YizUFs8+quWjLXRf7OO4DcrIviIgr6YsXmHyXtj
kbzNwE9Hi/loAAUqn/gqltKMc0JzP3g1OMJoeQzLDeuR17uoSXsW2fSVPo5G+kamgu0zncKH36BS
uvxb4/dsADuXTYB7LcR/NOFLYkJ87YF2u9sphjY89u9VOBLnFFpPS1cAq61XP3a0FfpIUhiXxaj7
67Rv4W/o/mg4pijpNGP3jwgvxIa/iMluzOup4Y0CQHLwi9Bn4xnuAdJsgtFBzPheArT+71L8+2eI
aB9vNkaJNeOjhYSQHZ0kvIjiFq05v2ZnWsMflYuL5Fri+w9oPzB6Tif7YfUMFArc1ByVeEuFLMbe
vbamw887swy2srOwEoM95le9MClN+gfRuKgwxIsSFfvyNSnMlPZagU3EEBdOSSetm7xChiOUTitj
+N5OfIHYuxqezkNUDMslAFTKhTErTegVdqjcnfud+q+v2QZgS6tYpGjxVmPtbvfIiVynqs1eHBkR
lAxYORxgkYn2XHvFyKMuQyuT0BOHdukvG4mtT5D6U+3mwasseOWysOrP2vcGG9X2mvGnMJVSwtZh
fFaUW8ftRDc1lPqEp5JZ0Wz6Y2djSW5SwMjtEwLSkEfkXVzTleJH177rW13R1njcH9wMPREbNQ2v
/JRrqKOXFqSc56qyVlGa/uKVGxasgyYBILmkReSb0FZn10/BxhNKaoVePi2crWrqR5pUuMrp3pRL
Z4E4nhmpK07KsO3iT4j4++LgaH7YOHi2SLO7gQWTkuotH3/DulF/GsYnWZxWg36EiIcsPJ4gGcs7
aLjKPLrhC7DAx7eLM7y9Sse6MwPJFLV9vDD3arTpqD3Ao6xRP7Hb5UO3EMHR64h29Un4AXTUhx4v
uLqIhpoFridsjH8xhNCzp2JrwmCc7Nj1ydXc7CfMikeg0ZamcNNKtSin2v+yazwXoH3hCOr12E5j
xg6fiTyLdi3ekGxQjvPXglLxxenZlpaBGuSZxbYK2H9K4dItGt1LicMpd0DY/axgJbY528rICxAm
JsHDEjtRobaAeW1+dDoaVahFxpnas5KJJ1E2PqUcsAYQ3yWsLDXUnOGJAs2F1IwV1x9mOBKPvpRe
Ne3UMwxsNWuQqkObWBr7LKxO6uTt0oIWL3sJW5ZP5Ry2GCEhe0HbW6VbPW1i2ICmTAUo6wJ/YKUI
lokk8V5i/hUtnCj2gHdUVriaV5o4Ia67ieqM1XTYsPkTckqH6pKaquqNYJ8TjKdYmQ7Z0C3vZwO7
A0gl1zDyI3BVZkZU/JGuW1cBioaKqAKcJmWuf/WtlsJfOG4qPMcxOf5sM7WGDVOIIbDq/cqz+dn5
GYOCO0aQIyxeyQ+SH1iuZePCSdfRHk83HNtJnmX1K2tjeM+38gR2G2SgXllF+H2ktuQMJITr0re9
/lf8Z2crSz/KtZXtXR2QrsGhHtEhHb8vVamqtsALbpB2mRmcUVB8nbB/YHg9TgqeOAjOygb5kn+8
tqx2R+ldVZLGJm4aIxlaAlfLTyGiHWb6ZmACmdWOoslqDzV4BDNIy68Rij9jbWFc8aKnWXINrruv
hQ6DA/ihVA0wUW/qHlBIv9U9F/TVT5bGw0RYcE4iZ5mxnlBo53ETyKn6FqdUtN5Rv/K45A2MI85T
0osnuVZGty6hp4P39CMAQR5eG8kpNfohfzyMR86zO9vHdT2Qa7rZqpOTfJ5lnqeepwuQMk0id6pm
NbiDrjF0uEtR5U7D8HkuLJFZAVuJRUgHFWKrNcsIJbnEhXojdCzSy3f24IzL3sJQW6lT2zVDr8Mh
tGLnWkvJ/aMF+Ha+ReAVxi0mD/jqnmRhxN49tw6iRYYYJWbjA/QD5B5Uq7vM2WDUz+hhGb6BhazM
jTWTv41VFo4nkHRfxW9ai1zdsEvJi9hFBAeAkITbe5fu9dv85uqtPiE2aRPcOncl6dcU8zs/zWtp
DNDCrT6GX+Ghz/tVC2jW0zxALcu2aBjqK7ZYPccelsAUmK+IFPOIi0ln4io/pS21ScmlZxzsimGP
3UhZPMdX87WFt7Nu/Fs1PeBr1eBfIA0zhT8nktK7w1d70Zh4qDwXxwcQeg8q5nn1liZ0u9QgOfCP
OrA8zgCnRBCuqqBAPfXTG6b4eAESV8YLWSyFpr/uZpQc9UYPG0l7W6/iOXUIjJFYqWLQlO4cAktb
Lvei4a6gO+Lc6aV6FO6IMEiV31ls526xKqS+/mTYqpEouWotdXSiLt9WKf6Dd8wgTOIwJ0/tIbDp
BiSe78XI4MXFXy5LkqFcT474RRZbDYacjQei8yHGlHrjfP41pXD1PXVl13QcRV2DzalmFyLJkdmr
2Lx8kjkxFmemgTwGYcsbmCyGcBbOuKccSEiVfWGQgq7DdYuMgFBCXQ1QlbrHJue4HzagmQHThS32
hyqIj91+LTOPaHhdRcGoSUlxHlg0HnuuthNVO+8LoTuTkHZDVjCgBTMyjyQGKhwr/d4SOIBHGytT
8kDSYiqyng+QBf6dTSXLQ+AZ87o+t0MNCCskVbbbttcqFRjoJVu+8j+m+EipMZmsCzce5sZT1V+E
mCLoV6tDs0tWOfNA1j4AkC/WmBIGMTMX7hKx8bJUsmjhInZm3g+J6zRsF41GLc39mDhb9BMfNFVE
2o00CEOzzd8/VSIVgd06qWbdxpgxL7Q77orfYPwwcqHzPg433hAktFgA4FjSZ4jww2SdO2ibFKec
slRJDZnbn3DjoxsOtOQE+QhKeqQ6a9bRlEUIkRapAd88jXpjnP/+jBBG9j2CovfICqq+ZTmkGx03
zmF6Yq2ywjYWFg0AEtoFr1BTHI8i12+zZZvPmAh7GlJF+jSJmIlsBZVUK3kfwH0sR4u2ZRzxVz8q
y6T4bVoZcBTmzJ2cfQpg7OStADS9JUzmxfo4/LPMQ5qQ5N8bdkNHyUAlopNAg21nzso3XRJQl+0v
sKuGgU02PIwEKu7eTN7F6zh3UITBGbmyes4oDZhcus2ACSJU0caiGUzY9jrKvwrj6yySvQIGF9pv
QBPv4LNQDaE0cTGTG1PLlEdj1PEwOzf9GjmCKucz6mw7U0oXy7sda4S7Bw4iyOvetPZMzyt1VT00
FjyShyl4Wd7JEIjC9v70Z8KzYB2AlZmi4T/4DsKzO5g1Oe7JroI/ADmd60EwLUZ+SitMRoMbC/5P
O4dOMCCoDiX8teQKu3/s2sUtYvrWFOAU5sK4jfGhTswOf717HfNX/1qgX2c6BxDN2/UmxDNAw5/Z
0fbNM+oI744/PjmIIFsa/x/FD+YqnQVCFVYuDDhMs35lC4SyS6uJwYCyBz12UlxXh7WgKNm+A7PR
Ci8oFgtYYqpn9ZspfXGIBJgnzJJrTFkSgMapq/34KNl8vNw+IVSqaYME1+/pZU2kT71aTson//8I
iHHsEVIJPGuTmyJr7xnpetg20/1N6YFe5JJIdU3L3iaROgUSk+3IixSuH22OiGZOlvi6q1z3SeQE
Qeb7bpL7uosVTpr2zVxLR9g+yLrCrj/9Qi5Lg7wz1r9/D2dXetN2dGCneVLwVFgMtcRoycePSxLP
0I0fAka9LjaExtFfma295e/U9xfPeCSAyNRGKub53L1vKOuQ7Bqan7d6Jafnml3YhRffiYAqYHa2
p9i54pNKTlr6X8HNJIGDHLjq9g1WYxzREGsXLCeKJliPkgZHk3MB1Vj5b1wyiQdSONtLN3j2q3lB
1JgO9TuJf59ckePFhk8WNbXd8sJ9ikzyPfjb5fMe16tMycoAm/zzhqX8dhSNVoN9btqxeKv075c6
oFzd9D0W4Vz7Bp9CB2djzi3yDLyJoreg/prQweEHAH1tAHFpszFHB5+sZcM5HQhxoXPD00iCMGac
lc0Deo6aEfD+e3GGNlhzpM3xn+B+kTC5Vwg9cZ32gslqSg/CkpkEDYjZ0DiessuX+toon0n2uE9+
j1I3Lw6AQidNUUGGsLX8U8mvh6dpNM5Z8sofLKz4ucsPyptREOoK3wFy+m3vM/CuVOzxJ0JZDeBv
EjB0IlHeM/dM/BrESlJD0dBZu4N7lFaEuwuPRTtM8wr5HNa5Z2/hnnXSiT4gy4lAsummwQl3t2IH
cqrEN/AOEVZm/7iH7ZrO5h87NQMKOCU3HyUUTCfADqFBTV69avsHfpYM+QIeD4yVagnNTuhbQ79F
jOyshHyvcn/TitSwGO4NTnEljNL1BMn0fsz8t8cX+3ryyrqrak2b8m3wEchk8cbLlTj/SP33ITqy
EZfAx57dwsQtvcdcqKRpduXHh1zycK75QeIRLgLOHs/CHFhBBabGSzO7OE6vsTWfgt3pYoR6kitL
vvX99Kl7oZZPywTdjpeTTipwo5z0aOeefD4iEWboXfZ0Xo7t7oA1O8DCrueeJVwvif6EOFX+NJ2V
YV14wL16bv843OTk8SDcjaRqffiAsdg5CQjEJ86dI7m9HAd9MzwU2hklFNrLFci72u+1KUEPJ4y3
TdA4E7XaCJKxF03Ag8PpCsmNP3+vSe+s7h6ljKZiT8BXzScBEJQMiB6lmaPbf+0OxUdixy4y//zs
tVKWXVJPGUry/mRjAI0CRN5erDVs3IP9YQc77XrJbuiVXyJaFqpJmztYKzYzU4/mqgOKYAngRZOt
uvRxD2ApIq2pa59VtvedDaMZ0AlVKkaK1j3tO/QHGkWdHL9bxsq4sjFDiHcMos3Pgow7D6l+biVI
jJXwWl58+allewI7Z2iMOXTNm5sHEPILEIIWTYLcfQ99P4+Xdw0tdSmgRccT2JhDqEhW8WWkntte
rSlCPhlmLGOSTCJoBYMyCIi2HmI5YHz8Npbz1m7zvDxdTs7eBKzEQDcRA/FXnc21Mk3N7AvaPUfx
IX09boXSfC9YAHAjwn7B3vnwgUnBHJ4L06ehib9rOtw9pBwgrM4ZHYJ072kueqNEumQNq+jkiuv1
OWaJS8nKrUvq9rmDWv6xHdm9WaKQZUzEe4lQuPd2Tlit60HU0ycyuie+RSJtIXdXjga0mRDVaCKu
uDZjLj3WEoKCriasaCJfIx4oTI7eKByWZXzaNJyO6N/7pcZEadF2lEwpsYiavpYwCfp9SDydzE2N
KPoIoUkoMc1tEeDCcw0EvCHwQlG6Nk/uLRXrpQtxvTatkaoLD96dODtAWCRaC/Nd7RFrBwR0RwTk
Pw3LaN+ZwwmBN20O/6iGYG8MWMlFo93iIwfwrz9cSHPX9I3TBNOaONp6A75TfnOx6IpBQ/1DUlyM
ZPmFKrSaolXHQVKHJnvmvrxgUxU88PuuJKxA/6ToEmehXGzRjUq1aeBx40xsU2jQz5ytw+nL6GpG
/vd0gzfqvxVQz2D0bDKSUEbyjHGl6HepoGHi6kmo0VIas3gXQuY09aRisDaFBK7S3+A4k2OW/tPl
vrkSYqH7sI9Jax7I3e5gn5utiI8rFOK2m0EOtCUgNQx75GaD0Vl6adP4aHVOh2tWH0S5yqMwcozj
jK04GPaOjPQO5QVMVz4RmqdJlUW6ewkMMVrDVaEHh/6Ewr9DqHty4Axf3hrQvOc453WlrB02fRxe
ck/PinVHsHu95SvikJqu8ptD4Ne3EnG2FwCY1TpRcc3VxYiFVpCVL+vG1HvYybmBn7Dyav1dPy+f
TENpot4rt8gEt7ia5y4M3XGCrHxRclcKQWIrENkdFPWLP9lDnUz8P24dXzkfsnuZG6ZeH/gKghn/
Ekunu6KOLfQIXNoHkWAxTWAKJElxLZh32aeqG+4GHTx7wbbyLEc4q7DERzOaMdzPww/skLQJDlwo
YIBlK6vPWb6KNoskDab9h637edG3WSYFjOM1aM+IdaJdniBHH1Pjb+YrVmWrcf5LNX44imGvmSYi
EBll14Uy5hlVrqx6WpEWSh7jm62IBvTS8qdjAqGMLxfTjlREor2npxfaJIdqoO1ldWpwiu3VLBqN
vRI88JH2Q5v9wBj3tcMYwciXjwemcziwjmRZ8izP86D+5hV09FAtsfnkm2GCZyJS77+AQsOzZisC
q6jvcx0RbrsoAlkcYKF9S8f1PuntbKMe6f3XseZ2k5Q3gY3euTmLBXYfbodMzruPRKCm93b3yhMi
2kgYLkYG1/H/x4sRfQ6S2194IPqT0DRvYNvmBx6m1M/Bb54My37j+SofWfbTOK6g4IwesUw14dIa
ITKHqBrbbnoJ3lQGenUr30cpDwa56I/20WFHiWWjo+QChWvhNyN7axjiQe67ENb0xMmLc1NAYr+a
hJMrtRGj11j849NFCilzlzfUo0d+DRjmCaM0V3o2TlsnYYEqZ/jYscKNzv+Ziq50llNOwYqB/Frm
CcDXwGpG8l/1JJlZR3zlYq8pVbN5DsK0CC24q7x0Gk3CpunHQl7RLTIPgJ2iu0Bgd1dpJspd4hLU
XqQMRkVd4KVc91ZQi+Lziz6bhsSd6J/tcDNHibCfDoU4rRMWYiBJVrHP/jcZGeSJWyf4P2xdU1g5
7o6HjV/YMWuO0WAvZLj7v6iFIKvQnis801xaxc4ehRJ13Bq7xb49wPqvt/bSSHFG/3X7Z3iqA6F4
L2ifsFiVlEFacISF3jevYGh3IWS7et02aMyzNpRHFNC2sQljNzk8cIEOfeJ2ruu0UXXsfeeg7VXP
SOALZ5MVVIu3Po2rFsOupPrUb6ckN6iYR9IB9qg8jTxL4fpIMdMbKTMsfVmhc4moKZtoxJ27bTpD
jGHuYOMtl0BX2e44kufKr+0eccJ8y9KqcTvYK9BNo1LMCtJZvilEu4pQNiv1x/VSGmpJAJ42tCKZ
XVHY158wayxtP+MhgCwyEAu8s3uzj+N7Y2Fjf43g9jS3SYuYiKsttdYw3CgVgSuSdmMZTgDsHlF7
E/GhY4gLzs3uv4VHWP7215CxTHfxNHV9J/Eq0YSraYbj/2N+uM9eCNKtsWKadGmPo4zAdIcWTiqV
pEMlGcWG+ivOIGbRjUnUV7L8L6YCwJ0X5CfpH9ZECEhj/ttS+OH4/JhGXiZ88A+cQztLceE8mkFQ
4RW/R8QSwKyCMihWLKR4MGYCRez0Vlwx+jRPzkxyGw9s8EKzTq6ujpaIbA0PIg7LDuv62VLZlSvW
vDuOSHPoGXF9iThyq1EMJtP8d8q8Jo6kgalHWDMriWLB47sc79zQMRaRLzEdZpSoOJMI9AvyuICo
4vcjWOm6CiA3bCdAITCft/cYnc1TcC/0r06MdPNjU20fTtQ02LRRI8c3nU4x70TwymFy27643N2N
IbNyGjwWac+yEV8zJSgRkR58J1po0B24x72/998YrNQENlXoYMNentfH1dr1GZLuYAOx3gWoO8B9
DyBWB834Mm5bMjIQuEOb1WjtdF8FEqTfwaVwwOamCnvHVXuJS3ffQjYblJF5w1n97j5Ustgrg/hM
faAga0tQ75OTK1xnPFwbXrmajMsF4oAapZ1hu2HogMT6A8jZY8WxYyaMb57RxzGHFKhsyU+ONh6w
CljMAb01AojaCU0Uvr8jdyIuTfAxGCqc/TvNXdJB8VkaE6wjKL76MEGe5h2Vix1ruj1V4fRTF6eE
cpe5ofEPX7O7TsoJgP7ojlYZ55WxnFY1YAaH5EyoTft8IyZ70aD22pPmKeBistgVOGmSedWGLzvF
KmK79cG/X5sNBtuZviLRgZ/I4XL8v7+ATfCsmRZKy+qbRdpOEAWfE9IYQG3Bi/XWga/NlvS3YD6Y
EvZajyi5a6z5xJ5C0SizCNvAf0+tne7gaPOo/5Qk+7FKQsnmC1v+0BRxXB80hW+mGhU9Zxx0V3da
1yQ0NuAxfUMGL9PS1R5uicUkXyiwEGtF72i4rDCB4/5sL5U1yZhSEbpTti7K2Nas7QdbmG+DYXKF
PNilTwtWWLLaFTAYUsO3TnotYYE3Z/10zh6/rJj/ex0bfLH5m2Q97Pb5hQhXM7qWaH3L8/c9dWg/
+zdYQd8/bIZPta/n5+Ics4m6Dl3wmH+zIMTRTaf6+2BzarJRa+uPRtErKxNCWIHxoeZk+qi0ihiO
iIjapLiC0WsHVBNe/UsFhAuTIWKgIDYKSk9QQeYgs8aL3a1tiKTwUizqG7+QXhbIQPKWk1hSIELR
0KCn0NO17JEupNUdfkKTvjKUFBF+dOerFZoCNeF3KKIM6IH857DBpQIsQ0n4iwXNhFt5Yaaa0mpk
1/UxcMsFuD3EWQEHGtkfFa+rTGd+0xNlrsxpf6xt31Oy7x2QpV7MmMaN5uGu3U8/J5S/RQOzExuU
2NsyMyX1+uSr8AAnjjKXYF3m21GKiH1oPK5+KKuLutMCzR18jYjErwINM9Yv22faki5gyo2ibg9p
COA/5VWctiAcMMKBk+KovSKxymViH5LBd3t3MEiBlaSCvageenEwBigW5mhOu6YQajJPjM9ZEU+M
K+RBcgrEVSpLHdlRWHyeEEm0umt1RfNEtnX/Sli3d5RavDViIjHtfR75896IMFPttDcopy6/WwWv
ey0F4gJj0Jt85KDSo1U3TYNZMVnRCbplphUvwEzEHl0MfLS+UcysbWGQmYB2Q/Nj8gpafw0g9pOG
jXYQWTGjdQ6t6qh+sdQiJyWmGLVcspgjZ6IiHR+SbB+13fZLOBbb3d6QVOCTLG/KS9dqPBMcNlj9
h35/fulNgxB5Qf8S2ABvcyHZ03Bs3orxQcchq7NJgJ4vXqgpWsI88Taw66/8IXPcPOvKLss8+KBz
uw3TeAnldKoxi1EWUHYHp1yBjxf8T+0hw3nSbgA77xHsVI35cgIvfoxOzAwJMsm/Nunaw6Dm7+Ib
p/6gRq8djrdUsTG/e3bMycwUumTfUn1lP946gF2gujC3Yad+hvAjNBfoz6ld8STTKpkyu/yIbgGA
mi0GeiXPI5Oh1GQt/2+/zwYwPGSBGk6NuIY4VUdb3Q5CVAVMVJpjZVVIS6JmZ/MScv98z5Kl/vuO
Rl9x/wU3kJG3CHS2s/Aqz4QVBAcYd4lq7HocihiC7S39kEmkfiMS4LEbsJfrWoaJR2nr5Jh4oyv6
vKuzuxwTTJBOX0gTY9lX6eICcGeZSf6K1DHfwekXAClpMM1WB978asjVphbcYtM+vJnfYEogj9Sv
2GoXrsbX/TzsuxpcZtn4UbYup27vSrHMoZHBcQXwIJ/QbbNYMQ37INOQrYLKV7fyIe6TGTA0bg2M
bmi3c2PQBpunvc1N0ZGpRjikUnUxsWEaMwqYOJqg/mql23SnWmtzVTjnKQXh0XG5v+iU2dfOFNEj
FHsHgrPZ7NKQeLrCYeVh8XHM39Y6r5pXewrxNFtqgueoYPnCvycl+XT6ww6aNdVaELIlnoWz0q2W
un4fYjJDfITll6aAe4FDd23kCGHny8fNtEIxTYdSUl6nHmqsTgN/9G9NPHzWvGt98r32m4kFSKEz
8Sv4RLNEScYF3xHD+pjQXujtGexyJrntLMTT4AD2Z740GBVKefLQQ/lOv2LN5w2dDEKyHNNxQIMG
nLARaJG3vdPUq4mYqVAb3jmFSM6ZSkWieWioUVUCY/H7mp/M8lWP+dpqOHjwfEAhFwJttVPTrnum
bC5DEWZseNePGVUDVeY4diqpY651iNbiynb+Hh3xJJvXXj132VtCjBftuwWs8XrkBSb23szZ8Tt/
qS2g3EoJdW5UrMVey4ztCA1Ba5p5QC5+zG6uiUDnav4xwlV9bW1Lg6pOuQEKM3LRX5tMy9ik4osi
PwD9yQEJN02Mi+4D1lnapYDz/QCJY5GX6BcICw69Z2yq3RnwsKEcWLQVWkPIX7yVhdqGu/8Qk1HX
/aJc03OOMBKO1iAG5zETjYeB6/8fFxbHtBybZAutBW+OvxXfRDgZyBOOhTAenuEWMSOF980I/rjk
Yy0KIEV+IiSwjRo9baLMiCo3BbsN3hXJUzOg9D6IxS7S3lh6phbeVM57NzfDJ26VpTv9bNLCaJoV
6S7oFWRkP8VFUu36Wudm8sScXfv4K0aGGikGvlrVDMRTL/VAsQks1HX/lkSJ0vMa+YjdmJu+DXFx
JD9lXPc+0RVOBlJKKT1fpot95dwk71jz0+wJ9rPegj08r4Xan70KtQ/hJHLvX6K25IagmRfYILir
BmL09N4SbwwTkRoQX0zTYKpstp2WB2DiKjiva6rBTpCc7uqseVttkoFM1rCxUlgt4JXMp0g94yjh
YT8hcmIv8s6lMjhqlpN1SmzI0quzDu7+pBpF/l8f4QOQ/x3mIVYZJpSQ1sHaH82WoWmbk92btRMY
ejB5u1/jA16Qqcy1RUnL0+X2CzllLqmblYD3ZqRvWnHqlKtqwxhf2n8SmbUROXYLF+FfewersyY+
KcE2j9/c+00M19ekCWimw7ShHAKZhxZqoUFzqaFQlrlNhpjNlkCN0yCvss87itPP8FwOFtCLpFmP
6aNUcHiOqW4iQ25LkERYIXzeA9Eow/DJGGWjbi1GaxDsbJ2wZ5SRLa+p0okj9zVX9v8+xkCpdjww
xbNLFT+rE0mdJiG419YoF3q5kxFwF0L40sl7oIk/rhCbdotykdpBtNd7isJCkukzUenLMw7idmTU
64XZItXU74a8juVuOrJf1caCMfFNJ4Bcrp6IHuXQBOpLdxokD3zz1zmZXcRxxR+zUwuw4ZihlL4+
cLKZtudocP4ipXoMA7qdRW9L1scFo5DFUwnTPHEr3YJPLf7MIW3b2D4Zvlcew1XtZVKC6qLCoS3b
M4sHlIFAGWxGoxd9zNlb1e0dj7luR0DJhm05QwfSnHUvjz3wE5I6u+V8RltzV2uWiMBJB0PM7LPv
jXarv5/yVzG6OJXz/XQPhrw+9jIs6uZDFUuVNhre6tE1/ejtoxCGakm1INspWHPsUxpqHdhv/QMJ
4GDoWqMBY0xjR/TWXEuHA1gS09CkQ10vjkS+XaHOdLrBquBi5ctVUlgoylU33mV0wZqnU9TWnbHx
4wOXsjEkpC8tTm1DXAlKAPU9acV1uXuubd48OlCFLabnhPqby1lqPa2UX5WH+jqnXxyAhZUmtTsu
vEikfUIAZ+enXMSx1Cs+h9abSiJSEMca9ZKNGYifvsuaNGwM/uq1LLUBVWsFlrbZxyef9k/XNLZr
4HIBj+WxL6+7UNU5SdixOD4NTcMmT9LFQqT2Z85QwG4+Iy9Vz1Z16xzsqEzJA1zkbxzAU2zqN3mY
B2Q3qMIyU7hgFGMVKgGzh74g5pBiCrhoevqCKXevGlT0clqKe9N4uHDoEZHwVOLTIQBVNLXP/R5j
08/Vp8MjucmhTS/MGeufmk4jWxF4/6FLuLbVMnmfpVAN8RBqgOrur+kNv7rrEHfolENlsZ6M3M3u
olDZV0MCIf348t+Qi5dr/aSSQhZaWZG0IZTe6lvfRbj8TJopTnA3Dp5v09go73SK2KibG3PXp+Dh
8c8itXT/qgYejxgPVNNKeK/bc8gBplVGh1S7vVAXHZRe4A0+cxzos1IYygyJaWfrCSqXkjRZAZss
fZipZzevxTOocyUIC7gXqhHqJmpF4Wf+7FjrWVSzbFOyiA3SiGfOUPH+uYIGji2lYcnF5ED+RsDv
QsNphTTZsEJbpM4CKQx2f9BiDpg5ouV4FYGaGOy+BsQjHpXSJ7fPe/CqFZkYhOa58Kpvtlm0AWDU
YdPIBKI8VmUo1m509a6t+y/HRU+qCPQ26ZwufQrVgr3z/r7MGO60wX+gdKBhwTRCKwI4oYd6qV85
UejNcyy9v8o+CDEwiZV3G1c77tcMDcxrvfYNLyuCFIRF6PhiCdKbRsslI9vHBFsZ3PljSaFVjp7k
jKok/waOVSYLDV4WrB9r5DgBYpzQs5JRb2zNPqUmZFzrq/47X/j7xXuTvK/Y6UOtbPpJUJ7Md6uc
ndBcEqOuNcf+f/4rXQ/qWAvKmoV1FJQ/onM9G3cokrYLw4wNCAplK3r+WmWDmgbNWN0hMBv1dl5G
/yGxJ1xH9tMqo5yhIYOQBo6uoBufW3A1xe9WHMC5wSRo833GDdmoqfk2ZnelavmorpbMGPVEdF5B
YYs0q+mmqV4wDFgdmH8iOcTgxT7xl5B9+/Hnf51z9p+m4CLlgsKPQHoAdEX5RV75GBOPgu8K3P/n
Z759Sk6OPBlRt+ifvbqXDhj11yCnI1XpJKr+R1poKpY73CeCyEi0J4IvpntKp+CIxr1FIxMuYuRS
9weYDvlFCHoPPpJI2Rqewv5xVaTK9DjHnyKRCu2riNqqkj0J5tDexVa3B9SIpu4Na9kfMs7nHG4o
VWfn9Jri0HgoxglIl8BvBHsXqWqD2yBTm9ot6URie8eykBoy1hvXHaWW53RMSNFphF/9iFNSI4hF
LfsX8NyHSOjumXTThTx5Pxb+gW+8ktdI3Ofin7xf8Bj9XQysQUnKPZgO9c9Gd7XPs4v7xcNOmEmu
8FmpB/NYaGfwW2TEVIhKHlr4lYp+wD1Bcw9yojHjuVK6icLl0qRs/m34MtvVsjQkt+FegB+xcQlv
Vg22Pt98PYNiRT64bkzAHpd8u/lYi0FELXsM1jpW61pARwcITbbBbTH/tJ0AZF3EEBtbSYoisdlX
rMxy4tWL0CHTDPgtR8bzFrugzqd4LO2HwB7+J9/0rmEv47qfPbL7FUknQeppYhOILlirpxAmG2h9
aIlv+zHDncooJa8f4v0ovLb6+RG35Wres9fgLPpmGXeo6rrdwMQ85eNGmn88nQ7javzDOMkUK4LV
bEIDJrF3YUkMRr2kA/kOO535bCoPl+vCROc97WW2TgQWks2gvfVGq1iKGQOFk7fvMQfzJcPfCiO3
GjFXhnKO0FEOrC81YoEiJ3rDxWJNhkPFMKY2hoKPVYmBVxWrVYVQ155P396/Ao9E5GsCYNHAWQbR
urrA4avLiaXtwj9Zdc9Smx0Tn4tjlW3h19TPmuNl8PrbYr+HuWJqJz2PHTp4AAvh+VEUUHhvAEdx
uQLKmTXjqdJExjDY59UPF8ct7HNA3K8ElNR6wBMCQOCRAcTIzxdVabfgv9aOu95Voizgu3bsBP4B
URXyqVdIc6K1l1NCKYJb4BYgpMiY0/KuGkfVvqSjt7Ypm3ew89/XZCyWznWmJdf/dKRrtakHpWVP
bcnANZJt8vrst0GCHDnWaOEV2JMixhh7k2BDTEDOKmq8szIGg9E35IoGdNHuAQvVp7f0x6hCaGjR
nnDYdUnSK/L755IlprDchTyX2SRm0uLk89nafunCMdHsMO1QZgG7kr6ZFedWU4LdvcH+PzVV8oFK
g2PHeYgdaTmPZeEJh7hK2ih7B3CFhdBKvKcZUGKHjLA8aHHxKGZOXZCpv9MILoUJuMJmHcSZHBte
wENhFqZJTdBrnC6ma8FprYmq522JPXk8F74AHBIXCxeYCnnAHSyNooCcen4paZF7JPkJ4iPudahZ
vUoPYzn3OJriTnYQcQuskRFRDq7eo7JSpJssMvyxWepO24vmTSYpRtU8I89qHEv1oeHIZ/EaXiQb
+Vh2spTj95Bvbzi1DwSBTbawnAVffBT8erMnbQmY0Bcxj2WAXzN0HFlGtWIm13kRpoZNH+LM0DfW
3swUeFMw7VuOO5E8DONsALLUgtDP4yJ1OYQncoEfndbmIQgXJD1tNoC3tz0Fpp+EYLAdKu9sfeQV
BuJnJ5eiPFJXxKgPe7o5IGKhuGspkdywsYvejFjSg6M6zzuXWEKsxw8iTP8IRMjYQzPIIOxjjffT
AlQfzBOVu0HCaYr4hZQiYpRZhHHNC0m3/FGknH3nWQ5DThWqyudvJd5hiOPTc6xG9YGt3MP58Iow
gdiKvi7QPolV1llW1ZYUeKuCt0aDejz0PIedahKNpZ780GXjn+r6+R1T35upxQPXPiHgZ2NegGAh
JSXVLn8jb0tryVC66FGgszzj0cI0M7yY7DceWttShvujXSd7CoW56Lq2kEZssPUtU427bsGBbiFO
1HmPZLeVOv+Y0ia8CE4+gCheyuv/G1zsQ7Nw0HoH6LgIj8TENF5mouIvmJY/79GuVkSI+tShW8Ze
kOwys95WbZBnW5WjBYSac2ozLbwNg/ARe166Q3eKEUNVkDYCzhb2b4oCRSyuWwtw4i+gHp7GJhxD
0h5W91A2orBiCwi24qZUpWYOXBhT0ncn5FGjGDURanojXIX3u3XvoJZKKo6rJlNqcAz1efYfFGtM
T2VvB43USoTyD+pWX5j5i/yDc1XSrbJZIzez4d/mSTFxiuQOxySlKfpccUi8vWN4j7T+9iwgqboZ
RWKTFIwr5nD3nlJWxGNJ64Vn5OVEHjb8qoQgebs0LQvmFFzs0KjLq8QCg8ElBZ+LIdfRtIHo/7s1
U4AFFHSAZQYu6/4mYuebPr2GqajEuOFXEv6mzmxCnbsf9OB9MBQJApUlCXYMnxaveJ7Tf9ltGEb7
T4H312rwU4kYKhudbd0XiIfuUeEcyq9HEe2wJikwqSNNA0mdvCPH++q8jzG/d2ObQxpKtATZWLm5
8q0v0TarpmAwlubpUGW8d1ca4yM+uwYJv9fFO6D9IcuHZOF/lZYf8jDSyS7iD5VSHyK1obleBZgc
hgY9FvuD/1br0TLvdd2jH6XrIJxr+ZPmmBj2eO/9sKf59uoDpzVzmG6nVaj5h5jMlHUfnc+K64qK
82kMQtxFVHMHqwB8SkjgtrzDsuMjduv5fZU8ngqu4menoznPjaD3oluwKUL6ISyxjm75GW2rX6Xy
2phElR7n3G/JMeSH1Oy5ZJyDmRLmocw+dcYQ2jfzc0r2QcM/7w02sMj6FLf2kzfy+0UTUEs2TM+w
F1/9uABEkIjpB0g8nff8GtfIXQHlWzhrj0dxcabMzZAzq+HlfxNr+4wFAsBNA6UYlpBsOlTyKkkl
dJCXqf5svfWirq4CrVNfCI/nnF6gknTivdmMelveNWy2LEtYbwrRy6c/aFLK48eyelqcJXW8OXcp
k4LHANSc/K1XDX1fGwpQyapMniPJfv3/UQ+HdKELug3inJ/dNwWMS6uqbtQ52dN1cLvY9jwXJyyE
hDJA9cwutHvHRTDeW7vm5apWCKzXEShSqsAXYHnUAnnsalIgsOmwVt3SpYZ8QGHbZH/IlU4xuqp2
IJS3oGr7vrOHf2oK9Qg7nceQ+RInaJYScXBTINEQs4iSb7raj4Uhgf3gR2jYHKWozpBJnX867CY9
QccSufRb64wmJh5Xt4LYcdx8a5ir2gn+wOpWEdJpWYgJSvJTA/U+jY5ePnkYcRdgV2R4NF129p9R
71KzwLGKe7jnP8iMLNJ1KXTt4N3Jy88ml+6f9gENPq+QDBff+F5RfiEZAS4D/s3CZLmxDOhlPatj
DkvImwV4uWcpihO1JZ8rY0CL4ubmqlyCu8MhrkevXU8z6peOwujdGaCehZaCGnbDRONJXNq/DevE
Lw3W9Kl7LZ/KQ6AI2Ey3goHHUlWwm8TC/KC3rteClGf3azEbcmz7BQnz3xrurkWKiLwxxoyBqUVo
+Lb3wEyDxF5INhI4YwcRdFPPzsgMt4BghqtafH0qr6W3XQC7OczVmeu+pOcwGrH8UwgbBiyvjAHC
dvBR7pNMW7JAOIL0l6PLXqN6rRwaDLa5uG0TGoZsStUBhJGfyhED9iGNKYvDHzBXEIUiMP5vXX2W
3W/+TQ9H/FPXsgum1zhaIyVh1MFzoFdPrwmQ8ifJIicUNJXJZdBSERsraBGMsw+7Vmaweb4Xm7ft
H32PAxM9At93hs4u6EzlhDX+kuUXJI0RVC6+Dutw1DqKZ8qAcoJffE6evLEbkz0Y93AR32JXgzrF
JNLC9naBH5XjaNcxxxmzBwZ7ApEdP0XRLNESlT6zDVAJi2a3nHfmOvc5pA/rvp48CJNCu7qfZrF4
I9aqxrRItvEESMLbQsXFzP40vWKkDugrPZUC/vL+o/Mxat4bmgXTm+Eetb/oOi5WGb+xgyeBael1
hCvfDpiip6/wp+eIRFnrXJpOe6NsF4ayaxfh2+UAKMvtqCLWZvzOBvJFlHJIFmoeXWMdZbhK8hKV
xcioqTm521ouP1SLf60SDBEXwW35smtPyqfb5Vq0s1ACvQva+bmgVxNLuwWX5L9iPdGeYdsY9+Zt
+4A4jMBvLaJjG64UUFboZ7MkTFrWUzCUOdsq/CxaKzBhlmmbluuxGBIBxcpPcIeyIiahV58QX4O2
yA6wFNr9Kge+F4XYIIkSxgJyKiChw1awF0txBPO6tdtMN1NmjSSgukSwUIkchgWnpw3mqGmcSE1B
ke+aMksY7HDsKJyNkG6eOtNpodi963xMdy+o5QVmdEwpHz6oCFcemdL/wuRhjgTG9dy4mg1KowdQ
Qa5NNkGJnqLJEzTNIKX8C43PaSGD9PnzeEtNV4RhR/l8+mWtwYHX+VVxededy8w/xAoBnokhoD25
54Fbr/ustvjeusdfxraA42W8eHGVNPLUp+L5No/Y014kW0sfHqH54E2YgTvtOYczUTvrftZZhQuA
YgpferQGxqdg+lL9RhP+H8XCITkQN9roEb529ixVbIMXzfdE+h5MF5o5U93upeW3iMWPP85upUPo
xYg/elh2BBaQyK8fT4Cszyx5PXASdTSXwilVBWwxJoBBJ8MrzlbRUZT37tpLIuK6t+0ENQMGYRYi
Zg2kBuNP24QpJaIZt7ygrX45L8GrxihCgRVajCqNBzoTI5SGQElfiNEqeCroZfJ3ZXJqE6JFkt/6
AexW5gcy4ROnImHfet4N9jWjY0tnTs5oQvUcHEeRsVRPI5h7EF9xTFNkHVofPWwpzIwL51/dNkKq
up/wnwSFEDq7G5ookJ8jM74oLRf7Xxmw1h6u9torVhvYgEZMtVeNSGZTJ9j3S9jUeucG9i/I0vgv
Yh4lI1+2bVIOJxuES7yL9E7L5S/Ket5SpuMRQcKAdIaG7JqPQSlPV8dXA05HTSy7ZGWQFJbxPl/Q
KEmVM5qlbYVI/oM2+8rXcRcVhguJ0pAeCf13W2+H7OKeB8cqVXj7GGj8m0qlctDtpigG39HzVbo0
eHAIQ9hgFXpBUjW5KHpSoKhjJ0tC4kflk9Pi4/tATuPMyx8w3K8UPlK7jVTEAAAmvF56hTFEV8Fs
uGy41xtSRsWwRXY9rOBMBg4xTbSqysINMrxJ1hVbglZjNS33mxE5gpcdXHhYS7q8ueTzQjDyfA+7
12I9yb10f0fEAzMH7f8rF5xfNxz1w4nLcBKiku13dM6opD6O1IVry045w/zYi8hKGpJe7pE4sOJk
hPrPkN9Lhzd+52FpA8RrhpbZ3cl+e290pcZCFnmou6sppdd7Uyod3mG8HxQMSD3WsJNcpivdKPkh
Q6nP8jNuITKn6aYY6RoP59snLSh4ZZkH1O9LwhHNKsAsYN8/8+GEl+RP6HwRYBoSQ+ZvJMXZzG3R
tfeSAUJ4GbRt3VwZ6d9SLC122YM3NkMbGJsXH9YG457Y9LztLfBjmuE6S44LwS3ejvhZq/D3viEv
jqi2LhpFGA8yEJ38PTcYSTAjwPViEEpnXMhVP/t0RQfY5OFejTdi7XWPZVARJ9fJMgmrn1wvEtkh
1L3xtGwtkOp5IIPEDixeium82wUabYR5uq+MjafVJwTQ3CkPDCKdm/bIxadpgg6Nn8Z7eR4FDzVS
qFk17DFrJmz/eiPUFtxDuYnmrKsPUp/tXL61ObOscSM1vooZgoUSLJ8W2kaMDAFOXdMMJnEUTbaV
aKe4cSU+AHAb3DgFgFQMoW9O1SknRJV8co1vHeCtmOovKgGwQad/yl7m5UufDoEvWXWQ9+tBQdvh
4jpXVYC10SYdEw0pCD+OlVzh5MWGpFyC9OYb/mNHI53UdN85fpt959A54zg9i1/MGOlh89v91dDR
3ESxf3mEhwTntJMNynxjnkizTkLxdcQYSeXmI/d7wt5NvQC9V/uuHXQeCcyqiP7xpcWqI5XzAb/P
T0754GOs7X+aDZ1zt9kyHX7xKU1B6L+nZuZIAjkvzwfU7PXN35WBFaNTNzvD2JJXq4+bbDcHdhY4
2GdHAZVzPn5lIFkt/3ZN3smqxwRnGqrCK3yfWzy05YLSsJWkbv6yzoh0vanfuKeNtFhQN7kB1dq7
aBlBKtX4Vli5E6lrHm9CQCS/OJ0yLFgjkGQ97nsmKEC981R4gyv+mCM4cGEfNsFyIJGkQwk1Z4jF
Ene//KTQ6/qb7LdzIa2KwQ3jyLmU89Uix3UR5Yt+5UX/pfqWwTSdxouwm8J8FNd6fnlBZsafvF09
7NWwsGmMGofA8J0dW6bOL8frd6DxkPvtr1r3s+KX807mfU0y7UiClMOhxjT9Gh+D+sgqBxJvKdxK
le7GQTGRUZRgF+IfhXXPCAHbh5d6r8aO/Bx0EHz6X9+SRZq6Cw86OPwhauKH3kS6fWmL25ecQ424
FEaGfe0Cd5+GRKEEGKqXE2XT3WULyhcMcBIddph42gFfLf2IQSOtvCDkQgu9FmvTnnyym+KEAuXj
AolMUymtSUJC8axJkNBmST0sCMTViH/dwQ5Gdz5ToBMlm05Ks+ApO0VGLqWp2w226FuyDbzHDJvQ
FypDh6Vtp7DK9wfpfduh/Xyo2WzhW7XCTKpjJgD/nJ2zLq2g52GGrT04puCjOBmxX5zzX0rYmka4
x/+ieJTOfOgvocerfb5y7xR/7nM0j0y5lGi1mQ78aNBnoMWw6QirwAqpRoppZ7yJ51GpIKazATjD
z2FtvXF0RlqlxSPGlWKsjHschFr2taryUeccifhhvEbX0OAaK1rp5cdOfO7SCpT3kfVpWawCT6XD
cVmGsoUrd43U9UNJk2PeA2tJCOprCpgofIs5sZ2xVelgLE+k5CG9pX/Gh4DgBavATnmNPlbmXCri
eGTMAp7TzdTXS1c3vMiSPk59CGxToGK0I+3HxcCf7ggs61jayGdnThrOdd5mr18/blzAnjMEqShN
UyIpDiOP9yNFra+1LkBclX+SwugB4fhFNQKobdXCMqTg9a3R4QRpIx9jK6qELU5K2GRU4lmZOwAY
xw4HfFqzzs7ilgSjsrhHuK5F6+FTrIxUkg38VsWt10JtpmmHplYSF6hj/GSiOfwEIEl51BAluLLW
mzYNfJFbZ7o643dz1L5+TqIlfkLMWzTpS8QFy664lAMD6zFXlqDqzROigTNEh7acpeENKvJKami7
OkSe8CjOhDkZzIVASUmLkqSUmTQSqdBvu3GxOMBOGnTXkJ1s7l6R0toG4S5lg4RhIgAzACyVivjd
BN/XduWoygs0/dSg+rQxQLnPRjZs1c5vytvme7FuG9kEfpTHqy60W6KDmg1PGTJNNARGPbIDf0ba
cKfmEHGbEdINo1JrAlIz5ByqjY0HRX9MHbD48SfKCckXrjel4s9IPvGJDOfrpYAjhqThXtW/eJSr
VsCINUE850hV8zZ8JnUsWt8C2BHz5ZJYip77v+cja4hPztYh8OrbPbjJn67Tsm1+ht4JbcPgxQt5
LemtQeL6PPkVFc0nWL0NQkSzAuXFzF/oyOuLyZ8895MXj7YKuaRBOXtI2LFY+KXP9Ex/MAv9sM9T
j156ZqNfa3kIxDEILspyeF257xU78+YJiJiO4T5vJgC/Lm9rbvGqBviiF6CFVcjTTPZ4MEBm0cUX
n0FnDiDQsV6/XEkTH6tmYzp7iaGTZR9d4ukOau70TmqIhpUMI7Of4LbObhqOGW2wZHB6gGXqG9T+
z8cDGo65TTZyrqVQhxEmvmByAZ2UMBM8XJ1lmyV+RLFRnvx3dYRGazHntNVXsyNVONqQKd4+qi3d
TIG/DOiytD0LOTzCI+eCi8F4I5NnXMKGFBuQF8MeiuAfNokjI7CPXA5tQkS8BihAzMqBjERXgX/9
k1umPc36HKZ8LnFMtdI4n9fND8xtaoKWIQ/+bDySKMkirwmAGLbVC4lt1CCTLU/rMpJdBiDnLYOO
T5EorWHHpVy9Q8tApYtBDntKnhRCDj03CjrZKSFqSCZk6UmPrvxsU+prNb5zC7AeGGQplaB5UwPT
wjiBxL5cV8Af6NmmUv4vHDy6iHimOuQkfd7+24DWhhz59hSV2U5bBpKc82Ezebp9MGaIRVVmPXj7
I6NxoNKzStp+OSvgIstP636ttydIpkSFsfO5Ax4pVEsehX9zngz9H+s53JfGlpzw1NxvAEtXIEbn
//g2JvzR/1wDWOhuB62oPZUo3ohyx5W7/uK0zEx/3zwUUhrm08QUGtF4+46fRuzZJ0pKX7xPd9iN
6NMNAxPel3p5/zi3YxeTXAt+BKi9bKhbldDIXKFN9U5DpQ53QX9K3rTScJEDWX9+uOkoU2hX8mqX
LtNt7MJ0OKbA1LK8jNqNhaCZZop0zNcn5nW06OfmXxBdluQCZA+kJZQKHqRycOxrSuaRIhaTIqDG
GENsmiuHOBQm6PUalCCBY2ccjxLL6LbevmA5lWwz6ZZPMbRJ9HzPsTjhR65U1UptUVcd0RdGORyr
eTe1vIN+nMzJChHfSFBKi1hEeIAqFfoae7PvWDR4eO4gcBlOE/C1ey/aHsPB5lVKITliQCQNSM03
RYPlgGvIdQYu5CnfknNSmMK7fR4ZBNvkYd3aFIs4BuOoE5BsMUEsxSTWk6z+Rt1gwvxjf29n43cw
bvyK06ImdTp2UnPL0X6oWgikqtqiCSUL//VuX6DSDKalqu8L2zSPkKvHrjNiM2FMy2tlkopUX+dK
7A4vOvtcCIaiYDwJfy0qDqkzbS1t33W2zdF+YEZZzXYBdh2vBfVVnsybm2j2NoHrr4wQp75p9Rw6
rInjtcpKPCBQMvBur3ZnQMK0NovqpIrg71uqmn65pOoRUTnu7wsxal0mvWs0oFwAYJWXDP1E8V0J
nq1HAZXKd1Vm8m4XR4MRxEOy6IAqgYbtPajbxjKbtxhSwv3GPdYAJoVvBo4jB7Ra8Y4SXHSBgLBG
Higyjx2x+9nzIuqueQLrKDrostZbd0QTNYOvh1iD6f8FLNw6Kj0X80sY7clSVdTyeFnznnfG7N6T
GSRTmxGPO+BE9f2l8Ab8s4MzPnz7efMD/K3Bwl6wxB2DjguHyVJqEzNqahZmhyaILiGCkuUEHa0E
K/LETeDsF1HlJQWBdRLkBQO9klpRJC02RLViQpmUqZ5FhJACdDxPyqZVF76A6yIpuGqZQkZgKuuA
gu0T953rk79AEUrCuiOIRLPwnETUJR82g875ZiNOfPqTW/vTuUE76PWf0FNaG9w19Os/3mDLC+S3
FPhZeIvpF2X/BADFiSugu5vmJa4ZCUVDXPLt+OJfSETw/l4yX60KyAXRq5WJBCvBxfhU9bzxMoot
5DnX12TjWVWHuiVCd2pEySg2iRWwx+aDTNp7JflCaTVTjWeqe4F6ZPBHQFZDTWnCVeyNmVKwFUuj
ypOmInUE5qPCM15f8yyl45/qAv0S0a6vR2s1HcEh6BBSyo74ZLlVGTWcnbtjNoAzmGJyVqZ/lhHs
iBOoNXD41XU4dvszlmzhV5o6rnK0rfunp36Sv4Xnd43L72mGuwU0QQPktznfi8N8Ltw4F5kaudQZ
9Zywz/Y9nOoLSaLXhcsznlwpkeGNbOQ3tFHUBFUVcr9oLhd2S19T1iDGvyeO1X/tZGzth40+simU
tPHAyQ8OAru0yFpp/6K0QuLg4xkP4n9Um0QBjXDoqhLSCyqxme/Jk7DAJl8LLUCiyc1M1BacVHIu
TaauImIInWycgR25kqiOdjehaFEP6sGI5sNAAW2JN9Ekk0In5oG83Wo1g7jTXk+sqvXHffP+f0y0
oRXSdX9hMmaRatc5ht0Pww3784lUMncj+5bsx90jqZO2rcarQVjJ1X18z/HRADjPjyonptjZg2CV
VSzovFIrYV58hqfnE2YpYGA8hWL1U2SamFdJE9g/WFBRkKT0Un+oa74IVhVK4S1cwVCRWwfGKFU3
0HzOAe2UxkS4wCavfEjnhlqJ1X6yymY0+9gH0c7jVYC38LioTG6jPw3cG/+VmaG/4aeGszoK5NKr
hQZXUfnmP4SNM2vGJHCPOequWJMe9/SZqwQShou1KmBNqIJ6fc5xFIP+XXkvXrKrUD/aFDnfbbUH
5AfWuh8obw1U+dcb0PlUdlE7TBLvMlAvnLyRterM3mYkeiZceCXbweB0bt3DoDZP2/Qf7r6Rdj7H
t3dAG6OQGXtCVlDeBTzzvzti3bx96NWxuJWZ6hqURrQCzHkmIycc5FkNs0AMcaekUam6xoAplTjc
mCWSyttZRI2aPxOvdi2iG+h++0nDtpqr6PiQqh8gFTbCMRUbnadEU3Iv2VhW5vTzeRzjq49yxDRr
BBXqkFfvMtT8kUs6Ozvr1On1bmyaEOTHmFRyNhcP8orJRFMVpFna/JpfsQ3VFy1bJLliUCZFFBMM
PZXm62Ez9MDYIc3WzhATnvqwMWK98L48TZMu8sh7cnD3HZpWnqcv/1yYeygHi6jONf/rdEsWxN/0
4DhFhzMwnaXnmB3BHBj2IeOkbJVjRJBcdOdMtfwRSCEd9aAfVZ/KzclozcV2j4BbsflWlvvtkhQz
vkJLyMrimqF5ZCJ1r8PIHeQg+SLkzpuTShNLpZpp3d/JsNk4ah0pKfPQswH42lajNfdj3Xo1vzoT
Scf0Jnxi7XLywxk+toqg2oLtuC9OpSRLtm/5vTK8Ob77xnBGPuSKk3D9TCnxkOp5u1Hsp1HWbcXN
kaTCzVaWRtOJEgfo2COQ96TfHNqLeOpRBXWzp/AC3SLlTfqerSuDYhO/Ot2i27sx3FqWlAwV2ujJ
Y+PFskEkzu9xCRLS8mz222cQ6C/fxIf1eQpaZlT0yIJWbIBaR5BBTtDyqL+gx1f9wNzjSnKPigfu
pF9SKtW77opLXqn8EUb6xiWd7MrrSQD2+bCe9y9S1D6xAvs4aQOfdPu1rmf3VqNsQHVuUKxg6ZGR
Gjky1pyMBucVc4qbVzv51MFDwSKsGjhnTT1HixWQoJHAmM+Ash2UBCCy9WKKJP6wQgdoNPXh67I/
uhZbVgQooDeu3g+vZyTPir6V/PxSlkGQYIV0l3FrLoX/PPgOO7cKPEbxjM08gVJTkrZhTyAqT97H
eQARUn7jSZCGPhAbJrU60ZKBZGNzx4sBjH9Er3sDiTLkiZmmRQelTBkcr5TnlzTATEcK7SH5+3os
LrGViVv4v56bEA+NW0o0h7kzHpkUmWCZodMdz7t/EB0CkAdL8fjDLtxYNMDECiHZdsAjWjUaXKPD
7gKBAwjWxCXvdDL8LFqynYHl4uGsV1J8GEi5dfY0djdgCM5wEU9/NnWPWKcDDBv67qK+/nGcXXRW
ZxUwTyY1BThFclHGQZKDia9vkN5n7oW7IUZU5hweADW/oAghhhe2Yhl5TMcC8Tb6FdbX9nAT3Raf
eHuA30/uy2jGMHWCNmXk6k7c7DthQXUj2PZ1VAqbV/TsXiKTPupBfSlFLXh0jQseff4PjAZVybby
GwKKOkEUuY4Obi4rZFNgWOjHhZ1RZKkl3y9LT3BxKH59oOX2LkXYqVpKM2KlSDxgFlyzgJQeIicW
yB6nY3rSXRQcHeSdlYiRgVP/wTDsWnypraKxZBQ3ae3bVUG2u1K7lXtKhs8vg2Y68QJHAq5YU4FW
1uGgf//yuBY9FERlHAWR73Xt7Dmb3Pr60GrQxaoDSgAH5LRkHKGPUJ/YntoSlDPWQQNapSUnfkb2
04WPxSOG6e7BZr0+dehZAib/4KfGBAlX1/NNKIk8nkUL2TgWuehzQDM67Sw82VCNyJT6/2e0GmZu
9QtFGGmGeV1f9UY+I59E0qJM50ixiwbdpQHRIIahBta85WrnztuC1uoUcDF1peCDLdTg7yAQF40C
j0DL0i7lYmeCgWKFh+AXf5Z+IL18/g1CaBPDjYKQMpIu9ibdA1wtlDrOv2Cedd9c3+4rF88mVFbd
ZY6tPbI66KkGZlVRrQGDV7GUGMNyOMC0A6O4dTPbHbCj4tcWLu2kF49XZT1sswL423oiMRtHDRM/
CBvvQIvEBBmsz7oYxHFBqKCN4hbEWWDPkxRttYa6hcwORrqVs7AoRvKff8YOVtwiioKY+vOLEgQz
9sd0qfoCsY65jwb6RsJ44biVNSzM3M0fpjPwY+2qC+ZYiXeg6sL77bYWOh2GiEaNOb72ezVGak1M
lrwBStiTKlMoqZH8h7XftxJMKpWRqxLSW/kdvQILZfiPZmwBpz+GbdpqOAXMa1AgKgLREbtbu9tt
4BpPmZtJgezF9byijCP2aXsY68aMCLMtIKP23unSs14uYaP5etci/sV1cuZnNQtClYuEoY4yJZXU
KOpzR7bdXHr4i5rC2SAydYdrM2V6hRGzjZsCpbOz0hwe0x+wwfvmZqLL9bDVr78FoJd/YlaC+2I7
fC20P+kwWedDHvMpkNDRf11XkwPvwksXwW0iy/1J9N/vEv6mP0IaJ9Jj2ruiM6V1CtFycKuDCnwd
5K6F7X6E79Ro0+2GEYwTx51dflEQwL450A7HyYsyEdNem7YMjb5mG2CGqxuHWGU/I3R/J5ZA958y
N6kfA/2LcbAsaDx5ndWYhrpVlUgvzxa5qbUdzxw8BKil90PA3YniPB2OJHkCTR2FuSSh70WnppbY
x3WUEqL4XzOarP4rMeSuFDBvZsI2s8HkbAHltOXtBEZIh+iIArF5Euf1E/gw5DzrHsUimqMQO0op
xiOgSMna/fSOM20AFSS9plm6B54i76e84WMx6Ud/RHwacK4BZ7GOP/0Nv1wNkiErbbPXIgCtnX6H
cIyRof+CZQ8wiVYEFTRGyLgHxwpDma1m8I2dUUwFb3Lc6z9zcKVVjKfcqEZnVcAzWEdi6oUpMxm4
K9zj03mUit4kCpcqVEekNaXPLKJuLtnOllYMw8HVYoSaLq9alXThJH7rPbGSafJRp0hVD1iR76i4
Kr5VwacP7V9cNlxRgiTY7KD24YX2ZfSBo2xnsKFZRFrqgU0MUpse7D/hdCHaOcB7RGdRVEBbeY9I
BX+9Q4jZpKVHqIC4OvkPDhJa8b5tfXOshmHko7DzI18vGiRKwIvCb7t9gS30zaHhbARWsqsnyoT0
J6xggNSft9FsHg26i/M9sK7K/3Jag9XZ8xMoS1n4hEfX6pg2APrcQT2uE/Njba7JZuor/7G6IiPI
vdCprcAxjwcX0ChVg4/ChFtpH3Yob55AcAnkD7Md1BJhyRp25AUJiqsdeATiA+L5EpXAxqZU9Pz6
+jS1QkbOMynX3IaAoGq0BzL/XyxuCTvA/ymFeBUIcH+4/5omsnu/OqoWAUrNUuwModeMvXirXdKI
Lm95c4fSCK9qx7OAGiYvvXI06GCDSqLJ1GRUhp6W9tDf+GFLqR+xuAEoQ/4oJTTIBLWHDq+I/suE
WIyAJSBfRwjhT2g7GqpVJL8B7iHFFBKJWDzLxV7lYIbOurYUbAW12iwcm4odg5gmkFhFJ+jUJsWj
iLjtRBBf37f1XTp22MocYJMvderQdRzyAkq5IDefZL5emhoVl+mW04cy2w5KVWWI3nclD4DSX5Bi
T1C872dtPL19WuQ/WoHh/6Cf/IB1bm2kt/ez6GAAtayu6Vveo0JL4lTqCX+VD1a95dJBFLhoa0HU
0WgZAMn6CGuSdP6zNOy/MOwBkabsL18QYmyWV8VO6eospcOWDpZJQL3rMTftbz0H//XMCcAJE1xD
wMPKgWtCjm+qBoVGlK+Kl1ofOFd4hZ6HH4InVEQG+j3MdUpbBWrNpOMYIeo9sZouACzT3hrNZGUG
G4q5xcJs1fmJlq5R4SPqgx90TuRTEliq/rRnpaM5uY2+NR7Ke4cxHp485eyM2QoTX4N0fXCmOjft
HYFnPJWMVz0PtrZ/mHFASRFyg5gikm9VxHtvbS9Sgv/aZbcErP/Yllo04zeJSnyS9j5KuxvJKlX9
cLoBjBX3DXZGwULwthLodR0zY3x2KnbZnEHuux3MQoXjAZxXZO0/8uSDLPnZLakb0p6ZrPFYjOzQ
tzspnxNlJByZBoqNV+kY3NOU1aiBGPrmkTNrFNHhy+LOQMiXZEWadbGXe3fLPwtb4tn5/RLHWaOR
4o2ACRebYjigCtZ20vdaA2ajy3QQrrQ+MsPufRMPRKBjVbukJcj6h9n+99xCw3A9cHUcZRrYtss8
Ihe8KPREVXTV/thOpQOLPP7W2ui7F2IrY7CRnfUF0kNxuJgdpMD8a7SiGsenG0Ni1zRtn0ZS0fOC
StDKJwY8phQYxuUjV9IMEq++oEze7NnEc2ZZWgeiuFfInodyMyL07Fawdvmo/p4eo2J3tLi1czH5
YMKyNoBIXTMF9zFEDYheQOW+Y903kQu5Oyy/20cvHaxKwrsjMADqbyirZtldF6SXBPednwiXb0J4
q0xz/UntFVXhWiL5PLIjwVTLkeJ5LYFsQ+KlJi+GEFGum56VjLXZhvX53BVEEGml+U4u1mYAoHGw
pn8IY14Od/3OW6R+WZ81Rh0cE0sN43HOjTwcG+JtDxsQqHFJp6qjFYCB9Ui+QZb/G2JFEGbQvmdI
IhrAX6uccVC1EC0av264jtAu5lzA9sNvFI/vbCFNtr/MnwC7z5AAS1D8piO2xTxeDF2eRJ+MnPJF
2Kl8U0S2Ty7pP+Rb3gZuN5TGjDeF11goEVUHP3BQaidx3vrCGPoG54y8ESS7hFV+InsORZ42myHv
73TiGOOHs2RjDPVv3g94Ul4dLAXGiNlWMT6t/ohdQf/O92IIrdwoUTfsD0EYLY9Tv2SzvUcywLM8
QpV3fOMH/mzvUrerDdb9YBYdT3c7fUOx6/CD8K8VLHv6R6SKxmUSLG0MVJqCQwvUjswYqLusIlYE
tDsGRYgtCWTQqbI+nruknrQIs4oRrsmgevfBqxpmBj3VXgsJc47oebjoYh46InJXAqInRI48/5Ey
3o4G2x/Nft0MvodiBsPbfc5PyymnQsjD8tGWYDs3fd6ecpGyF0luBsys1qEFL32BVXYl+hycC1/x
T1enjrfL0zFfbqG+T5OXAUqj9wy+d6B0Vnq93TDTpl1/mn/67DHK4UyYc5YNbCP8PR9Z1DsGSWhp
S5yBvOyyDOCC7SHMDmOKV33KkDge9H4/oqIyHOl3MOvlQKM0eznw36kXj8wynnyAJjZqI1T3sl19
uJYf2kMDm0vpPKkDI+xCVNA5Id40KY73DrMwdHNeXD7grmljYPEOAxrrNiBF5DjTNKFXkYQjLDBL
eNF6JbSEpMzNkne3Nypi/VNAHnKYuwQLu1nRVJ7ull5ZboGXOhTMlayD2WWmn0ogkVyn2C+p6QgL
En7xBrV8/X+tvT2sFgyXbKXYxrlRpa/MqAVKYvJz0qktpVKT/uPTO3hdl40yXVV7EkPpgqdyd6fp
LU6i0Yk3cRt4SCGt0ZWC7fNRY4cX7XeozgBsNKqgEhM0Nwwlbcwp9kx+vWTXU8K/tfJlNJFHlWQQ
dZEuB6oeVLbXWRJTArDJdp/AsHbmUaddmQrThjE5lSU5GIOqlhXNEggl/fX7QR9s7CeVLZiZGC7k
lXoT58wXlp2115Dy5hrqXHIt5NU/Gv3lTVMbGVoRjtMCgQZfUtLIV2Mr67FsJR+q3W1v+xDw6ajy
zKqwM0JLhzc+kAD8d2DkhbSMzT+aXEIg+zXnXnrfIWaoFH8Xeu7qGdKHXSksCk90F5nBWQhj0gWv
suR8ohrAo04rxcdoHDalc0ZK07mfYMOInBws/sM4TJzAxr1s/QsvBYkObXXxCGZ2iCGJIDxjSWNd
Uy8qV/dlfOuCCoGA6Iw3czxhA1/7WvXQlrAqTfoY8QzqeUfjcTf0ksJQdLKK4zDgMVc8vjhsiOgx
ykWKjlwI5abFFyiZ4Rf73uyf4zkOwR2sOqXCIOqSRspgwKM52fngzyOTOBF0F6RDWtNNXotIitq3
pKqkshReGzE7zHDT0ANIf9IHF5/dsBikv/zG/+udAGkaYlsZ6GUHA0wZ1YZ5NmiRmiE5tWlgjuR3
XcxyDgTE/iSSxdS5YnF3rHwSOHWoL0gYvbtuyM1AHtBPXkuFrbZw+Gbm0DlpQtM8t0GcnX4rqkP2
wkvoG+hgM81QAYgrHn4KpiwdfVJXB5xkrPqLzA+U+eBSbrYue/rF404rw3W9vU0pvdBsbWm2sXW2
QXqq9D/BXT83++yYzYPOM+Z0CgB71Wlg6Qf3feXaamoXyLkmDFputwtDnyDQDOfxOpCo46n67XGr
xGyQFj25OEuYt75zbBUlrS9EPMgDDL/YCHIge/FnyDhiH0XQJcRmlrKc4epMAK8HAhtVLV4onIW0
CtNFkLFW5la6svL5yYPWbN6LeA1H6LAW7OKGb3Ihj00HdRzHzzgPTTzfetze4FHrl6290iy07EFx
tWW7ygWtzvb4eLUC2FQMJuYR501dbuDWGQWw7m01e0vBFZud6tC3vtrcxeIb6VwrBenkAL4JnmNy
FGy6g/j37Lzf8ouQoFqTSUC/iKXA3HjaMhfbkqCYMasDUUr6maxV176aMDh7Lr44uMMCRv2OKict
kQt3OJOsqx5CIish9VyIF20drVaQhv92WEdgUQG+zuGm2GKiv9h/X0nuDh4wY6USfryJoH9eVGG8
j2AB/KmFxW2mSC/pSjpO1oA6zsOJiQE4743N63ywboALhOXPs/Lq4EPA3E8Ko6rQ9LgvO4qZmkDS
85a4WT8ob358ZdLAnqaWZJkBsfHoJ5/wu0YLCucNUxC+viTLzo8HRnLZzsCp4UDHKLRREEzLR1Or
ltZ7U32Z9Q9M6ES0VJABmTcMBTGgnXz4tqnKN6uGSU772jvjU/XIUMlKiS5vQvsL5XiAg7HNsnrb
N6H24eqf17UTXc93t3V4BVHtCuy4jxR7YdV8lkTkAEns1iK+VcxPpJlY7SHhk7vP7WgHlDGr1ZXT
it/x/StrfYZ4opagHZVq0xHx/Fw7d7RY87Uc8uKD3pYdyDuJtq0WP6i9HmkeRAlFm/JbTaa7VEmI
ZB7q0Fi0TkUJL/mIHWv4Bqd3xVwNvNmeS6D7a9rSDtvZyx3TI/lYkMVakycTzcm8y72pVrpydpIO
Az6tKWFuOlaR4QThXNoV/y+f0IZs3DDEPDKEX7uOPLKv5KtWLGQJU8v0ANEMsKIR8RKCU7idBg9Y
IqULMNA9m35KS/UuhNzlxsWPviPAdgAcsMffrgdO7rLoMf9y5PsGaYeJYtQdqe5ce/LFpkn3xS0A
mJH1zs72HiPGcQ5Peqk7amy+PBYVPiTAxVrqT9jmE8MWucCcjlP1ofmgmfFNuxcUps90Q7VaM4bW
89CGUCHZ5pb0hzTNsQyfVm56zAE/vESnzcS/eHyyrQbHq0x+rYj6pvKxQesABJMw2xGeRixu/mTm
xJj+knRB9OgHKt8aINVDoZvOT4pX1NoXslpVJbOXCrBJqCA7qXpzD+bBluq0km/OpKLru5dbv9/X
IeMI6kD46Wfu8oN/Gp8c9BwOLCntibcmHFjHat3hfBvkfSUP+iLd5cUMAxMH8/jIYPj20L/+LKl2
NFN6QP//8RqRHyJM/xu2qbHYSvgF2EOxM0VkMUl/8BEQTku7mH4tYnw3+nkupTletzRN741znrT3
UVjLgI2b1FFnn0UQwcK0zk3a5Zlt0Sqm4T1vkFO5DWh7/Haw8r14ws6YEOBCHI9EuY+dy/IF0PfH
h04Qp3IGWxQG9/+4rieaXQ81wDKuFjHMUywZxRHriipSl0000V3DdLfUlnJBRpk06A5IkKOQctj9
BgAnhpFwqUfgrVQN+g5xy8u81Wtmx+YpCauoqgW87pDtIPG4XcQwLsvMLwKGlY/KZuwwA+n4j5Xs
LpYJjUl1slISXwce4ZMucrKv0xMkzOQJ9Rc6q44yuj+IrRSW6MAIuExBldaxYB23GaGmqV0kLWju
LpKZDShfc4jo1kxmMcRqrzV8tfxCCbhOxZ/uchQZBNnyw4K0EKb1aAMfiia+QNShFwlyVwVnvk88
6qxmKy2agw/s/xpssx8d6Gkki77NoNnXmFPwv0gTBMl0owXKpEPLMHW+5XQNVchrzidi+Dm1x1JV
g33hCtrC94s1Ov0i0Af0lQMXQe2PXWesM6YaW3djvTEGswmbtRLTfxdgmllXLhzp2lhaW/244FQm
VFKI6Gir89NKGjM2mvWjoT2d7F/6EAqFvzbgnuA/XeBE14t1v0DsYAHUWvA9D+BPjyZlitCcPvIz
wMDdvpa19gtiC1Y54SJFQVDv/l/9C2I2551hCaN9Bma10EIGMYFaZEeXOZRVrKpDjFhdHYUQgNv0
Eo0wH4y+H5bi4CAy81XCU6ZXzHOJ7rmcL1H/JQFtmzSF8ZZjEAGl/Y/JIp9VG89eWDVw1axjs7hW
6G6H3IsgpTyWdg8I9cuELDRs/7owBni9aE/1vHmXmCHruSV6EcTMQtt4tAc+8+m7V8vOyppJkV99
W4hZZa5UfDVOYBO/3ESxaB+wj9qkjucrr/88SwRnnc85zTjZmcLguFw69ERkHZmBv50DoMu9DImh
sNeiucDUBixkV8BWM5J36DSilGsOVs5huTB+DhC+RfnkniCloZFb1LBQRBxhPk6TfLsjWcUApIXV
rNi0zAHglyCGW1DZ8LcqnhuNb2rpDxugfeIXdIMFDHDlznr3z2bbZIKfnOIwViBQN3lK3xl33u9x
UuiHBpPrI2qEhbfjJfHg8v4cLKbq253oJuIYv9eafbKk/KLP1+yzhLmnmWEOYWw5vXRinpUg+5EO
fgIveqN8rQrU7MWrCcYjeJfQiG2LkZUMyaFCQyVD9QgKH1KTvrPv7hTnbI5jKsnIEX2OjpM9DCcr
F1XeoG7Ay/xpFL3ERS6N0uk/qjrxZnOT0G9hoc5FNcejKJxbLE4+3c0gtsWnWFzPz77Jv/S08koU
Sr75UNGbaYUaa735dltwyXTvOEXu0td1acQNVW35S2OVd+K77+ATieNhkgcOKBfI07N+yEMP6zTF
r4yD1GDs/UeO1iY2+uY3lLtZxwQYXW14XWKBNPyowzs/ScVpWbafOSYYGFslTRCbyttP+FlAdeM5
iDtOiSfo0OYZ6JIJeY2xZm2fsz2iF2sOL3FKh07iI3kqqlFB+w8Yo+apG941f3DTWYqe3H4HV5kj
D4Fe/ifU9n//bnGhfgVz8xZx/EoE2s9yvEBRbBZFPTMyoFBY2aj3Y41Z5+YVtJkxawFExNF4exU8
3Kf/HNejfi3cnFM1LoJyB4258H+LJj403M5v433ucEN+oL1uMtKysiVupfF/spyToA+L6/TqEKFh
s4gjUHX+Tp4CwSVhYOMEvPiEn//DaHf/76iEgxZ7vXmRSwTaga0ONM1B0yBVBQZ9+6i+8faxreEv
xLadfXfT/DsiVTrzCBsJoEg/FKexYJRO3lKnzs5lH48mvb0XYQXzDkaqZ68BotWGPrfe6UVRKNiw
xjMb8Hb6YUrSWp2CqTz1p4uPfRZYn42r1YbtN0d5cjuRexXGsg0uPsqrzKrj1JUVNIiOiOrZtiak
BYVtGly4h6eUX41dW0t+bLjExfhB7mIa1xRIL3zPWqN9ybgnFfFv4+2rhzJ2d0fCTTbeGvlpOl1Y
eycFnI5ez8tW7uzxMnx+cBok+5PZadpIaqTi/FI4Gtm8i+bzfH3A1Nn8d7UDV+mjMQ89TBNe2bem
pLsh4iC2gFvcgres3Mh/28+kBN6p4g5BPBoVitE4MEAUDAIeXhNF+LeD8QjRSQoVzltNJZ3sANSj
HvpHIijTsiGNOYra12jY48UkyZx1R00z5ckeVZteuif2kXmXDwZ3qaONmEw665SN2+EnR7i31HdK
AvnQdW30fGMrNWckuKjmnXS7flblm/hdCMmFmrn9H71KnEV41ff1Vu/yG6fKRqPEscHnAgsOL5gl
nWuhIuy9TQEcfUgixFT9nrYit5BMUn3eJuckfN+Q2oN+pL300VH0U2Z7erJTOA5bK4XjJSAvZrMk
5u7JTmcYo8bjHCtZxTxd+KNRX2x0bt7aUoqfj2rgWCb9aaVRnWDroURjbvu8w35KSQf+Bac+ZuzZ
VXp9jl4BA/qCIcD1PELstPkWFTtVOyzUXPKTPR51TQsuBqO9F9oRpw/toREYu9uoOB98FWat2B5V
nt1adWQ+sZhWRXqQuSNMaY1b7BfNefUb4HMma/ELSGEudrrJKPOLg9S1f4IZgALfcITwVmh5xkSK
+oGMEA22xtXRDI6spR0NtTJYo9ETBC5ckTfIytWeAoeMWBurrwmoB9u3NECgLArvqunzy/VqcOxN
HrJMq4Lf8muLdh44OECpjsZ3xvRfSLNZwrs1bZoHecJuol88k79tQF5pfhzoa8Iroog72fsmV3TM
jjuAQVpiVMGY856oZ984jo3vyTdksz1idq65GwlmC50L49lSIGn4lMKdNR4GJ4wOBMgxORksBKyy
UEe1StRfw/elmwjW56yFnkXQF6qSUdczc/rA9QR8iOwemQJjZc7PcAitEBv7pih3XkmDa8y3rJC5
AN6Svc8AKtGcPY4FvSogcvamOksOcRhPWI9AmEXfZsKDsii2lspvU9XlUbPiU+ChR0AROqcMHA7w
VTTqakME0jG6OFTE6oHlKlfG0lpTqq9TJib+0iiXlmFSWzsTvl9snAN8ny76GxL4xy0VrfTjU19A
qwT/14aWv61YDdK10eidJNrwNLMM5INjSGOnE1DOJtg92oFgVz01DEfAJOn3OLrX68L85yPNalRs
Pb8knoayn+1EcYTygh2M/xH0c3esuq7YSSlJByj37EKBORKYzEuUEN/KoKHFEbrEFdSY6IJ1RwUL
wOeHUp3MN8Kb8Hevw8Il20pWN9YpHZ4VnW+NxE7pHGQXkMGB5QZyBa1lTnuht1qknwX93EhKqMt/
O+KYnyK/IHmA8xr67M1Z99VIZVVVBcVazscaDp0Z+V+yRjPUms4tbeL/O/mF6wR6aQmE3OBy7Qsk
0HIkEI2w5gsvEmJ632T6wSe0TF0dkoJUBe1tIc856dbnLVZkzVA8of9LzeQH6NEq4FT+mSq0B3Nu
FBAEDcjPMfKPNM16U3/LfqiZqWzOsvwDY1XB9xbl07KaxQyyOTVD2yfueF8lDF58UYKidpe0mn52
6Fj8OHgrUOl/IBsYr8hi3r6GcQQ8zWzBqaVg3RD1Qx2vW+B0Te/mwPAYd6aIrcSJyXpZcDdQ2cIU
e3UB6tpw3xJZzsX3Y9/cs9Umu35siKvMt55weLXl00dDY3So2mi0KXyi6sG3tPM0c6pADxXSVgDc
S0P9njcnWqwKdJDbCDBXYTDEdlJlyg1ZWhVWxYZgzYqU3XInQdGRMGefhDFeGpSJZVM4m8NvXqi2
MuDHLzlWIi6K+rxkFAZHGpxVE1VI3x8SVxlURFD3YabtmUEohj187Obe1RolbpS7e+4TDemAc73j
j9P5NeVQn5ayk3fp4uCLdh/lQuzaPpFfNYyak3wHeSHfKMejsB1WhYQL1DG3OBJyCOgGUzb2r3IL
mJ7sZebANCMmb02N3tt03Vfn7uq5vxdeuJZMwzz/g9LtINULoghBbujJg2Kyg5U4lAl+MSuOgbSN
9qSwbiN58KY9G8FmBPGzNB4zqv0k1AB8zHP/Pi7HigiTShNY5cI+8foYHRbI+MrBXvxoSIMrwyDX
hL5C9tEgDC38J56KLCw9dETXtoqvWyGyWQFCFvmx/hKqAP98sRLgcyfffm7q1tw7FdD2EeFZclAa
JwZys75R4K5EFktzAspjqkVf3PRQLd0VH1dCM2sAtHz63TVLL/tNHRoR3pJUslk1lq/GYFs9AzlE
rQJiPOjMZm9H108he600+VaYRsD9byyGdD7WpfAwjueTb1mXReP+RkdW9m+tHne4/3IY3KByNalb
tVxTR6CzhhLuiCAsFcd2IBDWZ2K6QgIQMAcWAAkC4/9RWP1kD6hBQIdY9EgSkgVC+Q8ADIuwALmk
+QsWIeKzPelsnzBk0/V0LcL8mrU7sw+YU6dBJMIb9wJswx/icrigM0L46v0emPjkYIcRDQDVL43e
3omxv1HlnPyTbV1jP+ONY3T0OM5lKNyJytgFsG2Clyrdi9A+68I+/9WmBGMZR4zo9sLtZdLlxjvO
xXfYJAodLopPwSG9YkoQ8+tjo3Uzu1nYJM0u1uTW44GutH1H39mYguV5QL7DYIrgKzL3Xz2suKMv
hsHh8woHwlcZXyj3wKltzLC71+u+248ca8lBW+YqYfGJ+VkCZr25V2aLqiZtB7avyTPFVjnqC3YM
c3ib39hmnyL/kcUJkIyVHW3mRE92NVCDsggWM9mIWdqsMMpCUgde1c+jaLjHBJGD18MymCCTqIcE
v8o5HqMTot2ivNUGnqpkLwCoIkmt+8ztE8/6Gn3dmijcQPFY5oPrjD31wTq4qTWot61t/SvkJa+l
fkDAqsBV9+iC1UWC1UvfgedZ+7MjTzkHKHgDJZoXYElVE9Q39xfkF9226Jaq4owqNe1afslXGGPu
bfHqyKfer3PFyYeHd6PtAoc57sJYS0+zgzbJkojed3HSuVok/m+EdCGk+8cF5iNWRo0QV0ABvqW7
SAGPL+nGxp80CU5rC7Ls1xuOAkPPAgEn8iU38gQrmr6gRwEsMph7id8bVbp6zRfGXL6XB0glMGIB
sYtaltq6XUYc39vkoNRlehI1Bj2znsJ1XKIllqeILiDylscV8MqUubAtb3YUcYsm2nG4c6wmYrT/
fk9fLSf/Ridcnm4T16hCokWM858CE6w0czpEDLXoqJKnu5qdLc2y8aRFjr5F+lAv4AMbG9MOIkBd
D67hWt8oAFYDyqRm7l7WyU1UfrbOhzxyuc+g2k8/rbunfs2s+WG3+L0UmJDtemXltBZNGwpluF85
/gpKZmlPQBdKpFTg1eMoEL2cZQroltVdpkZdnFuE9g1n96nnC1CnlILc1h3EyASSzTb7aB8ZzbD9
Q+WEaL3603IFJBIETkYGipJXYZEk9ps7FQMIXy4/te1PBj+0xs/pRgwsAxXF8/nWRaQZJACqIFW3
Do6eWF/rvGiqJ1iuhDD7rmSap4PZlvm2l0QYe6JJKR4DRfpJ9JC/t/Rvz1DxSp8437xfgWQOCZii
RuF9EMfSzzgIpBRHEJlrSVsFwgKjnTW3VmO5jocAAv2lw2dScZ0L22nwyBtzEx2nX4n3zfoDmj+Y
Zx9B9DahcTsorQQ9a2jSoUi4hpeaJGD5EoL41BLd+bniJZ9d/NyMZFpRqBAf/T1BTEFCZaMh+Cmx
W8PAxQjjhtM5cyNnh1LJZrUlVRlTRFsmeRGOb3Avbhu9qH8VSLNPDBE4fsbvkmwYObdnNaBfOPvS
sLqyeitM0Im39UWTRK3O2Jcm7piVn3nBQcFQ7gmEapVEd41FXX9icj0YqQXun/Dxp/wVWs+jW/vq
STvmGos4uoc0dADut1FEoa7WLMCMwxDo2cZDc4FeIAwD6U7JyK0dQ0lck5s5BMSBcQIZhyZL6reT
0l/0FiMnBuFFd0aX8pr/tDKRV8PgsYvXfOIYqyeScsY7OJmL2fuhcnOWxdMvb845wYUbhF8LEwjE
rv7WJj8EtwA0dshWMmDz6frprGt0XFhjPjUS/Ug91qITljGdahH0JkJpXXvZ4uL45y7N77Iq2yRu
wJvbkQBiZLJAe+410nWVQ1z/NREaNlvb4XyCmGdPdkYuQog+6kgCEKbUKLUQGosI4qiob1oycX5D
2orLae4hDFyup9Z1mRfWZNfqpAPPURPMLx523UC5LIZSY6kZYhJLjJ5THi9Q2RGmWJw+AYWAweQP
4hVezPE+gBjstB+ui/E65EskQTvr9mmU6tIYsg16TMnIjWYn5WwAc+k1xB/kQ1jCSBTCWnWNeFl3
HnCngIrPvp+Y5PIW/CkqgWwnaQV0b5CJk34i0Yf7aZQjzI2vXs6BybEJ8NhVci0fYRGAkS/Rm4G2
jtq6AnmgHPSYZzlTr5tgunJMGqCq+hanZPmHgy3xKTSZn13urKpmH8PkaRHCLJNrK1X6geGaEpyR
wRBFnh3E81w31JMVvVfLjktu8ES1rcK2KCm7LaO4sp7VURIFAX220wA3PHeQWxBKVk2SGzFELa2e
AME1J6FpIkp4+iIMDGnIaT8gWnxhxjBFldYQ+dtafRxcCh6xtQEjmb9XNXnpxqszoYpUhmLgLD70
sa7Je6TNXmAHVefbLxaKBEhjRbwPxCBjFnwBWewkYIEmkew/MNUMktlt7kzJdpqWZjllSFM104rI
nz1b2odZbZLmVf/Cq8mt+iJP1TRXajtTL51bIZSrqACxobk0bBrJfHFFt6mI8Z6TUgk34zGMaE4M
2H5wZS6FCF5X5wk0zQ4oV4cXelaCbawl7HFMMvmY3g0UP1l22lcC40Et5YEVn6hLV472IFbg9+yG
C+CEwOlaF5DMjcpW+PjMnbsowMDlRHtVbOdAjmO2RJj0Cbx1zSxpBIKL2xMibrB8OS2pK/PdMcFC
/A3kLK3xv72i1hwmuf+PrPsSTIbxovCMsKdQ3A7WsgLfuU5anQtsnP4rRGl7BcoU6k1wJFIRWSPk
6Oq3CgwIn3wwkdEI2XzwNhKUiR46iD6LvkJL/EB4YcTLGd2NzJA6L0v1BEcocUkvcMbaVqMWzKhT
uUbPUXYRJxXhslWeVzZuUtSJaMtuZftZGj3zJyujkkD1uTePIrqpwKLNah0ZgyCsTdTVaqrs+Nt4
jupsDJpEv1agvImiqaUMmopwxDOCA8tDFOguVH9FtdOljIACOGtrvOQGl8Dd3dN639VJuBRtX5W0
U3Wrp+oqCsv/pTK5WmKOKISuW1fv6BI7rUuLTWEZs8PeZmiMFZty08OMEem8URVTXAGUX3U0K9T4
a5asQWml3GPVsr06faG6e29GU1rR8P/oyHBJSA2dDMsYmMtmuqhDIMPMuqmw7mPQPzCQHTEkmosf
VjpHjpv5y2KPm2EBVQNGZHTML9/92ARd7HMm1tbEq9AXSUwwubyEGZnAK/RkEIf9Qg2mQkZikt29
R9zppJ6ntj9j9dUgSmtzI4FdxGCHSfdkPCna8G0b+6UGS4F5PNSj4BPA1nIyTMuDsrQAwmFJAXaX
NJ3zNZqeSYB+diZH+/tTBqbkhBeRsWFl49rxWzvEecaLisGlvkaqkgAzenAemjkC7JdhuDyCfIji
lrkCYIBsKG5koUXXM4QG4sBT8q0OS3ymdtGf1Tr+mP3LYlAcKgCX6Slph4ZXFy1XlEAEiT4NAXoP
2fXpfyqFVH664gWblpVLovw1vxZFTiXB/a18DS297vqasYxBIPEdpL6t8X0qTjVLdQf8docQbzAn
us5NnOmmNQvvc5yVr7JjYY6kM5yyr/7IzAVnHsuS87AnZ/F93Yg1T3rvRmDoOB99RAXclv8hTPt2
fH2H+b3rv4h7+W6XIHCNhqIxCpUscsw38hnO9CUDSRV6otOK9HkyMS/62H/QqubaW2Vb+w3qyhBF
KU3RxFIw81OvXfsOLIvntrWEofmJJq+UDnHKTNGhr1VgwKuEapXeT53nuoUwvyBvRuuPGfeMT1jH
U7Kq7FYPJwKOBAOdARoUKSddSodpFeYjEH44DjvmQpJ9n6wobTelKtgC5WRRArY7gLV/XNKXrJvB
qG86eu+xkPW+ySAAVPlWMKfF21PUI2ZC9Ts9RuY1MEHPVcknlw85fIFYu81c/nKOPo+9pUVh6bO/
LjkS9G673RyBOClTrFCg1e4rDl2rF5QpJg9hrGTdxYHRA+lytZ1WY2HtU6Kf6dx68F1Dw+fqNI8T
wHUgehA5To8C1BCl4at0Bw6+MCqX82EleT3Db3IqEXW67dD2pP2DhqU7at2NEDRbcH4A1giiUuNc
cpBbyqt9Oo7+ulT3pn4jKk9wttL11RyVf+9ctVmlj97+moM5ZIls+fFt4On3IY9Rc8XyYvRNJWHy
2SbCf8MENAdCR61Yy5WajjIWJCQT3IGi09+Ena9WEiXccxaKp1vlEIqm8eHYahQsqlIeU5q6uj0b
kCb7IBm+39r9zwfT5EFl8qKjHJCDaIvvuCyrmt/YHjDrXf1AHXS1IwIl2iTTqRa/fG7nskXzKjyn
yz8Ve+Yi1XNjCaaYPnzJv92IiifhC4ebjPIwdaL6l2lWSayCdTcNTTEsTSeIaAukZziRf2Akm7bn
TJ8+niV+zMyb1HqEgNHNGqUXT7VV/LWLqYkSYu8vdZciJIOiCAIMGypTnuv89MrZ+XwGMyYuucHh
BNb6ESmbCAsFyCSUu7UXDS9w7ALUMdaN3f/WvFG0MrOfJM6ctej8IAtUmWqz/HtTEJTloUafN0nb
A/Wjj9hs2akICYinnCtYJA9a/Bb21wP0TGYmmb+nT0Q0S7sNZ5HrviFF/32y0gz7vZWOBhVjWyCn
g2plF/GcWlj+AmGgtC8wT4ThLf9v+CdQcd+WAA2nTA8csPiJxi4VDNWe+loFR1P7LJUl6E/r5hZY
IM2G0B47MpNX36yJTBGVXpN5KQpD+8T3cy+5jHodU4EEECUdSOhYyZzTCbD8K0GS4xd/FhmNNAVr
5Hn/yvzP8Su7yzf7vq64g37o6Lgvy7CE+oJQMY3EJQ1djtmAe8VtfY6Gzlymx2gCYmTCoYUlGuei
2EGLbcFJ8fyTjmg14yzj+w+NRJ3kiCCj9K4fgLm/WhTn3Q9UnvfC6r3ga+8yD4jVFm5Sh9CcX5/m
sQxgU3aOOZOZZJDlASTmaT/rQukdPHRacRMfPYhXgtlFh0+IeZErhrK65n1A70OIwNrnGFp/CL20
aLNEtnwLO+VdVdyNWAHiIvmkCYnSyjwAmboACqlU1EDTnEAnzPeJAAci+Qh39ddskIFoom3UxjvE
CjSsSHkF7vb4AmFhIoltoJazk8UzF9tEsVV6RAj7GUOS4hPo4X3nG9wpDB0PCjm0X9NjFsN6A1AL
5TB0Wc09laDsTX/AaHYFVM5RgytcrosaIwH+R0r8iklqrfFRUOKjKfSO0JslpY21K9a2x86OZB/q
FPZsMY2FR//qGB1J7Z7fCWh/Spj9h5gKbnKlr2ABy16NTVhRNy9yL13TEWH/KJzEFLKghF9BV6Tu
TPwGC5iZlz3Sl1SBT/5rAvvgEQckD9Ncf7kDTOtv+qG2E65RsgJybbKDKCPsSZSbXl+UM3gE3zFz
W/j4IgC45JlTyqA2zkVfBzmk3HrhES1tzBrnJdmXz26ZzeZvUxXpt4iZLtcU2myi466aZZw2WYjg
RGcntoaPlvg8NLxW7nvPf1Q1QQ6002q2GmmVdoZYisO6q8UYu572xV4qjRhX84usoJ9t+A46zVIN
Zx/UmlKsbj8LK/LPLNWLMIBNQjyWNFXoKPW1LbYAGTgmTsdUqKNffvw36Qe73cV+CUCXvi/8ili8
w1iuyZ2UU5vW6PdBdgZNVmoWI/EKqUGlaHGVzeBIr2ZpdVO3ixyiXxvtbo9CqpiIoQtif+HO/OYh
oe758f+Wub9iUe/MvEOx8zIdqKwHbsBzwDb4VP2pI8ELDbwgKHe2BaY2ACeXlfcjj466rkBTOKJD
cf4Hfh6Ula+QPWUFr9hjF51tI8lWiiE1dl4HNVupHFGK2MvkKnZZb9gU9sc3CuanSggf34QtXN2J
pKHgErv7Wvz6fKPTw7GpXRnQe5hzB9shsEFeO1r+38nnfa+y24I+YjF8C3SjdynnE+ixJtKQanjG
mydPwvkgOQYTlimHvcVfrw0N07b7xnidbNz0Ut5vmW0yrPSN2DElvEXszZlJgC4W9LKLtVzUVNcN
DzyOw1mjToOaulnXG0msLuz2KMgLB0NX90Loo+T0qxd9iOJ82Ec8I3sNk+Zv4XP6MAPbBirOwLFT
c2XHEbyjt/w/MY+Qq2V1M+tiqpEDKf36HbYQCAuGBcVqJbQn3ZxxG+ALzLeKxxc0Dj2xxDGpfN+I
BfYxACEahzvtUQu8lf2mzSJ43pxNftTKBlgkSGx+nDJzgEU4n+hKvDqoq7oP2T+CVj5afmgndmso
HNbkt0UDrMCJz46WnvCO0xkb7Ws1jmHuc1V5SbI2t+sb6nhLjNWfQ5DZNTDmkAj3svr8/NXV4WtS
Yxk3oLTma9ifBhq8ZXGq/gHIs1u4eSk3JADrrTTL9el3MlkTYW8F8ze49oVjO5QjdsRWW7JDBYNN
Cd+Cjx5jXndL6M1fvGRqDBXRru5fs1DJ3lq090mqIbv8ToDtmQZlabDr6wnBbPs4jgJ7+WQc55Ql
IPfo68V6kaCgPFuIeKNMK3+WEQkxwWsvVrOdxKzuMlij+q2X1mwehlBVc8avSV7bQzq+qcXLCTpW
jf5Gut3Gm6Om5iGpfJX891oROciS+UL3hTbIazwzTVS2BYyp/eDPpNd2oXhMRepWJKJdS+5wLeVf
UrD4WhjlJqb+jN8YAJFQBGRubR41r99Sc3zChPWh2QlrVmjRQygq59oumTbxSP0qdIHZkm4x5otY
TafeNfvKVX0yK7f81CAny5C2UbV6bUveIA5E+C0PQcTneaE8HKMxlLL0ZBGLxYUDUn4Qqfpt9PuN
+/3woi26gK2pVpVey/U9VSX0+X5XGY9SQLqebb8uoxJz742BLEHevsM780YzDht4HbDuTqLvj1BM
8/evt1dV6wVMXsBvTeEECXSw3X+On2LjP+N69czyMUM+oikPfGWA4BBZH//IsbTxVmIWehfHhiew
4c6lGj6BPzN5PT6Rp9gORmLccb0P10G9LLtfmoZg1CNkX+ugW9ultfDu2m/wUey9aWmFG2bQ6KCx
SyLZDhYWqPUzzD9zvRacqbVH24rnE38edYrpeKjJMADyNY/sb9bIWj9RnyFPYU2/yFUyaPIp7QhN
mSqOvhecSSFl/3wviLJLJ3r/LPBQ8dt5lIsFi5sl1zhoR9MIiIZDGKSohaAc28MzlQjgwB3GcIS5
cJ1F1csdPpoI3Mc6yLzIWrSsWWMrxR2s/eaT8LAWJqLSAqUxBr+38rtwQIWdKl6xkrtplnQT0u25
6EgY8PcM/X19ur8nq9Pjbb+zOiZxX14jNTC7NkxOOTZCv84Vu/BDAkDq452lCjG1Acz8trKymYMX
D0xVSsTSkK1HEofbZMiJa5kmLikFWq/kU+AmxeyyL6fRTGHl6yPojQGom+hYS+r4pkenk45XYqG/
K//blBtWNw+osJCrwZvnFRSkVqJC9UYNKWQ5CWQHT1vivGl6nUbix9LbaX4kJBqSWbZ3PI8NISqt
FracIg9k5gb+0DPNHQ10v1xKWI9oklyYRTwrJhxzqe9cfakmmjpmliB+4MLKmwM/FjtLRs7yb9sl
H1Kd/iC2bKJrXtJXHi3Fg9DXyEwmTPKvXxvA6dYMHHItzBLNZi4s1G58PhpYMYjGRv+uWXaxFNQU
DsGoMNN6L8ap2omMqjdltqbHjJ2nvAtGvIguFP14X5eMjR4jDcnyMjUxSDCSd1V+D+nzsc7HgsNr
NlurTziCwl4Zrv5MK5O6owGHETpjozu90KSza04CH3cY6fV83sg2+kZ43UKrWdKkRqXVhsF9cYUT
2HMi09nBkBNBuo//tL2wIgIB/YGdDufuaJSH0OUni8F4Iem3B+hKjOhljAA9/2uem/MDXz+aoLgV
Rij2pNqGWHUlb0OZjK67NC+dJLv9jEx57lXb0v6eReVfubELgmm4cCtyke2f3NPinlilSb4MVJ0+
iTSvxRs0oFHMQS5xxUYiFeEcOQL+Upo0x8irrjaffwt+pgwtUH91awBXh7vV92k0Z0hrf8mkJzkH
1cIRWUBOs7wl9jv86jsK2h32iRQOD4EcFjVa7a+z+2p18A9ExPMIU0HaJzvOh9fZv6dMQA8VzWlY
uTZ2YjlPEGUifB+qSce841eMaa8yRSHtPhzO/lO0QsBd58JGyQ8HwLHT3hr0RcspN3u97jk+0EMF
2jt2pAi4vzdkTrxyg8bE0WShVj9Fl3GBxubBU+oaoax+fpJOiQaCkAkq5evaiAWcqUP1vS/hExAw
7sQBnAu5n1CM0sViaz/VqH333Iyz5oHXGHx/12cb/F4sNHTGJdKqo2nXAXIpoRSDXbwzs5i4GzS6
9ifSVmMNIJErvUhtX+eWI3yi3x60AYbXQLHPXCHuatD16u4k7J9pEvBM1fUsFJ8xKiF11ddNBlRs
bGMkJa0ri+HfhQpzPKPQBQe5YfQ470pIRreDtbrL1ZuYsTu4rb6OPllRscRshROTA6eSRcYdCZue
nNeVmCW3b8649Sc8PRxx7g60Fr7zJjYEid72nNORqHdPQiq8nLhVuz1fk3nJXA1/rx7qygEE7RNT
wwJles/ZkQpxpdvS9p889MxS2pZZ/MejuboJQCzQYwdH55uta0p82/+fRT8sPZMnABPkowT9XU0K
Z2ofES6CecMKHIPkCgU7CdlJVB5CZ6GryQ5pYc2zXYoFSyLA2NDldhYPWmEZodlH3aeCnXXWk84s
JQ5LbvPP0d93H3AEKDlmDz+F/3eNUQRN9qQRW1Jen4O31qSxBtiHN+Kd0UOkoXNXNlRK7MTQIu/S
Eo5DOLmdost5+yUvPUeWEojB0ROMn75wPxP6OYRPNc9a54K5hVFFifQ/1eGforh9zSyHF5maTOnK
er8+05P1YSP1flwM69Z7drcFr0qBQuvs4fQkSRyDh7jzN8ehj+DlMm2qjdRLzIjZ0MRhBdU1c/fP
r2lIeDh1mCrcnwveusV3xJRDMwDxhKKnrKFs3wV2j7VeX4HDaHT+Whf38OmvG5Eq9U2m89PCUhNG
3ijYBg+BXmMzHMF72gTJYSMRH+G/JtIgozVmgOsP+u6hD/kqmDlp0mzh9+hR9lnsFpm/+ez5qkT9
UqQCPtJG9JjfYqBhtNMHzYYfcnWc6S9jSVuqRGi5GV8gVP2ue4YHcYcp3n/JUWktkYK/4DIacamy
0qR/GhFC/jXkEbtFQX8zNDBVWXQY4DU03w6GiS6/p4Q4UuVaJe0y5NshfPY/6xeH8mwAvo6+pDRf
fJFJ7PnP6IQLTTAF77GT0NDEy3jwR9xAv968RJALrBpW0Xp9aBT73X0KoaBU4a2gqmcUGtMsGfHN
23Qe5WvyNVXYUaHiBsFevcLSUpUgJ9XW6bbHDJOEzVsN5rAaUWX49CwtUkaC3N9pAL7WctSv7xrP
LJAYTO62LfpzJepUgu2VFs0O7NI5FcFn0bYXoqQkLbuI5hvtbkzUA24tHLQvIIhqT+AFBLCN9MuP
Wk8kAruwCCVQOTJHVc2NCMwhO7X+Wpe+ctJlqKzCEJBteXlwW1U+8lEkGXwUCfSH1j5m8x6xl+5d
Cdf7ALsE0Qrjm+Y2IW0Pv1pWaQc4+M/pdc0/3md2f+kd+TjpyFsIQ8CjrkkHVh2IBhTsSNGZ3Tfk
oIrYLg514ltWvPM6b/kcnwL+oCP7+TBoJ8NIGQEyPAAY9qgxqVa1l83SHIVeA8mv2Y649CBP19HL
vL6bSf+O/0JEEkpAGsLjhRYHsKSKtrTOj8DFwWRB9tj/hJB1ay0sU9Ta0733xiX82shTHCUCc7R1
qEJU8HpnhPK3yfA+R540gICjCWu+lPigwn06KjLkosMvcYfAwL8GvyXpr/POC3j87aajKY31si65
Q1VdC59CVRpcDDRdQJcrsXrSl3TCt7KPaHc16T0/HT7KOfl+UexJg5OZWTCFLwTw+Na4ovgnkpQZ
rRrI+e/PCC2R4taog3GeEa+PhhvqAKJObuCDZEpKEfehm3XqpWmvtxsouKcJdD+B8m9tEUhISiHa
CiW7J89xR4UlU3+LCe5EbzburhKT0KyDlxmMKmQp/7GbuTUvyPHltDLabmX+sx0fObkaeNV2OPxt
n1URWD1JpJiF3xQ12i2rKKRPEm4zTNAxIiySXm0xFkEYywfzgugYiQPqUaKBfIM1YXAHAVKD29+J
6K+32K4zGtAt8bKA2IwL5gbSt6zGMu4US3kv8YLN/eGJriUAAtxWxp1/BrYhFvzIPUft8hbQICj/
QmZ8ia/+zCPvLUd4sIJvS8cnBbMVsnirLSRTfuh8I33kJX3R61CRYhV4B/FZu40mF4p2s8MYXWCk
KbVSAoTRLBgIiw45aO6/7QE1b6YUW+SxXAHSMT+z6eqHfuzeNzWSlk2tDyM6wFCS3ngbOycPGk2t
m7ABdVrtX8dYuCgOc4T3v4FbSp98F/6EQ0uZl1HXTlvOkgDKTgVlsOln/ePtlRtFBHdc22DKp5wP
IuvFXSN0X0ly8/dwY1ydjBZ0/k709MTRbndpwLigYoTA+X9d/rooQIGEelwAlWeujZ+ZSs9sJ7xd
08UUKEmbU7InSIUw+3vPVonvFGzu7nJV3JgDO0L0U4TNdORrNxEze/YqKecj8YXo2NjWQIIJBOA8
4lKDT+SNIB3gvL3LNcGx85Ar2kuJO5auaCAF41wdLYZO04o2KJQzRiLYT5gQU4zwG9vHfJ1IKYlz
GnHacyhyPWGVGdCEmCKJZGhdLLw6vtApGS/2dWExV+NHYiMMuQBi3XB50VS0QEoIjlQ44EJwl5op
FNflWi1LW0wBGBBAK9CWpaj8ZlNkAt+M6tSl9EGlSzsIn20Dl8iwZrH4UeLwXub1Jlf8ntvnHzv5
bbq4b4RZQ7UbasQYSdqyEcbstKg+03qVYKLy0k30Zb0mpWcb8Yg2oG1NRDy+dzomQAjbeq/xaq1j
JXKuC+CXwlD8g9a4qXK6RhG2196qVEzW88KAJePAlB30bC+8CTZilNrJ2OzwkM1ssWvGqLp3Drpj
3t/GTSPm8z++gMBKvxAlNudIvm0kZQSS0O9ygFYDzmjek+bVovqNO8vRX+b84LeB4Lq9kf33Kb1B
KIH1ZqSuZ1PAjzqKpJ8rJKEaZ4TJgetzCZPG8dUWStoNRLllBkyqBK9Jx6GGeOoEZ9sclWVYDbci
RI3aSRECyBF2UyUPgN79ZyV1UPUrtLaN2Jf++GoYI01HcFxAZiauvqDuudQlyB9/NBGLOiaHFeBw
Yxs5cpdCD3P+fTj1K0XwnROTlYe8PGh9z9FymYLfRAPn6xzS30L1jTjJ+OHexD1MF5UCkcR/8Hd5
58jOtNP7oaN7FImu1Po/+TGXgepNdVjpnctzRu3NuNDSdK8ahJgVW+FTjJiomSfI0cJk9KSkX9/7
7nDNlBjpwbh+X/sWjCt7hheHL/+XIUi4sRZ3a46Z3GrgEud73g15kuAI0Gt4pLRFlkvcRgD5TaW6
WlC5JzJ0PFQiN+oG95UNhvoJBBrI9jEbl2/wNtNcAXa78CsyReWIjzaoU08HJAz7YDXlN/8rVY0C
AWhkNe59xH88GX4Y0UwTPj1Sw8DiGbfyld1SvsWIzeTtN0BuroQoURJ5L7UOMd3a5VGJd1ChauGO
hnvYhvhpd3BjizcXsrXrrwv38ynLy0KKInH0QXunMPZcz3Fa4MEwjWbPRUKmoGNfy1bqBa+Jt+0m
4CFn/AjeoDsisYZvbVcGBhU+53QT93JAohWfN7KVAoy2KOuLJwbQWaCwhm/cRQY26zAjZknwN1fO
rkG/8y2gM8AvirBmREOhbM/LMxPZ1MEDoc5LZEbV8MwGLGrVz12UaASgM06TDb4nSGk6NgasUixX
LkGZgUhiAtuIrzDT8eOKYogedAdrf3IvwJag+kxsrYYb5ZjiwhfygDcwhuN4l9BrL3wwIIhMUeGl
/TxaglTXb54Ar/5AXlyW3rKh4CrpNOeWM8835BieWP9nXuIzLb1YRgj39Nm7rf+7STZ2J8GIn1XN
swxZ3JXEx4MrPlW/HTqkfXd+0IwlPBbyAKSlMs4lWjlA/UM0gBGTsdyMEUceGJ7i5gJD98888Th8
q/C3llZnrbBUbM4xRI1uAjbmcemHhKssUbpUjaf7ZmwF24yVLyU4T00tytSAYSc9makRlQBUoNVd
eXeELcpQPCsDuOoSBR6J3JbBtPppZKS3s2ST7hZLQGQuH5Adkh6v9XPSB66han0QiukbxEl6ElKG
cjt4TwbDBYL+XYgz/Yxo/XXdZylxuX8oX0r2yg38Dl+2qt9xjvntNW+HZ2blsXuiOQDmQQixeG3x
7R/BP36XjFNrypb+gvVwqQVmK4z3NTlPg8nXg1LcVd1xNxuqS/jP9c8BxAHWwyOBQgydKf7YxOxD
TkeHIMf/wFRiOusnqkAGO2EQbNEOZpel3QGF4BIx7h0JhQM7B4JzygH328xRzAlt/Wkn7EghjB6f
dP0b5WQCLq4iqq2TRxjqAtJadg4bOMJsuJtdekW+rB+JavTReJTkkQeT6oDxCDE5v3N2x3t33ctj
oS9pVv0QxIIeZ+dYGA07LkqunWUVdOn1MarqW5CdMP5ZyZggojHIMLYcn4sdq2JLYMY+kNkwDxQh
0lLXoS/Fi1UlU2A87K7lTaS+nG7cceDikv8LsW5WrY6VBGFhbyowMdnegN9nmi9rXrQXQXiDn5RZ
87jDzAlTggPKqIns9ysHFUi1RHraqdZdaa+Jiya3364Tq5GYHHc5cE3vufeMm+a4VuQ+gOI1nEVl
Z3NAfjzjTdtH9GdpSzIQSAptTYGoTVgkVzFOfYXp5/Mxir7A+hwgA5fv0V7OVXLuAn9lTbS9WLFH
kaFgCJwq7hHt8UPNaa7nQlkVYbiYN2VILOu7MEKSOIZ/BFV55SFND18n06gxE5NWmvLExDFClRO4
StMW1gB7wOX/BITRlw+xIL9/R5zSJgBWCD20wJTVdXf/3jwKaM/uRjhqDshO/dw+w6jI6/rPwVGq
qCcSh3J7eZMfszsnwFIVdFDJq4moG5koViota8rSLjVMBdp40GNiMd7ZIcuaIvorZh4dwcwji7SB
5X37hERJ3olVllmZNjpSwqGMdGvh1/hzlPmJfxl4taCNtrU8yclU+t0Qt9TDU4unsTJD1oPfCTcV
Nu4z79oX28jnPpfbjXs5ZyPx+cm3JjxsG6zKoDJR4fwsRbCtNP0NR1XNVFzWDN0GZs+B7VgWWE9L
Y0pXvCYWnf3jfWL13o3cKm5mvlHUcM7mlWbx1xRdox43EWWHhKwibXOZ8YC4fNn3rRLJQkeRwx6O
6gVkM2CLpzvSn2a5ADRw2EfBujqaqfynja8ReIv2jlVkJupcBOWgYizB63MKWRK/MXNKUWQ8pyVe
QdU1YeBfFK+vtuOgCMFFA/c2oVuwEfoKgFi6f2QIo2vRKcc2Vb+qdl/OlfKZSjHoodidlqFyJqBB
xh728UFlkaieCENdd5JeElsJtC6vrux1rmO+ftRWd7eVjSblvEbZbY6SHuqghAlvMkR2TvBWkaiG
ZGy8fKFAuL0M8vcDCLPzjWMiQD/5xHTXZQ09D4uTqZ67r8XaOlquZY4cvjsD+L61F36Q+JiLn17f
xLKORfcyx51UPzBfcqWKKvCOo/zrugv/9MEc5lxU7Yste/L1Boj3zo8uh+LL0CKu2a8DQCnZQD4o
gEZ5Zfk9V04yjgjuWd+/zqbeTcNi13H/eAcQFFO17Ezn1b+uOqI4NfuqDr6mBJ6xeC/0bU43lg4v
Htxsopv5QepqxrFZBCQqui6roj9YIoaTHdSiITy0uuZxFORkI1/zPwUJWvAVDv7By4zyx0VlJuI1
8iHggitvaNLYp8jyZv0QOwPr0ZrRd3wGEb1uX+r+bWdTYhelOtPA4zAz/rU6ZRXjchZ1ljTKViRv
RxPDfIPpj0uSecL3hacbeXm4uoSVVdqjoID8VMbN+izRzkumj9pG2ZxEoyx3K68wV1CblTMjvoih
StU4T8v6c1Tg6b9JTZ2839aoCUOHFoxNe+ykD+EpH7zHtZXrZLu2ZUXm4n27IOb3iwXETJ/VJsc9
U4P76jZXV2rK8+AfhGsJ7n0/xUvzzecsa3w+VUs4MVosV+KZ7B6us0cbCJX4VJ3IpmUsD3BN4rtI
pcGH6XC+qAvRSRCSY5mCShew1ZrIP6we35U0VtriijZI84fu13OiclxZYz6ZqpUK34pGKLVTwzAP
l+famGFXI0yDKM0eioCTr5sMHYsrDnoOkNNfPDP22cQUjqSutKV1GCZcVHJu+GZSc6UDiJ/D8MjI
HXQdDMDA+RR9WCQPgoUSHVUuHVgFCMPGmNNJiv/byU/NpZuSan5TWzlEzPDfPMVvSBi6qwBaBRk9
5JQ8TLzsou/7BMoYCncsaic9T4dFESR71galdNjiQetlDg4NjAt80W3iSCjG/wDfSc0HEeikGczL
52gn8Zhl8QOtihuYxAbtfWec5MYtuj9OU6gx8n78ghcifruneLJm8Hj6yB/Yx8BTh63ge9ctf0AG
5BiMhvpsLtXQRcpnCTGmHliz2d2GP/YBVXUWPYfIz1eYoG49I/mT31VDOKxkavDfM/+Se3IdRSQS
Ks543BxDM0Q6tAiq0FlgWv+eQcVvnqgB6w+yztw69KJMvFMOPdQAxdjQzlfZH8C1yiu8a8JSx4/3
5217Q6+fn8mqNeTw8tDa9HST90BEKC0S7tZAUexBd9OX/YKydKBCTyzABr1eRSDSHk9NfOwcbQPQ
d8aus5UDvQd8CaFcHPgcy4y5BVQTA96ttQKB1kNGtbsn9lNdx1IdjkqpeXlnXJiRlbtrgAJwyBf3
x8Ph4IbxE4JFLJfFIh7dp6PifB6ZjQ4aZ5eBpLDI/e4iwCDIsphgVEiJZjsANj1hW0x4gRupMz/2
V0ooZhctWH9lHpHzRh5WfFJn6DW37abc31fCcuDO7hez1byPtb8jzx7347oL0062RGCciy7frHUR
bWfSazubAslPUB5rzkyMhtdQESp1EGJXi00k42kiUxFYstEACPbcr9WevmRMGtCO1GHK47oO4gPF
emAns8lPjozwDTUYeCfMmNSGMQ9+dX5Sr5cchaE8y0pEgZO33OdYKDlu6ZGgXBoYMt6nZw5mQ1ji
Oqxn4Lln7Nf1gz7eKVsT457wC4GFCPot7tv2cxgtPZeHOU7WPjBuzw9PgaEVnyw2EZixLIujXYgT
tiV0N4E6WijAu23CEGbth09pgPYWhqGd1L24nHDinN92AYJObFbPkRwHd7a5MZjobijWRuMuYccK
8A8TCIOvkUbbzSlvit9AX9gvVRzzD6nI2PlEtyz6/gYf1afUwRCmn2f240ZtlkosTYp466mSRxor
nsMd2CgDAjc1Wwoy/+92x2Y6v06mv+jQo5NFVaGyNrRi3pBmuzdhN5dxKXKWstNb8Q2j1B4u79vc
+b/m2PB5rC0UWJzFQ/Eqta6vyBFwfdhycMUHIufVlzYAnZPHLWuyIlh4lspVGC6YehKVZxFds8zn
CPoTpx0Oq+Ah3X0YAaXLam3nxAdeTYLoFMoiv3rHNVlrkvnFN8RqnJcC+hTgHjYnpqObxUhdhSWK
ycYFkYycmLTwg1dk1f/nW0RDUQ+DqTGpr+17VAr7ZD7zwSa1KYyJdV4WmvwA5IttH1rBeZeeSE5+
qSZvo9Eb6tUh19htAw2S0x7Dcs2pERYoB72+QdeVtkFVf71ynhCqQcQR711n1/+FXJYyON7e5Tk3
EVjK7ukFSkpfkAYzxhkwhHaG86UdPdtkfhy0UldejRTGirsA/SlaQuFhgbq/bL3Lq7hr9Ja56w/1
rVmjeKDGUaJyOeO3hV10iOYU16KoCxR8TXB7Pd2l9bcOzUQKdbwhhq5j/u6rHxy8fMxnWQJWR5d+
HZ2Rem+3tnlPBu+CqgOEH9Nx9Pg+s4ZAJuExhh2Y6uH86sRJxxEsjc0dVWSDGanwbP9n3AA/ACTq
wtY8+9ifWGjOq8a2wYdXMpywMkmz9zbgvZiZSrrrLwClFWNgbuLZOCtv79nTWkCMllhx5MlNChZp
3lqs0Gjl5uImOupQ2xCryZeuTQMXpZOMVG7XsctXlV/kXgn4r9Ie7accu3qvmaKVm2ptoE3sb4VY
B3+0c4VNy7jak73Ieb/yzfFIP0F80frDqbn60tOtbqCAd1CPb6AWPm0Go5DxzXbsh8T1puY+Tbo0
YhHn6ecu3jQmKzD32t6uFr6MLDXBlIcwVQskagrQ3dgKYX3vbXXzje//pBgRdWCZpTDsrgSFFcsv
MKNTfW1qkLsbMv8SWa0eRIWmJdDyRe/SLGAtt9kj60EO0i22gl/GiXEtN5V3n0nokZPcNAsG7juZ
LGAO1Bu7zjCcJy9sT3RMVxeYaGsmbZrqHx5LfYeHnX+BD+XZ8o0cexr1tPAd2d44zTEz/tqLOkv7
derkR0d3lXjeNrsMN/ofgvACyobI6F+QqLbb86FjwBGQpCtSZVIEx7c7mC0JUc79487+KbcpDg6z
AAPwIFbwN2kVXbXAKoI6xy+giOSv0SJCUqEvt5thEdvAeasvDb7cEV29ir27ibqGAlCR+Ho+L0vu
4Sj7ByYt0K45kyUcew0XEfiyDdXm3ZYP20fC7tsA0yL5ZfiDafOXhKHcj21IFtdeCBOH+IrFA86d
xCzz5/j9r4Abkdrj+CvYecQDdeBwbrHCA7s3544U8uSYEYeEvJGe4dJ/1WWxhLle8vbdOnV3XiqB
OrezTtRGxSUATxBiw5I1Ws7AZrnHw+boY2m9QgMHUW7cCSMydVAWHnVK6pRJi8QAPXYRKGpHDauR
PF8Er/vprX+djXXR1BIQg30CewN4jrn0vnvR21c599f/51EsPh3tlNCqlv0uJwOmTxIOWHg+lEwk
y7M3B2sCWmv4kOlVeFISedV04rQBcMu4n0CmN2p+vXWPh5L6U/EOO3jvP766PWyKvzridayZUw1q
k2G/8iVXBTDB84VgZ27w7z3bp1U7BFV6tT54SwPAgymlIaAdGrty3XlfYDveoXHlm80xAE0z/ZUp
HzjgHm2G6aMr74DJSHprlXrzpEML7CwQTwWkfmDcYCQTiC9q1fr6OdiGI6OUaCuHVnT4YUlwEQOH
KwSYLNQ7tqaZnjfsCxg1nrdh/qDhLieVNziHiEQudV5dEJ6qXdvCc+EN0wFJrW7rLudiLZL0F0Vf
D+vNVY+kJ0v918cVJXMi3ZYbOKnK5JA2sWso7MRQwT0CfXUO0ca8sKyu9DQfOvoSIKNP0BFFbYw4
MfyqZtXzRv+/6rI8jBncxZ8SUDf2naRPmG64DthJ2hirjS5bE67ECd/a/GHN5lpmlNgPEdag4cIo
BE9VZsaETRR4uOMWS4a01TOF4aulXlCIJWCxsL3j7KIMR6CjGiyY6+t6wuFLvh9uVNQ7hfFoiBHZ
1284Tvd2aGqeRB/wrM9DpQ6nSUWhIhqofW7PsHyx/08CE/AHOTYpkhcI57x/vBpg3/J2Y23d1XZ6
NCae2FQTTBu8Men/XfFf/vr5nxPeRWjdqTZ7dp8r8fw6L9FKkJQEm1DH/YPb5muir1EKypOCiYVf
LDF3ofxqtostZe/wjtwMsOCetM9zUBG8znpPNW3rPgK/sBlfre3zjo9yPk9GGhQ2u6l0wYx3XuEk
FpScnxvK1fr5WYfDC48dC1QV5W+FqRzO5NXyY6CIOP3s3fGgpPM0xpBZt+1yGexZ2TftUB1ydmoc
3sPFbdCkpifA34+hjgT6M1DzGQTN0XakStUFi6f/+UlOq+JJgm+4JXPX8pTOm6yDVPLOYaQ2zo4x
0Vdjxaw/8B0v8PpMwny1mayDWhfnQnYf/8T0ZTstzgZU3VB1YpsYyJ/yHewjWmRL8IHBCLY0XpSv
YbymCDkLpCpIRLstcRRE13/YcvLbhy05UDT/3zvrqD+y3DGVfrOlwn31M1L+ZyCubFNDopTYr60+
8T7V59Cog06bVypx3oC3vzJmt4YEnVortnqke176KfQMuJRMYBUUdShjvQlukn5eCBiqBc53VzoJ
t0NcQeRHjUKcFEgb80W6SIxTDQtmImczyAAXO2NTwg9mc5xFhso+v5PgWv95XOTSxkRf41phWEkz
hdOCUeWWI7Kykw+7Kg7C5G4KCdEx3xV812PUqauHs24I4kS6lcP7RH8/y7SNeRE3eYKaAa6k1bFN
wOYmQ0FH/A0FPvEpV6XcJR5GhuArPru0zh6jXg8c4KcAAIh3N/ALThPmuxMA+q5ZL4FKYrLS4O+q
ZiBKyXXzEkanTLbkxJoU3OGjl+64BoT74C4LROryPNGhU1fwY3GF0eWVsVqQU4sPQanj9lW8iZym
Fyyb7yQUfM2PwZdHfNepRr1GDCGZU2ucuYRHrXumlFZfqYhEX8sUdknjRWD49zFw1MnCRzvabKat
13Po6vrLTXNoGfAP3MiaHlS68RcEp2AC3D8nAUNJoxc+m2K4oCQmU6modg0f9vmd4Ei74UKWYG4w
bs5ReWgFbsZ6dhd3NrkGVpjwqEsRC1VVXmAi/dUYSKDs37VidPmc23h01WBO45jnVZPUpYSd9Pkp
E5QqMOBci31nJ68s+cXoZ6ZGWqAmQb6yYd2b6LHBAGRaLmiohr+wWVyPTS6JrA+XTpuBkPaYPmv9
4lox0ip6SP6zXmenmCUxnXt2Ib15kbR0hyqCuu2ID39joyQiCqJdta9xglIWhmDZLsOx3jPSeybZ
1ewRLiMDwBQt4kYUws/fl3flbvrVsXVC/YiO65Vhn7sTqzFLiCd00VHpZReXWoTYGHlA7YX5fbXA
Pd+xyXOlAyzGSIXBaVxigdsRpbZx3hfN2drLC6mqtmpj9tUCI7gs+1Yy2rjSSRDtaMZHP9kPOQtx
6+S0U10nmCibU3dFabXVGhXzQIDhWnpH8u++HIB2xsWZbI9Rm4w763PdUNQDGJA6wioGzlAWpUQ/
vqj2Yqq5dti4aH3aDD4RgefS8Q3gIb0phYAJh3nc5K5T3uDcWE7F0b3ZK6/wX7nqI5p6Z9McH4vs
OI6fSC+37d3kMLxFAfRQ6UwCmHboyYDACaK714PddTFSJzSalbIDDM9rmHikGiEvlzbnb1prNqd3
Df269bUYiY3p5CW2QlsXOQYXMaGzb97Q4sGa8D+tcAgpenw6nqJcQskX+XRbZiHjVPmXA1M7wWGr
c7Z524PvcTrv8Y8CtdBDn+R6PcrztyK964KjCXO0sFfr0Rj+kj1KKqCGDOBwQ0x2MG9cAQTiwkK1
GIfHz6X6BeXTsyeuSx/suCnwskUpMo1ZOzntZCI8keMoJTLMKdA+Nkab30tBSoGSBP2d5qCMdVVm
uiYmvUBwGQBBtyu4itwI7ZSfm95UvR1rqEaFjyeNOKFkC+x9Nn09uyjuFRmiEDCZ5Ts22G+k+5Td
BgSVRoSu5EHcaYqL7yFgbzkfrwlP2kTOLt+QIfEAYcYtgs9uvbDS4WGYY+qaza7sMEdFjuN9HZFX
1MdLknPQipYldsaN0qeHeXFI3rvo0P3I11HEiEwzCfbtL18BnKEYNaB7pSZ9ju0FYhTWpcHA/Xgo
WiNtRwS/ENLdWCi+wUIR9+9RJoaRVV0Xt4DYWVYTQI+TOxfmFo+HwAX960iUI4QFlBaXJYjMGQ2B
BH2FG/V+dHt12tc+UqR1Bg6LiBwdtLqKHps+p/Nak0O8aBRMH2r4wAjgmNtoPl3L4X5+/VEgLXMI
rcbFYWVSJGzI1Z58SR3vwEdjH6/mYfRpjIPnBGd82AlxoYQwBUkmfpS1ZNQm0ViamakaO+3DKF3Q
V0B9hQmlXreFEqpTZRhG7h/4Cd8psv3AxIalvl/ukqG7seEOKXwu7DwvFIOmRzwdunTZf2MXNJKv
CdzrQn5RP7c+/YvzeS+dkfw2SqePSAStUwuSzU/tR7alEMnXn43Eh+uyyxlmb6fxf3uggS4hUSlf
rkjs1K4Z1uny4MPXXSTjSQnmv6IrksNITYavt01cRfuJQWERdv5S1xKaVro7LdmrS2QgOcJQaiQP
7MvUeBQhLgv1zJVBsD1CeU0qc6IuvxrRS5DTabVY3OGkeioJKtqz64MvVRXK1EUsYmrk3NWuPkBW
ikVRQ0nBC9D5PnH9B8GpcpJSvoUCcSH+E9r5evTuoRnzLxQDbgFt3s/liUCVzG9Z/SLR0vr+WO8e
l70Wr6Wy5s9p3QYqsxpoiBgasDnSvQSpfK/khRsxjr0wu5dBh9Fyyn3a2D3ua8kX2pKS9aQP7bAM
SxDGN+A5xNP+zUVKHEEX1Y9zwRlWVBspiYcFJZShjNbxOP1hDlMeTpPw+4eEuCVTmxIvDwQvmS/K
NOqpdTOjFAdqrvaPKfnelmiJyK1WUe2CXOMWKp+yLrlHvjY32WRFTlD1W9sJx5R1zpBM5Ss9jfNe
EdkmMeoZeIvyvJYjlC/VLL71qmWgE0S0ThFjYbL66vODaj5qGoiW2zbX2gvVWYhBUWfN1FvpKtAC
9m8/UWRvw77/pyeNRx313M89F6cKk67BpjOOjps2bylntmWAP1eb4+nUVP9yvkqAHhIqRcz0m71/
QFdYIX78cwO5Uub4vMI54Fi+4kPL7DgC83EujLMVxom3YMg9HNGUK5J7FI+lG/enPJLiT22iPXe9
UCtSXmEpNxNsMia5DQ9RiTDNvs6+8ahZ9EODmO04sM56AkLw275yh/MND4oa3/FSFGp+w4XALx7z
NGx4EAW+g/tm0D9EpYhmkkUwI7oG1U7JoUnYhEjjLDPT9AO8mdSIyK+7Km2RJ0khSbhJ6LocjYpI
Ta7Dyi1MIa40KhYhwuKzTvnEuG74ydRf1zS21HIm7ovb7LJBbpnPGejzaFxSp6IfKgmq6mre080i
CE4MSG4cJedZEhGVNqxqKg1jSxeHXmbQ8ZzxbnDhzpuQgIXMezfyqZDYaS72jNZEtr45Ohl1UKf/
XODxsA45YqGm7z8nVSbnfrHR4ty/UNnPN7jDSlhW4U28So5Zhj1q0UYLCnFGycvzYBhxwmhVfXeg
SlxeGdSd3R82EBxvoXuXImgtzzON7DScKmOiWOS1cg76s9myKkDD8mPgGYRSVQXtvbmF6SbcKFEP
CCs8mXTfSQeLsd4qM7g0F6BiueCnaSUid3ZIs9lZ0RtU/6W4AY41KZbVSaaEJgMnjfhfesJAYdLt
ifxoLWPl09Qmo5l7jWFn0wyqOEVldIIy2zZWS52cl7i75g1d5ytIjm+k+98ZDNZ0Kpu8JFQX2sAQ
HzuauUMIMN8Zb2GmlGdvsjxswPnJDq/GHgymyOuC/xywyZNVhiBqrEMlHHTwMyaZesgtzM5o48GN
6FApxq2mVkV6xPRgmoK6EdPFdJJIY+B3093+cPZ6JIkRYiH0Kt8bUEHUiXC6MAhB0pp5T00RW1Hw
JXFQZiHnGDXSn+pqDxkRrEJ5TL+HJNvvQ3HNDWxCAeDzWmcl/nsb30UvMpHSfPttds/BEeI0AnmS
kz7NrR+dkizWuy/PLWXPJDE9JToGMDsvi+Y+VcFHDkaLTe/bQmqoOntn9LYtzqtXxiqutkTldD4L
LcsJMriQSpPl3zxYLZ2VCnNY9X2ZLMh7SFzLcxQsJ0+oYyWTxNV8zmf8PG7za63ueVezuo/PMKtd
4A0wYHZ/tzqPyaEdeK00eq9Iu3tAUYuFgMLv+XIBHlCZM4SQJF59c6G7tMvj0nZ2Bdgn8DwPD0ZK
g4H3eb+eOTWAJuti9TC77kf+waZQJEGRC8QEGSx8p1vjaczqe5VULvurJaAS24s8vfyL2LUdOmUJ
ljAd/+iWZpyWW/52xLB+nw6VbFyCXr7uM050EPa47xTowtcJN57g2xWvfxJNsRXOfxqOml7s4tyY
jmKJx3Ih2C4fxIWqY0TjUWv+18ezXWZ1Xmy5nsrJBI12XDSbEE871jpXQk4OeJFPw/+KQc+rD6XZ
XMy4cbKzv91+WcilKMxrPU8NGYvL+RLT/dtFTV+OiyVJFnzY5o1nh/dvkKfazFX8PnQmRXqRPWL0
nygBloUBKLag9CbrT+T80oB8NVOd6JaKx2lbM6e+KbEfMufrb9844RYadouTWbSl10nzLSKZY6EI
zAFRSH4Qb2+PBCTjhM83kyci1rV0akulWujvwm2woowwmXRLLbwScEY22lwBJDoHxf3B4y6/5oJ7
IWpnHfghipqpPg9AAE5Bo8cOVAQJFM6v+q9OT9nWVv+ixKjuiycL45HGe+zhx7GavwuIO+E4mo/k
B5sj7VLJSIbLXDSYwSPuUd6tQGLhBPuxRKzoxnacWhEP1I48yOJwcE3gwxOdimgvQZJtOno1cEri
sXtQJ5ruFTOadfJ/5er9peLSLwZekMAcbxGua4VapKnTYCvfvIZ8JrKshpvihUPFehTqzfD9B28r
5XULLHSXb55dx78qLhmHLERhRBTiLZwCtrjtHbIRQC5vYdMP4shEMbDy11BaLN3ldoTGS7riwNWh
IyBTCNogSsnf6YV5lkYp6f99zXpt1w9xEXKwGz1W5lDpgS8hUKciObcqHi335EiSJNmrjPrH9xUV
UR6miv/P4ePoJ276HXDrH6NQRzadUXduk7gctGPcl/uZEwd1urg8BIshwF39MykU37y1hEtJgm9J
/ymbwfthCgZ9HOb/dSOwJ2OsPvJoR/9wnO4eRZSVLURmJQPhiQQW+cFwApdH8YTwex92LDKXFZYi
Fh1CpDTB3SlbFva4d+8Hmaf95FHUlwmGWMuklQXo+W01vYDhr+l2+5FUrI9rnw9E/ev0ZpiSQfAw
cVGPq2f30y1emMdwqSzUi4L4V/VFttAidITEH1bwaKdtBWMkWwKVi1NCwrGz6ny/IwYkBXS7eGEQ
ZT+tmH+slGKNwSJLTvCi3LMAyJlCY+huFrF9/TVXDxBeKpLATozJ88it5zM6kBHiUAWibwRupfg3
cVuhKh0kBKMRPyp23InCqo8ZxrElLLnqvFN8h16vz3FOG34QNIuVmKV+dQZkd9miRq+ccl8K2ml9
yhhIVu+3x0yB/v5Ulr8k+TTobHAkTwlUY9UpsDsryCKshVeFoMxd0eUxpb43z07C2bGvU5RlsPyD
l2qVS8FXUNz+MyBhwAg10Bs6YFpEegR+TU7Fsdq7WaoPJePVZz12vWlMitACJzHtg2PUVReiPMHj
Ny0V3vrpZR1KSGEIErBCTvrW+KrjTknByUX3Z4RAETnO7yENmHJ2DWYSJZBGH8Vf6yKsx1ZvzrYV
M7q6j7b3fad4qjaWWqmx2VAxlqR6M5ZzzpcSpCbffhVbQ89rcIIZMuYXl5EGoYxSHhajreEVWssh
Yz5fj2h39fBeyQW3o+q4tKBEl0QQrKw9bqXGkZn0k+O+H2nDz0cMdOfPBrcoEKzPzRM6hetlsxS9
OLXtq+lSfakC+UbUJaS6JlqROrAX5jewe72zbFKJY5JLa/cTH+8PjQzKQIXl6JXHzRMQD6zp8DYs
jCkfyW7FIOZxOkg+JR3sDXM6dIDm8+KEShJG9jhtK6Z4NDmuK47P9mvdH5vYv85DBWcI4tOHiBlD
LhfWa7tMLzMPNgvzdLcNAIfFD936MnYB8dWjvZvYtpeQXIdxkpGq8f70Sd+FHtXQtmRW/w/CRaR6
9s4ptogevbBUWkT+6281ZZzgC7cmix2YksUsoVBTqrhMQkXWdj4GlqPopq9K0s5ZGDn0GjVAbI6k
y1jp+hJsusK8fq26bLfD3RDr2t3zfu5DVt/2dPnIxMOOvzB9REfN2u8vPGp71WPD/6deIuyiR8Yv
5gDXWD0ia5XafBvA7kP0hRDfPFNXQazQ04yby5dZyWclbkbUpotD/iJrxn9Z1Z359+ZJ2B5J+eB/
mn0ZqlSLClGGnggIU8goL/4GtaEIaJAea4kKTBElaSGBNyXKRCby4bFZVf9frnWDenk2VhucrEAq
55NPq29+DoXDEn9KOaq1jL+IGW588XRHVrsFNv0yiO/GADTnXBIsvFtLNZ19kxuU/kuhCrN9X72X
yDa+LnCCxULaCYnCAcx4D0oYwS5Wl+/K7XRgP9PtTnO0C+HQGMwkfVVKhUUthJRO08tCiKILcXHW
Edeoanc5GOB28X7U3RgKX+xQJh4ygmiJwGhM4jUXZXYSBfW/VS5OBePhYQ3aE3hcQ1NKzlR9Xi1o
16TItMh4k5kRbzpPYN43Es3rrSTZX2OwQ1PhVjK5I3l3I55LA4SC8yD5MM8E+TxoacfHbO5n5Gze
k81qHtyH3KyU4Ee2v6QrplJ7vhm6RRTeUdCxBNZrOaOYinhbSYvMriSVoxybENX8kGbppnoc+FdA
BghKYt050UZYPNNGxcfUw/+SP4D/pLLFVSG9ROaKTxYSnr8TGJ8H4ev0PIRT9ooXTbIRXqyQ7fhR
lTx2D/KbUmlPu15qqKdnliv+aIC34SA2MsJIcVNZY2dhyD/IbCEqVs16yCYppJLcLnKF8TblSj5g
SfGttX/ME9uJNi199Xc0IPROkOAY4xOeyBOlW0R4h+3k2yAdG1nHCaUsjD06NRbpBAK7mGo6btlC
Xpx2LpRq5qpN0DztaxLYyJlQT7VtdheVyHA22B1DtbsHmikOp21cbTWsVhl06wWm/Ga0jdczeoMt
oDgjqqLeO1l7UYLAtCH0WgLh6LZpdiLMCZfP/E6PG8qszW/G409c/1MwjiUDvNtw5yNAM/IztFks
5CbHhhE0VwAO5nM7qi++yV8J3f4+YsdKIT7tK36JvdFAvQHXkrmDngtxqvmG5a/KLI0Mb4wViL9m
GCRL4k9PuRR1iXE455EzaD4axHsfeq1MPLKbMhxMNf59zEEtY1HoYAtztiwkOLntEzIaY5FBrnFl
gvJ9ojbe9PIKGS7fITi5LMkU9FNHN2T5lKdMQ2oArQV3aebyF05A2Mlun7/TFv39n67yfwEklSWs
oovNvkT2tmQyTlf7b+pl9pTDjj1SvqD/50GKWtX8qZx5nxwx2exbks98ZtpZAD8kmuIYv8FixF/6
v3EwVZMBUlED86ZP3fs3sbXm5yBBl7VUxMf9neshxIrktA8DL7zW1q+7iCEpE2ASjQmReU1pQXGw
LrfMb1QDs3YKJ1TieTVzsVwt6P1f1QHlSy41TiAHObsRf0ARSZpMSqAbclEMGjr4fdkOli6Yzgpd
FskkB2Lk9UpKVmkyeEy/hiKOxIBPQCWC59siMlEaHHCv2W+LBPCL+BaByVF51cF8zbemtuN8KA5C
gJlhPVqvYCVDj48DO412Jw8FNJeaK8KwW+7rKvjGjQGVFRueHAwbVPH4yYwaruVKRwDUvP697/05
k/TwQq24WV6bd8s816WUoUhEqXRv4ArPlZyUM0jEUiiR363Rr86uJmuIFtib70TwaGdvLSoL80pF
AEuM+Ut9aqyhFIyicBMVdv6AcEO12FTdKXhA6Q05MwcjthEpIZYxxzjof4cN0KGbMZ8SPh4r8ozW
P3dHtXvh4Q0+A9MxEQX4wuMdk00ddT3jgGRLxBsgxU13rf7uOEJeBRlVd57xJfO/ri24dgwSplPV
tV0fRA87LG9lRN1bWaqi0I9tWQulUbGfM1SUjExx7886krFdMIR4hCib4bB5tPfh25YolxnTSmS4
R+5RdKb9+HKD7WGFyH5GWROQ3Dy8MkAKhvTuxGHTDv3AdISS14SILUy8zhPCfJgfmFI647hyv2NY
OddqKOjQJSV9c6tVD6Jw+AUM6T/HGj6O4M3kpC4+w76L8mQRnAI9VU3VfvwtAswQxPO1nSgwlft9
1N7DfAzQY7yY6NtVWf7T8copp/+ImHmtkfeiWkY6EtauPcjrbqcxftNZiSi75MbudMKim/qFx7K+
pmqxNQ67F3/8WUaFaHKwOLXlfNvENqCosgA7T5oyYvNB/rFxUKw1vWxuS3mJzqxnTEYpDXUkJIoU
FtNlwYZ8NOxnTTLGz3nGX42CNg72uvKjxDdxqWnN7dp4ffd9MsDGz+2PVEdcEoXShIIeQtxBobyd
FVxIeAfVoEQ7tnp3mt+ZL7bFOn+BCkicN1u/I4vwBNsb1KFJorb6bG2zUWNDo1zzCZlq9+i1L7va
sScQc7Fj+JFtfdF87CWH7FKfp5pzxubCIAj2o32X4vko08DJ5t22XEDczgXsU05vpFE/LhAIT2ZM
a+Q5uUXq4QY4Uo9FzQu+uvdT55NyKw0Ja4CtyrKZUQDoKO7WyTFoYalnxRN59YMczbU3GucZg9J/
L5A9U4fQOy+cT8k0Na4BT47OQc7oYA2m98Cafxd+ybYsUEjDkJEbWvJd1PBNA6SdfhmpSkG6jZjJ
3jHE1Op2yaCYtBW1ozxToSILA8+hgof5ovF3Z9btBnhtoeobB+yaWZH8/w9VjPGFnN66IOlWQfvq
Sju3JzX08C9CcIcx+NCb1OBiCFAGRk67gR5VrYnQaee2lfPQ0vyjqE96TPZ5QVM8W3HI02gy4AWM
zD0rwoblVX0fY9aIRidWK+f14GvymfeVCQrnJe8tmbf00eQDqnlrquwTF6bu2kYaM3ASw+okHZwO
OliWpuq9JleME90WD8njottD1eHEtvMt+ImzLUaiOf6K7hxyCkr4y7iC8ttJN4UW8wqynZhRIXaX
BeeEXzFyOe4CncKIog2PAN8Igf5mUJkmiH8lRbw8usyVNOS4ojgK/qCKPxpG6XnoO2xgYrq/og8G
h4NGodSVjHdns9yLylA+J/0IOSQo+fx7nOfGEf7kiDIRhM0Bc1c67e/CjFTi+wW7AnEdTBM19ENH
W81HeqUkPBZAaDEed65a8K2Iu3cdsRon5WyNCC63NLMwxVi4RaLvI3um5iomjnQYjEoM8RIicCRL
wHHMT8eP1GiO7LkCV//VaHLcH1uh53m7+I/zhMA5PaYNAsBfAXI5dKawtvF5EQFeus33kdPtc3/t
wlvNmg0TLn0mCj6UkvZ+R7WCeJdHz2IILx0fJylcrNz7Vs40i7TaD4GCOdWQUnuuVz+igzTm1ZE/
DinS39n2KGMRCxEvQ7uzex6nG70B8DpqPfmdlagKszeZlZXQeW0VwYiQj6Z2YygFVGXnp7+n0w+7
e8MSYnzFmPgK6pF2E5YRVZkd1ea8JX5gyIXVIrFAM8I5jcVQqEzXkeOlrds3YVW3I1i3B6yYf7FV
lpeu1UO6Q+Zxanhm0N3oIfxSJVgnWG8eaQuYFt/EOrAE3yL3OuX96uhfXNYltl4PaI0xgSu812OF
ZfFChCn4giQTz3JHipvQdAl14IHNx7heIC20WJwF3ExuQ6YnksewUWe9ykAyIxmKKAYUSF+BfxxW
ckbB1tngQfm5zDd7+d/5JKKQnxtDRBKOaVn5Raz3MqODZ130aAS5afRCAM513tQe+/5PfgJjNaeZ
euZ5U7B2D9Pt2kZvojJHYBuv25fLS1Pqn7GsY5PqwqRMUR9gysbvqPyDJtZqLIIUGaWMHIh50KXs
9bsgbnhY0xGHs+EctQxdjo5i7KrnQtGQCYnlOf2kzm+h2wiYWy7emTK5ng8ybSOfJRsAKnI14Xwl
GgDfl6mM3LBJwOwd7u0C1+iggl9oipo6Uklamf/30DpIp+T4IEAtSqCJJZmS1orpKAT3jwl6eQsS
PtlTLY1NQo4w7kVbH6Z/CGxqGugTBRLp6yX+76GrG7kLLY674d0pxE+TCXLJ7Ik7SfgD0mK9/g3l
RME2ZHAsh35XFxHjXbE71TJcbfE/pTDKBJP+UMJew90fOywrTyRnSFY+zDNDVJKhg9SQ53bwzYct
iokWVSC87DlHuctLLF6z42Ow2N4WOWEV8I7EfMghhLg/XjQxpyWVQKjSGvKrOqyOvpB4R6fw4Dbu
hgkZVLK3vB0NWFoiAXgmu2ns2x+EO7nlHOi3+q+1fsG6yIkT/peY9IZG//6pVYgyepVgWKKiJtpR
V9FlCP6KvFo1Q04+I0al2TsAssME9+o6Z/fyi6PcHhrUcKvP06u6egP1DsxVKmVuw+ptcx0+n5V3
iKVgVTodHsvVBrE3cJh/TUC0k4R63Es1ucrzQBK3rJT+9+Gf6sXo+9Z5MTDIbAxwpv+WdpL7SUhk
B5I2x4CiC9N7/J4tOCupDFaDiTOrqxOrwC6Ut+wTZ7vLr+eYSwc0A1XbfG9Tpn873oknbazlF8gs
0sIhOyNv7MCajhCVgVQ4hacj3BqhQHCN758UML7aSlF7iOjW6YksdxHtYwE/qPKWARWg/tSVRNvU
idMBhN+frS1Wgm3V2U5cx/nZIdPpGiRrXEWDqTnK5p8IKDvRcMpwMO5PI2S82GvSurD+o4R1ve5R
nUhA+L620ZeqSpl8ZOOsP00ZY+TFqSitR6lwJuS9QKX85DWi+ZfYo0V3SIvb/CYLqv3x3r9qbEPi
itojA4bfOLRude0s+lOcGrDeL/sOUQ5uTbQdQMUUQ5xdUwBvNnuj50E7UUagzWqsm2HVQQzYpLE5
4AoAfKkra4WDcvKIHUG1gNMr7ZM36ioVmB54GiZ1eHIFtBw+PdGEluXRfEe8CilsuFKn14lhZsZM
tK772V8sOK62mS+35MPCN+rJ8Ocmf9IQrbcGB6n10SNNHFSXfcc5wNxgx0dCuzYiz76+aF9mQm1j
yrDPJe27R5YOmbx/Ijosr4RDa6jTN2lG2SiELfJnbujg6SBdO8W+5a4yXsh67nxXaVIXhlekndkJ
LUyRggBcu+RBCDp2OytjBxcNA8L2fRfGUnu2EFUvBp3mcNyOo2sdSZEZCQrvvd3Rv+nfI4wzcdU1
bES8ycGiox0ItTkFJKi87dSJe1SgyA/1Wf8vsjQa8flikRLB4TVkw4S5RoTTwV0v7vZWNXchi0C/
dFCV43mw2LONxVWRaExWWXcnd514yeBK49UfxOGgFm+PgEZzvZidWbAaMijnewaF96/QT8/eCxhB
87idmwwNsNMYms0rsr3gmjFaVbRx35Ai/5Fph6U9zlkUTxgfSlPGqEGBhHiwQzrqMVlay6F5XtbW
XRLVAJcAh3qQkz8d08eLhQaIni6M1I3w390cvMw8xc8TPJxB1E44pC9BLrXpphv0rmWC+XxePTiB
NswSfaOzOVnDgmMbRmEdfogbA4nbRwRjxxcLa1aLETSVbMdgvycUmptEvvhpaFzm2ID+tqAOFzh6
xJ8Ci6xYwr05iefq9nlWNg0uMNWgulz6e5NCA6LC1t62a7YPPIggw5DcYg9vPQPw4tOwyOHSv+M4
SLQ4nn1pqyr3z1gYipUiEHPkhGwqmvFBHpLu13MJ8x9jaNWTbgPbEzLDk/elWgX+WWEEUL5gw9TN
R/dGmBI431VmmGOF9p0q0bZYF88KCyeO6bk61CSGZuyBZaW6ZDNgd10yXQ+ywoCKuIXBLefjLHaC
VWceH9aSjwOXKDAgdektywJ/UrhviTkEURZmpnEWK92JUyqhzc2vnTEk7YvHTUmogPGsHWHHqr2s
MY5gWgWvqm3W8deitmHezIeaf0Eyfkd5/r3PCpTS5WFRkbpIoWhjTcDp3niEfVV7Z4/gy6nJfA4R
uq+aMeTK8X1b8Jsqf+e2eXgYIdRCGiZL6i3A/J18tzhZUqCezjni9Ix/rthobfw1PE3FA3+JjLte
g3Fd6MvnbKAlO9qqpjWB1jZu7zH1p3epoWxtVVSHC8V4GxF20K+bDmKgD+9xcLMzNceXrUrixp13
moLfiUTkI/Kk0YkRzf0TTvtDgtJNLBPBarVm37mivMnCAb9TgN52hG8I06o7JVi5IEA7YTkhMBsp
DQ/lZ9UCRYxtJkLCV2ISKYLEu4ryuzBi9qDyJGLR1wQv0tPP174xTWiKu2DNtRDpUWhw7cUeYijW
REWtsC6ZWVGxSVUVIpFIsuPa9hHdpkjvtILxavrLhYaVZXmuASd23wQMwIQjn7dz11fKU9q/vWsW
7KfwOauZ+NJZlfecthoVL70pv+y8DtVvutO/8WxKSNbIC6godnWZQVzZFg5cAaL2emiYTqfCqQm1
5+oeGGhz6XNVjttUhhxWG82VSrH95JTLJwOr5Q6L8Zp8V1bsgcZeQ2YUHDM3fQbvs9edCibZmh2X
FWkHr/fk6Nj0wbe4qxjytJ7ttTLw5qPocngiBFNtf6LSkQD7XapgeOFmzZ6giz/cxZGjrjwBWZ3h
w9Wv/4Dj7IDH4ZT31KT2Y6jGNJTP6N1uMk4FOp+1MHpzW/Yf5F4nqCiP6FL0QZIfBt3+JejDtgFA
CCZchTy1lc/EVKozG87QI7Q8mhfq3BRg2fWcu/QT0L0roBU56AAJnqXu9eOzYik9dJFx0Q/rR96C
4J9bAtBFAjx5EV1m9CcN8Bwp1hbYx3PXncI08EUBK+mPHR329Rw1akqgM+Go+Ga4w0qnwPOoRmPA
ScH8aAb+u59kAEBRtRQm59Dk+oewPpNf59CFwzl+f5aPz9jmHKChScOf3Ogfab8W/i2K2zqYpALe
Hx/LGMYQ7i3zGi1AYhnRkmyaWKx7GJQ99i3mxvSEJ+YbRXfL2KFP6Xo69isalCSbs4zZcIqcv/21
S8rz7fGAYYsYXjBkSB8Ossu4WZ4FkbrgWKde+QzDobwdi/9+p9GI+1wn6n7lhMVDa+rR6NEZgum8
4xBUp2PDK8r4zqCNzhSbIKpargu8LbVdxxGpJWRb4isZiKr+Y59+HeMiW81u4VEI1/3ZYXoEu8fd
Qxh4CiRxf2ZeuBInNUPcr++tdEdNJs1f5NKOSJFf/HlMqEgzN69TK9BRfz0PPHCxSQWMlW8q0AOi
OCx9aukUC1bZWuxpuV6tQH1bMKL8L+BL/rn4t0vuo8ZTLbJivFTDK6eEs5nAhYL38+2mj4KYR/8A
qmAkgrD99PJUzzekO+U5kElrB+JGiBI+xE3lLbB7N6fsG/YhWAjeg9btywnYPiS3rK/6bILbPe4O
APKsq5p29nQ7Z+L/hNZP2SnnkbFK5HmYHn5eb7zuu61SV0ITvwgSoEFoBKM5UBgwoPqHv6IbPbRg
ykLiW1xRAnokoCGHQvcHswtIYnBP5Fz4Q7K0gm81LsIxmb8gHksckJDF3NvgJKFG+bvzC8MrEgY5
fz/p9GQ9K1p5koYnMUaMWT0++7m7MSKmnfdSjw9P7+VF5yquGHD7cfx5BNHFzGWquoPUV53a0Q1Y
aoIQAyT/DjeoLHzp/gv8rUNbld0okc07EOuSLnFN/Ob7fvfypWZpgRFB6BGeQYeVlul1VEv9SjT5
V1cj+2ozAJbmPjjLtkZpk7eK8HhzLZ4bbCBsIUafIHzU/yP6mPQljRNb3GKVXcQ9+GqGQ6Ok89m+
3CnZ1QbD4V6KXF199T+zwdXIoSFL+zClPK4mNP2He26GQxiT+28v9xyIeOBuYlojPZRdOGUdTcm7
DXahXbhXZT0vJh3Ro/6MX72NV25geU3+7hMh5ZfzWmsb7p7I/USKN8Pn5zRwVo2jVD4iVaDUDorT
EUDboex29gtL5JtQYvepvnI9S2IDfNkSOLvMyK+jnuTWX6w1cnXcWYc0dIi5dnQ0/vuAisiuG9oj
FMVZX+4N7WflqekmdSCq8KEk2VmhTHSBoWSVI4G/Ja6sVwLmNiXiPNluCIUk2ASvp0RJHCrKzMTU
sPUItslheOdVfM1LJIEJ8kA3IxG+av/u3Ful/QcNOlqKu0yJqMdwBRmW4iqRPTE5Z5JFINqPdgsR
dnBrRzMrW7hq4Am9GjIzK5LkM6AsY1AnL1BkBqPOzUamLefGH6CV5D5jYsdUs9txZvPajukqqvuG
iehm6IeS8xS/A4+s1R8WXaxyu3qMXFP5yVOubp7Am8kLNEpmSFFSGvwqThdCrRcOLSIj+dVu9dIL
CNxCxMz/q32oYpvtfiApU8KTFtB5gjCHf+XRHW1qjS3ycZnoYx0fRegWhDf2mCYSdifyE/DEacp3
9WsGeA1dZ9UQifsdLItNBtUuAOzzauLpxhFZ+kfBgBcGDzAnlbHSqnbi5qvsxSSqukxh3hOIZ35l
N0nUlKT7ldJfHxbFEafy5O4yvg5B+V/RHR6qvLJXjtQFmdjzT3nOE3geuCIaFikDm88ZUskfFsxh
wQ8fjr+ZYpf8Ar5ZNoYKJSbM/h23oneJHx/zN/9Wy3xomtpLLST0XElp5E1oV3t4qKSzBCr3GKD+
bRExd9fIPie7HJYJl3iDbBF7aDKJhXd668vavLXfecXOpU5LxYARW/t7pZFpZVMVFfMs29t+r18H
aNZCAD40oawwfaxFEfoWjMhe/r13VvjmqQ9Ap9cg4TECLlPCkLFKWOKDOgr9RmxIlOIZsVXlBMUn
01/CN3/+Nlycoch3zhUgPd9yroKi/ENR/1YUfWfNwNXKzmwqBJZXRrPJxohcingtYSIAq52OjZJD
eUaRcr8qLxvuL+JlHolWjpOGHWmhsL06gnDfFtsgkUrG5BhqVi/Iz4C1fIAb+4YEdd4CInhbMHTL
JFMsiJeN1Wto8fwU8pbHRhzUgEcdEALU4NgLQ9XmAqUNrqdoNJKUDqldj4a//OpLSco5wJ87/vUW
f1gTgb0skxbrlZ4DwecKTa570eb5hleRzil9YrrwpzHNTzliwdmOo0ft9LS8UcK0i/ahadbUrMAu
8mGSfZ6tOMyX5dUC4xXEvyObyrAkhynSUoE9X0NAQU0vGHobnC3bsXjh12OXXcsE7FRXLyeVqvdj
+FTmcYwTvSLjIdrSQY8xwnoZNnPrw7t1Rui0DIKco8usFd+gvs5Ewo7hPtv9bGuKviZqT365yOCA
zOaVHDoAp/X7PeBLMAFJCrhrjAXt6RPUdzaNxYXVIFx4Ax+rjAklcVm7K7triT0tiEJax8qPx6eZ
OlY0fub7NuPRiE83nwhPqTQtb4S4xrvAKBzZmQ+Cx2pH4Nfwpr0VzjAyK00RVeygV5y10zV6CoyM
wGS9jmkaPuNvcDq24+ALEf9xKApZOSbA7zbUL9/q0nBYDWuEtI1/7PQRXnqj2rOPMvZZ7UHndFRK
Y0Tf/BUuQSqRV3EFbgW4kvQazNoZ+QfNTLpHRXWf23+ekOckglI70lhrGMSjlOINiZoFdY6cZJex
oolo+CpdJE860FnUzDP0a0SjRaEaHPjG1OLIANwQjkFkmWQACQbN2euQAz7hnJoywqIo+PZZRvyx
HT2j7hW8UggSXlunTX9q4QyDQpcQfJ7XhrwHugGHvoOZdvYojGGy7oil6n+0k+HalPKbIjzvcPY1
YZoJ+y27Yc12YEh/B5ZS8vbX/MNitzUzbJgHBiKKh4e7aGkH7s1aK5ulBBxQ4levYHbGeZO3qrb9
1VYkgBVWb4laaP4dWrHwJczuo8qlu6mhojGjVSzWKInrf0j+0Kl8hlGULJZrftKU1nF4KhqII9VV
gZttzmadMtZc9LhWrB1inJD+KPjqzrq/kKWYh4HMdcsW+HRkwMMQykDydHoGNvPurRXImceLwihM
1kG8Ig/qT53QCpccgazvO8gs6S+qjUWXsCzYgVdds6vncV+u7cqpGoImfEb1La/sPSossJ6HkmY7
7+54l5HgBWdM47FG2Tp26jDs9aWSdo+DIO4NIc/y9TuhYr2SAThuDfWtZLkS2yDF+HLXAGt4moHF
xeSFJGV4jBeem12t2nPyGLDKfYc8rLu1bZXYvLY8h1T+tQf3CK0YgI0oxxHHqwk+D0zulzcFJwH7
yDLZwUfB0Ft/QpEbN4y2h6giQmCGr/5e0UZ+RYZj1o6ArPGjvnQEJ+FwNNOMjxRyQ8pxV8U9xaxd
xxJxlYEsTRPChj3nnpxs9hfm4S3kESzXoSrLWnoUXoHwdStMIhY4gZIeJB92zkbo0/xnn39OcTLa
Mg9COT52JqKAdfC52+zuDH+xKeRr40O3Y33ls74VA3DOvbuTVsO2QvKPhwT/Ls7qWiuHZeGG8XwF
vUein4SGewggpXBuRLobuMHpWUd3kmQ/7qLtVaknRvo/3m1uv+3mYrMdPVsHJfd9flINGZLEFKiE
WjiZ7zSSES/JvSCjBboIB8Tf6BI8QkbADDGRb+f56RcT0cdqyp4ncHr2wkrZM+2SZKHzSFFvAg4o
+h3v9nBFOKz8NXGzQ4Cugj5vbeiYHBzJxp2SFvxjgcIds4bkwQync68EGcFXg8aD9bURK3PEXRGZ
yGMV6owbgnB97NVhqoaCSsv17J6iPxbNxj+5B8NsiIY8fY1Lhy2E2TIrnonFCKqw7nPESSxqZ4p1
PqgU2UpuuCtS2Y0Tc5ttfRow3KPqqLVIt53QMZJH96efuITN8kkKtNiXNl+aeBm+tct5O86BS5Mg
1JEzN6wv8djU+x3HZnnrlZT+9l/IW78BAq2MLhCWLmxkUVQczaE7sa2BgHkSvUFifQJOTEJ7pOXc
57VaZ7A8HvBbIGgWp7bKoL9Gt4JfTL4P59jzxAGQOD+GOlrkf3QFinrKB5ArtCA9Lctdzei5Y8l6
X0K6bOlRvg1sAbvkclEm5rfLTLepPRRnP5i1jsSsA+Lrs5S+t/TjIzOEHHBbOqSrim4FAm/97Xtn
JBYONdGS3KtO026320erZL5dgwm3sTGoiV3Ab9lP1fTQHkISOocOlI301uhr9fRd/t/Js9NrOCv4
IsGWhg0WD6xlgqjTYnfnZeAJmW1xjOTF8SIVLppjpOfQTnwhAJVfqDJ5nl0KD9tq7Y/vwo68pFCu
d/CoAunR61+55wVi/Cx7nJlN0qbAhS7ekLEUO6Ylp9G1BitrzE7F8dzGBRl5qHq/CAljGokFkDJ5
x+XJl05kV10fIo7XKKQB7FMvYzHvgjt/E8JDrxIxstL32oRVSE4lMKJk7HPRy6WkNFfRJf950OIE
jp0zNxExuk5P6G1GWJ6n/PwZlA/7VXhQ3/we1kzs+BRVL7de5Er+znmHgOysyDs3Okfu8dyR3pZb
vQ2K+J+3DAIIIfXFAw4CyT3Y5qxZpf9hq4+EuqfA7nmTu2gXctyyYHsNW9RFXGfIW3JwVVovOpDx
sJrm7FPg015U+4N6TdytcbmLN1hwo5DPrMzuiTJY5dc5Ywzqyb3R/loNYPKqyMroC+aB13mgEELj
4hdHQWIPiUTltNc+tt9vEshn4Uk/5TCe8mxtM/xN24P5HAtfMJsF607odjSp4orCbCFQfYonMgl/
Ou29ThPMmktKICnXvwUuKHqVhsP0YQXwiUhS0lqm0LU5AJQWWAWP+QlebfdEi/F3UMuz2RAM/5D5
captEhMV2LZtly1WJCdc1Q5S5RurFvLqD2fmWmAcKPSNkeh98CIfTX9dhPXDf68QZSaKmGx62qsw
3Go9tLL8ZmFBybChN0TCu0omCz0CsTssrEiarpCFf2d1nJfcWYVfCSuTLWq36E/lpHTN6BIh8sbV
Mg8ihigeR75q2xR4Tb7uwcuM54ZqSrdIJJ7Upbr76YpRtVB9VdXx3pdB5HQ1+QXTgJtuem6iYmBG
YVCbH9PqJpRTw4CEeyZkfBbtjrrSPSBvrlwZPVl19TaQtsswyRdsN4Hf+S0JRmP5BcQp36lGSKGv
YIpBYkhcDt3ZRURnxLr8JHlHSqvu3lMK1mWblivJxXap9Afvs5Bskvi4Bq1lUnSGjzZh1J3SXJd/
KaJkIPm260GrKNN8VX8aTCu4i7SwJFrQ+o/Ml3Xmmo0Rb1IcBjotlGsypNHq3k8DX+wuY4Qf5DpA
ZAYJuL7Gl0OfMNneX0QcYhFaQiiHWckloETNnEWLWU0oQGfmVKwpU2gsyYiWT3eYZKoh/kj+IhAJ
MmKJrWkDGvYuyb5X2yZKgzb2D3/62C18Pik4OjBspjGeBBWaNqmmXa9RST9AkpB9isbC4ZMx2YXT
fg20Oh9Fah4d5Sw0PwftG31arwuZvYUs8gNL8wfAdaOE35LNRRwaHpKK/aMfuJos4sQLQHOzv9tJ
moa3B/ZPhK7D6HqHW/jR6IV/Kd/Tz45JRwWksiJ3GQEVanDIDI54WdyHrcxeLWwNY010Z5NhP2PP
9IWeJ7+V6qF+X04iK09quw8e0pBljaDnxOZ+8hb0k7r9jayv89m0QJVxzw4kmxYET3VJjp4mSfqY
0LKw0TsPtxXKt2ZpoImKdLn4voI+ilQrZZmb/joP62kWVhAMVx/L2aRSJ4T35xsp21UaxNa2NH7i
0NAqxvRN+fGP11wF8aIduigHvrRJQuiQazuP91KRzu3mNlKTmANIQAFTnFtwzRwuABhXzZq8OFFl
nuHEU5ug2efseBaVjRXBHaclV4YkZGj3qzqVBB16U7XrlDLEolCj2WYFEohcSCUFm0OaZ8S1UxA0
w9TyF+wsRsehwc5rdLy7i3OgA4vls0EGKMCnMV85Bkuv0CYLAH8SuRf9J2JaNYrhgyxcJ5vK3Ru4
lyy9SZ9DlHOWiet45hUT8sNQA7u9Gh1szr1Alv7P97Pxh/WFXUypsinUVxtMYBpNWTuPRWjOEBQe
c9aBy8DhEzt8QKVDJTl95dj7tW67nCHD8b2RV0RxVjV5J6yp9IU+yUsbHyhnHRpRSbPuQ+SOhHLC
z642WETj5i4pX1ndiiARVgs4fCOEufV3XDurr6aRih1r34jQM5c6iILJVHvxKbBKtxtHnwbaqhzD
ulb+WMhnAr9sThjfeyjPoBaaguFsaGz/Gi0Vvyk7cnJonmG6dPX9mjz8+dOObQGhhmxSW/pUMy3k
NHwxjW1ndtQThv8XCNM4yQzYviUPCEu4Aus6q9iwlu0WYxUotrR2/ClMdTRWGFkRA5dezEttG/kJ
+wuO8qlphuRhDnADhmGRW/6+6QxUIixAgzL0fzuZp0N6ljxFScrOtwKViMD4diy9RY8FYhSdG0Jy
H0z6wvY3c2o7MJwvhvD5yd44OL5VlxsrcnkCfI0WZO4KL7EiEmfKDFMCZINPQTZ02/N2dG+DBFgF
v/bEsGwbmqyzj9P2lwqT7jMVxg3Jhhb4jGzWZeYoxoqcHlXSBMNlGJYoOOKEj2hEv39039EM2poj
y+icDMxn1UFwZRq7Jf6qG9X7trswW5uGuu0QCk6emhSZjhkWvRThJO93qJka3kWOljU8AoHFmq/Q
VObut2fuEkaNucPWlOyv8JK7xARP1TIqtGcQBALuKScIgJdL7tTJ22zbezG5AW8LinGBo+Edc+Tr
khid3Pc6tsCrx1MSWHf/N4JcXBQphi9G7yyyvnxgFjA1KXVw0CfnfQ/DPC3B6QI4GKKUWBIJ4mxc
DpT8ls8tSA7UE4c35/x3jxLwvPkU05O0d7n+oPQ9gUPzYpJvdx78DyAl4PmdGdmBzghCW/JLjZ7A
Q1KAN/Rh3y00gvYpiWrKSJqNpM1LxVZJjkPEihcn+OW97HNGGFevzRyzrub7kysVruyiRbVl8cE+
wI+qcHVgHoBp06bfPWeyR1aFbeL0OzAm7DV1a1HPyxg4usY7f+JfaqXW17sPmn+lRXPE7P+QSUiZ
pgJSQ6NNYrZ5hz74miC2qSmimTgbqY/7/FAADNdpmlf3AGPgaVdAK/Yj2Gs66ns/IhYf+exz/qeM
F1WVqfHXEeaIEwKdbrnqsSW+80SvS8tBQrBNSv5iduc3q8DUjnWRbxZjdjuhoHNvzSh9jQx08P/v
xpr7DZizpWNxt3ul6wqxTOVui2GUkzN6fzjMbTZ9y4txz0hAHdedpNPRyebKWvKl7mpESXNgvdn+
gxMhYUX5iSjT9cPic5bTTBM/Y4zGtCador85W2Y2KfUIyPY/Y7eO7+Xoe7m6i5GYNPSyGq6KyU0f
9aVryo5fWWatGPGp17rHrmniL820Lo8rX1FR7/1IveqieI3lj27AzjjCOaQG6B5r/2BsIRxWoa8D
bHkAx21pMTTZvL/jjLxz+6wTPZXs2PQhj8rMgzcPwTinhflN6B8koFGX8gLrrAFM6/W16WFO4YQP
+WcVow0gTesxFU8Vm9fZJtxYVpqMmy9in4j3XdafZpNRZ2YNkijXRPqKZ3jXlioEpCIQCOFIii07
5ths/0EZeNY6gxeQpRPjg2KBWcmAqIfa78kYiW2GWJWT0upyaX0qTf9brbIOQ9FKH+8pVb6Ajdg1
slRJonzXlkBMDCsq6Sv4zCro+YdMq5dATdQ3TeL8NrJEp00K6id0H3hUz1phlad4uSSQEObqZ5hE
o72MC3dyDRPRpLGHonwsdPrVLW9HRGrgv/SdnwgKYSMeJIHH8m9OKBUq0+Cvd1ez8BlqVQQxzj6s
UL2BbzkwLEqU4ic1zVvMmcsIU8FD3dn4tSCgXVoSd1wWdCq5G8v/CyCGDIEy7rUDUEYOq8AxUkjs
95yKlPd+KCRbyAVXbU4mmpXkZa60m07dk40ak4NwVXD8DrIFi/fi0q6+BmFF01KSZVCKzv4rNBCC
NumDZSVw4gXIgNwk6j7RHNW572ZtwtNbTtg1uqnA3itzUhTudDvfzaV3u67rfeL4aDYr5KeQKahx
7o5kieUNcYOlRV5QDNWKofaahMAj7kULiwng5oHKF85y3hOaoOG6+37pulDL+aixdzS1APBMsqLg
P7YkAJNV3qtrOG80fVxgxKy8nso/hH1wtSCedqD6bAPXtW2wf0QxMOQVaQdd8zKyys7ZMjNP+iOD
ZoeeUnTlzIPlEko+DzFHkqEv24iw+iU5yujijBtBOKWS2877NtRV8hHamSpwqHJjGzgZ4Ol7NoSu
Zfn7g1Sd7hgD3yC4w/Eb7JtvIolDTaCnk14LIX3P0VSMagJEKXsHCfYFPb/L/T6QvuZrIoLZTmL8
oEzLhbUWAxO5PPIgOplHggLXX7YLxozQppWOsfoFb3jGGvzmQOwxnBK9xLemKVq9vG5CBllv+urm
GEjqIjIRn+Thhu8vHFQaP9PuEpQJ+2Wyt4miMcsAsvRvzIF+kS9bHHF6o5qiyAXJG1jEE+TZlA4J
bxkh3Hn0mG9HZnHH8Sd5Ivnt4PZbtwcD2jM0QNrZROAfnsafAN8AXtc/wrecbWDPTNoz6KIdggw5
x2kxcBS4cIjgjxomaqu/Vy5+xHvhM2p2QZhLBukNsp2E/DhuOFgK6Vo/vCyv8MAwaiLsIQTcfpdg
aUUAmOUn/39HqUg8CXcxJS1lxHo5/UNihNKrK70AllKFsis2SnKUeVdLHNBiefTwT7m1kDNaXdZp
3/XDygjyzMENATRo5aoKSwRKnUlQh2X5F0hanTJ/g6LdnrlIzSJzDobOA5AaSX5YnpWrg6yYev5U
D7QCRRhG2bRVFTmKSGq5sj2vEG02OyRzXuhx6QL6NVc6QVaEHKlDM9i9AM2aJ38HXo7eGopTgbmS
jWvCQwTsGfcFs7zKowHvXXqh7Q2yPpae+GhFQA5V4dXouP4kXNDP6Sob32als9d8b7RUJ4GVXmB7
ne/rBcmVBq6i5F4uulKTx8/s9EdogRc3MRSRU73paUo6c3ErAuv9MUPIndz68KXDkzM/GWhEvouM
i/CjmH26INw7as1QLJA4yHYnFry2UxT1xEHzQeLGCR76MYkdvjQbsdIxLD2pvDEQRJdj/xjvp0jo
xo+OdsDIepmOc3N/JXUC+QnsdqGSvcl9gwdA8eYJW+YXEaQsIvaRN/tA6MgV4jIX8MyIZY66thQd
y7d1Ivd/TAyfZW+M3GzsAci7kGH96f3mMMgMF1NfKrOQiK5W+E4H8N//D3ilQ85Czp8fBRi/mCW4
g/upOo9EoGJle2GKzajqpbH7Fk0ap7OJtyss1m68/P/S3UmHjnG9utfDbN+lJcP44tuqiCrjx14f
KpLjQIXeu3a6kyaVIt24vBazmtPP7G0Wy/9NKJwnW1jXnlUKksJPgFt20WN+G8mzR3Zd8xyaJENf
8p9EYblXjoCZ3HBnqPrX9rBcTWxxNy1Xjb5RKbCPLSbSRHPtMnPAzdWwavD8ZBlcLN5fp87OEngD
NU+FEHFt377tJG72+qz5zz7YSbGaZr3v/c8xuTavyC0ihQAyl6zDnHJlOmev/m8IK6yNjR+lxQ6n
FUGlSXugBLJJ3NhODkHXVOU+HtO6yH8WJiHdqTzL2LWXDbrgiMbPqh0n0Loq8Fj6zmU5l2b+3WXz
m9kAjTKD7fbwv32ApmPOnTUXJHewIlp1JZqaKUESIG0L5Tv2rpkRCtjJ6kOvS75Z1fcNAFFEtqr8
jVlWsnrp9bzY1gIiBVuGgys5SD0beQ9bSNBr1cvaW19fIBsqkf0Aod1SZTB4sDQ77Y0tuu/puc/O
1ZIx5CJPnSS6GUiv+xCYAFcU3SK8NfwVK+g9oZhGplVmggJFas/VIxHQO4hAvty2Xaim7/rlQPWH
gn1Revv6ygiWPzvu65aY0H9vua99WtT9ePxbdYwWmgm20X4YEEpOOMFIrgdaPBP0lgWwf4WCXlHC
H/L/W6QYNeAQSdixaQ37Qu322BW8YZcowIcyLSVToZiTTLhGSwl9MUkB61xCupc/mAXF8RtAwaIQ
paLeqFWlpZezFjiQ/GZHEoXLesPwR1tW7tclDMSkJt0S5HZS/fz/C9W29SYtjq+tAFkom7Iep7qi
smxNifwJqdNroK7JZt2c+yuuLRE4owr2h8hr/vmwReJb718VeUJk7PyeWuXs8vlBcfBULC7Rsiwd
ChxV8jz2fi0Lfn9P6DYk0ywvN7SBPTu4Wq9qnW21leg/Vf6nPfTb6NcEPEeFNpyNuQMlJ6EG0zlP
ssq38vto1A4jyfvBvFb3x/0grEvJeutGotNAeqU+iBz2w/yOthfYv3tma/svQ6ujXVTLkiNJsZx0
fct2mrEsP8vtpo1I6g973iAkyQMrYQ6SwNFvTlgylg3sRPQbudyPMkLRBSe7MFEjp1F1Ddxo5aGQ
xTCS72bazeducJyLIMN1gPu8EF4HjiVa22ffruN8ErvGM9I5jJVs2K8VRWSLiCps+zBwHJ7/AznZ
YITA0QXzGSCwu3WKVrfFA0NiEnpmXVt/6/gyI8KEucsRSjEDJpwsBMTcVkXItksx4pF6FaMV+Nnz
EQF0ZWcQMtUbpRncvP4CIjX2z7lb58pycVwzblhXe5P31mB2AVWcSyrMPGq96+cNoc7ulBJlJdKJ
CgUTDlZ88cMhbF+vAHIexGU0mkVuEQ9seXn6DoiLVY06y+eFZkZNjoNkkJ/pXE7DQSgoBHfuJbDA
qoAmHymUKbtHWN56BNAIfRiIV7j52SXJ63Cw+1lLMoXIIc6w7041czZlRh6bwAlSCRq8JR/Bn6TM
jjsBFpQMA62xY/TIPnHpoc/XawLBZGx//hLGsjYHJLXGp944SbSzLkzvsTcpnQcJQyuLMG1E1rLu
NF4TRnUgGHAnuvU0L3bfyG6daRe6LkqO4f2BxXfzqVEY4pczuICzO+YwbB1pXK+UkzZkC8+m0Bar
zQkNF++jBxYpIKeBSWCksRSIHjYRM5p0vomqGg+30okXX2ENRVCiXp3lIbYT3OB9m7MSBdr/FarQ
+WVFuwT9YFACLnvTJKCkpjtKiVaOP+K3k6dHxMQK4MCeqF4PLtxTyKBoD/lkRISv55RapgxtmWCI
ZtheT/kF7Z3JwxXAINB1ntTi0UDoV8GLPaV6cfAcJmEtRtT/JdpGGDwy5EFfCPPoP4/BgGpiJT3S
Z6FdMXtKuMUFeAQ0G7e/JyWJ7gQ+NdThndhNyzMY4Q/HxMxJAVoL7y+xeiG/vcWuaBIQtY2/5ARb
q29TY2EZ+/lis1Xp/MfYbmWR5d2eUs4HlKZeVI+KtO984KZtUofx149tjLs6cTuaN0vDYalp4Eew
B9qUcqY30pIYFQ94z7YoWqE4qo6aDxXEHbJG5UrxstF/6bWq4RVtNvKvZcY2UFT3Kx9VuVqEhBiD
Z6/pAiMjTlKomuKkEoyTzKCzEh2ok7gLg2aH0vmQ/6pqADWsmfSn+22ycEKHk6FqSuPO8pvmQ8Aw
kasm95hb+pKBPl//3mbAlVIbVrtX8UGmJWUlBGIgV7l7mWm/uf7kKI6vWgh781rhRZf5apM0wS+l
QDEBhcD2cQO/ZWK2bu14vuKAP+J2abCpgGZTqmn5YXN11julFLRLklxpCXssOPvp3d9zR+5D9AGv
c/pDqXFB2qxYiQCiG+9YF3NZj4lek8BG1kPSuo+2w4icpRmyXEQ+ACLjP2OFR3/9zwf0SMZ0gDm6
ZDKHEl4bzssAp3jtxXiM0WBjF1s5wXkAMxnk+yNYcYmT+xVDqHBsayoeUe9qChpomkDFzKHXmuUc
qk6oZ/7QZ1OXxdqLMhll5NpGEoNRPDm46+uHiNQXLE07sZC7iOKy9fKXYRtUkuPpdvtN0TlL3y/q
1xl7phO0xB5n0mV8xWK9DsK8MB323JpNMTtiivOHpRxh1Du0fs+dSS8NNHz+4DtTm+UVZobMun1v
dH49nb4Pet8t4gzC5+ejTC+3hR81A735A6sKevQk9XkcEwYcht4lHTpHqCYLHNZ2QO7oZLOtOpQ+
eeenuuDLY/LYEqO20blyxuGLpiu5HsizJuo8AsaBjIKkACdMUTBnT5zwXublCr3liekMTmDw0hzF
sFirXNoGfJOSiZ8IgCsJV6ypPTl1hHOW+7elAc4uDEZQ4RMWWR0tQU/Zf2qgEXhXXqUDKXWxwvA0
z7R9+Hmg+kstdRxLuatgw+sVuldRu5Dwgp8voYjan66zFV+AFOpTfYF/BHOr3caLujHpZoAvCbTa
Zmln34t5JWnGlqV5W1Mk9e+xAN7BV3z+wthvL9u7NNQ5FxhmRHe4pvYHORRbMJDGh7glHAyEW1tC
FVm+ZYuWAR25z2pqm0hn+fBZWWDTTYM8AVAMpSsPzV7/CsTSFwosIpIAxQo8gjTjch/DqIopnhMs
2Hy3LnlhD1dn1jyH9kv+D2ALFI2Fb+caaFwRpZK8hU2f/bQ2Gs/ZGVlggD+DanL7Ekd03MTc2cDh
Ow4UpXrz3F9JEKf+udMx0Z5Btszec1kT7SEfF4yp6QN/LMH3nrV+KAd+WBHIQsvblamAFxX+X73G
nR5GxvFmbMg+49MMC8dxu1kcGKh/cph/mioA2Zw9KY4pl/wxVWpJ5gqW8n+Dt3bHTq+YLxxl++ck
ejtfaGnBRKKD2OXriW4K0asdSx5/NymltMY91XhOx1yO2GxOcN2/wNAgfxzY6CcTQl8ae4G/baNI
U1r7sWgQRXpsD6JeeF6FsV8tluLh6M3Rc4eDGQjfkh5zLK61uME3kmeJKpS7tVL5pKMfyBBoPfA1
cLFBxmMSNPYvoMUs7H5qIHET9qN8XuMtQHKPT2BSsEBc5lX7x22gQkbSHrOSZ8FpF69L6IFAaCy0
q2c8qJDCjQRSK2kEdgXEjULPSv0G8ajbGHcp1E2zEe03RzDidcqFCTdxIKybW9T6ZXn8uufVqS3K
l2SejYJoc8cutlgi+ImptEXMpykyX7AriXMSZPSltgdTrvXDDZyKmxC1OvXiBnk0lkSnZXLZ4yYV
uNn+ogBmc7NTbCUruGSlUVHaYD+GIGtGfmk7w+g2QxReI621szU2bQm35Ig3KSMN2LG5aKBdb59h
YRiTkui29hWodS70mCNoOExnjR7G2Mc8BDzDRIyqJ49CpY+0xDj+OJTPVFHC00HMrpvIq3uW/dSS
1FiKP5RADg9Q+EFnxwzRjnjju+Vvst8k6sQBavGC+qe22cdMVavTh4fhip6WZwu1kCophuVD3OeT
NRhkw+WgIa7grXousZihiv5m+GCFXIgYn3POlH7r0Bxpp+k+q9qfhstnIbAhKruDBoSCDCN5sc30
AACaTxL7OIOOyhiDflNJVe6hgPmHbtxL101yTjzGR9t/l8gg9QWamJQSp+tjOYEQUdIiE4QKPD/1
1chV3oquTzsTEx+3kR/sVLicXhkbWFrnpnXtejGh+Gi5jqZKms/fe+RHKlmewgBVz8DA5JNEiERw
gC6mFYY/N1kwJkxgLM6g/IxGq+MkQBafEyFdJdE/c/than8fAawrXwTO97QJ2oZOn/FGary4DhCV
5SWqdhCCzMIJKXOpdfdIPH4vUDD63YY+JsW/NP02aG71lQSOlk28k6TEPO7wEM/vezuVOxLwsXqH
DSo9OhDmEs7ieW34IDgN1NOIQy5/1i3ikf9dzX12maj/HaKQOTuVL5bN1bwKoYxHXXiC0hi26yf7
3JQRDuxpBKZv62JReqxIr2wDTQ0LP9W66D4/qQiP/tNxYFGQm1zz1f3EMKM1C9DQNnK2P6V/Fvz+
MGQprA3TkQYZJ/jSyq2wgAygyj6PRs65RF2zmYbiAhQEogIMMMBTKr0365tI2ERHQBAnroECrT8b
s7RSEPITUWTSeW82jnd4orhWldBOsEKY/r5RB7UDnrY/nR6BezgXUxgKwzsKNnf1cqSF4rwCAtLC
wZ7UNMRjkV4gwg+65K/T3NnuORD/wVrXPlx9tXj9Hh9FuRH3+MRQjkdX2N7CL86hF934hYZ5jzQN
hVnEriswltDyqJZrPhW3zMHxvGpkk0jOGITNHqB2zi9pjXS6CnoEGhv02n0YgFMiJtfoykX1Elwc
vv5GsbSpi6Ybg/kWFV8DsO/jB53V8x0crLJbbnnXBC8N5tlLP8GHCX91d7jC+WMXlHx7a8W6pxbQ
s+zgVLlRAoRm+UinfRJS7TGE0l0yTFF+cFcTasK7FZ7UEnyANeaAiUk+aWxzhiyD9d1yNjGNHseV
1nVaDeth231v5RBDNEGpdyZRXEjWPTK9LGOAbsnUb4yb1aIB0YTIsJVd4i4AyVi+ZXgmdA7laCAH
qNdtXQIzskUxT/JNcSgDArf7n9hQMTbtolnuf9xmAPvyc+WvOckMuuI77WEtMA3HBGZvH+IMc03B
7tqb15bqBW9+Mowg0HYmkJzIoxzez6VjLT2titRNrD7xMLTH4VV8H1xTBzFZQAcWiuplbZsg1AII
X01jmtizo6abd/AMBxexdDOT6k3yConiTlCK+t4wOnsAT9UVcvi9w+en3jmsgq9Vol1GemcIwgFq
SxX+pfpSB4LkGUUj8BfGtLyLN6XptD5UaWCiv6u0EXNLOGVdf/xhkl/Tott4RG8nNfCWDp/qVfAH
r+fIp+9h+kZVgmNgmDfF6cKnw7V3f3xB82i6t4s6yfWWOtLJKc3OF6AsFNmkZ/pspUTX/L8XMPrd
YujAdsYbpv+7s3rkClLMhntg2V0wK4MZr1mHz/mo2Vmzk7V8n7QIe7sebQTZMwO6GJ/eFdmrwJ41
zNL7I76rG+gf7SXF52QragX9l7ruIUMXl2PuwHlqZ4f3PEzqjJrzCb3TOl5Lz3Kn0lcMLFcbUAQv
hjRzse9kimqAmUJhvSsHvK47xx81FREdA6ai8gH85312lTcVPKMEt+y7IUs3aRRTo5G6lgjLd9hP
arjuPnnGgquu8KQqSH9inV+Zd9q1P46qIPmXiZaEefhbGbqBRpZPnKbJ4Nmhd2OpR6NEn7mAX58K
e4FmSJMas7WxXbkgpz4I0/s1pT0hJt1Stn8xd8o5vPEtA1TzkdFq8lv8ZBmH64F/8abcZihMg3t7
xmMSG96mCplw5mlNAeGEbZAkUlHe8VD2xXozQzZM8UE27dQ3Z/y3l8CTjQTbCnmUvowpykPkx3xy
uxJMwkrSv4C1bzvH7xmfrRkpTkVmB+vugM9cyf8p5gn3kyUT1sGZ+fAy+l9ZQXSpCoB4Z8FI+/gO
emlOEd5WAz7dgqpSWWbGPz472K9foKtTxqjiAEZEX/FRq8KSYptUeKbJmRS6/rexqFwtYbNyoNSK
kR0WHV6hs2vQDZG5M7fM0ncOARR7CSO0BCAWwRBzhTIr/P4S8muxZ117/Tmf12NDWnZXmPSRfkBw
CpxrMMY4qfq7r/UHHlGvphdIVg6kDuOvx9sh5Ne+9K/VFBGu6qG6fM2izLDQeAdCy6Clv9YQ/vcF
kHkXDb1o2a9DvhyPrKxepNJ1tPQL8CJbor/74z7TaFGXJj8xBXTBaceRQKLbzeufRCdUKsBk+Wfs
4HNzwGz6lLokMe2k/ZJzD8S2gkbpfgVCSjwvlUo564cosBMK6w/Q6X1l5dp+BMsNJJpDgPZaBolK
MgMGRk4MPkwKMlVSNOKB+gHwzVAOBP6xAMKRS7Urp7Aa6IaWOCTwr3/G7j6/MiuZn9Jjmtg8ONrm
gH3QmIKU9Q3yrb3p8BBFspGFijOEQv8UrMzZ7aQGrszYbunrhMrEBcx+HWd8NCqhp613s1i7HF7+
f2DO0pC7oAU7RWfuckT4trAFwITRy+7WNLTUPNgiOQgURa3Ch1S580ypjKEIganCRfal/amHsmQ6
chx9Qh8sNP6GO81NVLnDMFO9oywtJC+1qMjTr5ZB36JcpBgJQald7EtE6Ph6tS/RvYEABlcdoki0
spUk1dXXKSRvXNWgaTHP75aLJTH3d6uhk7QqAYmqUzikUz+KZC/C3exi/vG+ukVWOCp0rIN1tOA9
N/OzHgbiv0Ql3HjfOu0KiWPZz0eJkv1rVL/DViDdp+h4JC1hNwgG2wfqLtijOPTdqdIrHZT2YpCv
IGfOHCQZJYhQsvtIVNf8Eucqgw+d1uby7GgYsRDXSunEkgK1soapMFEGifUuaiphs/GFCCENhjYi
RlMaXQsSV+V5+lLhWr/nN05uVPFkrK0pJZ6S244SQsWo6HThzpyUxVmLwUcW4honc3sHirjoz1M+
kUl2B/9vS4Xw1fhUblr2m+wkA9ybVTuCRN6QwLdDyuHFCjbvDrUX1zV9Z12o63OJE48rr+duaqCG
tN+S+vgto+ZCsUjCzyLX4YmN5tMnXyZ+NeyX5E32Jd7kiQ3sMcGRehquLDl3QEhvoRy3pMv4/lv/
qT9eZhGLUael1OUOhCmlBOtgfUgRw1ZhsCZqDld/YWfXhonUvahtSuK1E6/faAzKuq3myvopts/9
W+cch89ISuywME64iaI5SWE7RLCe6bxj70xAO5am+Ce47ZHAoencyjBGZACoyySJ6XXto0cRnRVA
vgw1qpxpYo0opbwi5m2te3Cd9I0etDf3OgXX+KQcgXbuAp12WsEj0HPHx0EGr/OvedhMPvu+UFJY
Y00xNxxpTEAab2gOyXn7gLKbyDmabntPttO/7z3YxUW/xdL8i1/WdoIzySngZ5khQ9XQZTfcOW3F
Cb1xcneqz3dy5WjjeyuEJ6ZEr2jei+parBjmtFbgQ5x5TUneCPswxIWmX3o7ksJorW1zjP6dyFFB
L+ZYFon8fF+mNbS5cHEBzAzNAwz1/b69ASrjh4XDm86/OlDO7qH3Wf8esuHB6+OmggDZxInQzYol
rlk0c02PcDshzSZpn25VmeGrp9GxB38bjj05VhRttzquN/uS/PCj8xdhKKqVfLGA6QIzSr3Tf12R
We/+2VEhvGnB05KY22sFuvnEIKcWvTjYuy0N2fY8YFh1iv8B/YS0mutKo8XVZrW8j08LUUMwIHu9
eY8Sf0qro2tvltXW0Ochfhtq4z8HzLLj4SelezmUVwWPpf5hJjkV/EdxsslG4OGK9xrDQiXm1HeT
3TWrwiYrhH0qReAWCxiIZh9TqK6/x7CJu+3rJxci8GP1dFsO64lROkQ9/2xd7nNheLbCaAauduiC
N92tNi26mp+XtaMW7N9tL04x+f9cTGZhSS9oYuV8wSMkei9S/t0vaJgWsuArUEAj0bKcwaWz8pqn
t2kllf5WbNDwdcnFb9UIk6iU0Y+wJOQ5zisMbXZU071QRMvUSkuRrDiRiA7coSs8FAkEa+UU+h72
o+I6/D2+jZCJVtbVpRs5rUemg4k94UQZSIETgBNhhSZAsYlc7/49A/Dof3sPz3rw9mbm2p/NSeXE
Fb+RAD5qXJ+o4Qn98x+smpUpzcnc3P9ZBG53KXShHnmXuKcLyalhSKz9kbQUHja7Xwrka4bBZHA/
jiEwGOeLcByn6G2Y2+BAJRjavY3yfZynwC6oUX2hwpAuAKscfiLaAJqtCy9huCUh9BAC4rO96G4D
Hr+siOxb2qoOTrfZL47nPrJEAu3+YuhSWH6jZS9idgCn3MQQMZajruk6FfWh+twnGgQoiM4HaJl0
a9CyuudtaP3NxEEsSQCBtOTm1zEMrF4ormBA3dIrCYpyL0uxmNxblQiArHg2WUfIAdqoxV5XWBdk
HuqmLcKaExf935jZsm03seLj2NB14SNgZxtsebfKL7fE/gbuUNU0jJ3UcJjFAsIg7EpjdC5rgZoE
UWzwKGxMFRI/K3WAuYTYyd+oVgvKB2v7soILxsHMSRg9runj7UsJmQkH3/6nrDMfBgm+pVLdk94n
D2fS67ON8haF+ovbSm0jg3MpWYyrbgNWMAyPOxcVxeU2A3UOXxN5qsPWpEk7ZVF6novarXiR+BAJ
KCLkF6dzaZwMqlPi1XYPVTZMRiS1iMlmCf8OTx8Jup2y6m1gIQMdqkanzs0XOQL7R87/B8IKUPvy
xltyaR1hsdosv++nFGec1/LEKxURlPm6OCl/MuabrQsfMXKx+AtVMiiN8UnM2ZdNbns7ZUpoWpfE
18flyWcdRkYaJuqW9fv5GS7ErudrDxoJlxe7gzTfii2GjWhwBOzq+n8rJ/hWLU8GS49TZyghdgnS
y71wIf8SL64dLsgxF/2TSFHVSEDSC4I2vC68CA1TqYGHjx4mEJZFEIQzEUTsEq+fwlLVB5Gr+8Z6
90NvIFHuOQw7gxIJlq33CRir7UX00Y+5NxmTNmocVkTdJkU2A94tiTruy0+9LTRuaAV2egMkW/OE
/lGWSD/H+sLrx1+G1kI8pBoWfQtnEUOGMO5hwhKeQ4TTOhOJ6hxJvQvlwws7fvjZbk/U5tZPFnRR
aPxK+TEAm11YjABBQyPZwxKhnYS+nDr40nAEi7xFCalh1I0ug10O7UPNqY875FU+GHvFmjoieQzy
XrzSmRvM2KB9PFkqZrf9CeHPZtEp8Y8aTJhUu1yUfzakLymGmjygbxaX4bpUYF3xiKkntSytIIw6
xcF9Fk+hMSX2R+EfdF5u13lCV9AspxIUgOVGbn3mBDSArjFnedROiDhsVzyNoNwShLvt1JjIX+Md
JWW+JiavYwZ3o8TsSpxvdvi3saY0vPm6KI6oo26Bf6Hj2FsAqzzsz+PUlcCQ7q8nj2YhT+oAUPpI
0A5jBVnIbO2U2t7Zy5W1iSDpzWln1ijhwBWqI4AHaTZK3HlmLqbRWk2weMDtuNR81lSZ3g2/xjqn
sf+3Wpk0L3VFx0Z5JvOYuJGsayDXKYbCt4CZ3jjG6frbZkE2MvSkYjnNG9jQldW2Ncj+pepTQygC
ynJvgOOUmNyd9mqzunDLa7dsy3H0pd+m1m+hpabNCxq/M5ZkoRYa07xUFhmi3U+/FuwNgGq7OmjX
nZkZH0b6TWdGmqBF6581qa9svnxUAWC+m7nAUseX12j4X8pGBkmB7j6z5bk1BJC9IpqndvpXvZCa
bo6nNpn9WMfn7JTB7KEwBGcl9rZFVKokdjWqzfcjcBJ3s85BLyaXMKcrtADNaYTr4CUwJmHBXbsI
cBU8VoPusa+iRq2NnsJlIm8ftNoac97X2cbtn8W0VIvC2qweWxvDM2/Ltsduc5/F+jpWkjuSiM4j
KWhBCoxzU2Yq2ZJHCG8uNmMKuG8ue0B5N6aR4shV+wWqpN8vgipKnLc4jEg2XOQf84IbxXnt/hN1
BuV0mQQBSeoNKf0peFpSTZUz0pz0eGH7g268B7pLSFQ5FlleNCsW+kLiQe4pSO7WYSp7t09z+pff
g1RWBwrV88yMbd0ojuXUhBrX3eGKAuRQVW4mFQoBidAfP5Q7jp66x8/0gfvEPlpGP7cJNLBh4bn+
pXcj/bThIH/dV38WqgzMbXliaxbuI+mTqnxIAi9mecWK/ibpzttR+jSKJoe2V54gYh4cLc4cygxP
XNoQS7XC3juR+3wqS7FGoDKnoAK/R5fJtN7FqgdGgva4myXhUqYXOIiXXBDowa+QLFfuJlbTSVkY
LydFYRrvnR47OLO7Ewx0dq5CelZt/2kXQrjaY/xxHn4ixrkwFE/Xfp56gQtN0d26WuGEF4EX/93G
NpMY47A45kiC5F0K5fmU3QiUDFdZghzFfGk3R2v4BLwPUfflyhEfTYBnG2B9xNEh4SGvFGi+MAwv
xcaSYvRXd42RFl0wQIMp5R7ucEGmDPwcJdEUxTiCw6wwfK9raTh5i0kFPN/xYZV9cswIHZ3p70Z5
Daj8/U7sYczaph7Yq2ZjY5YrGLo8dm/zZfZ5sBoNPERYjdGD50yj3FnVJqF0Q3YLqPFoMYqTTIgR
Y2KymZDtBhoEmDC3kg9Aqgf/CWuKI9u9PvdH1cnNAA2EqBBOXxkFUE815czEDWQfHxA9N/LW3K4d
yC9qIVrbFVL1YcEjE1dFp1/AsfAgj1qWPCBhc9nu5/OoEZObVn08XONrCqa/WXNxJ1ea/y9y/xpY
B7kj1yC+uc+/9FAZcnKOTKq3IbgbIrwdw0lROde3pv8lIuZWM3/t0iKWYYpD5bdaqMf88qlQIjVQ
P+9dFYsC+xl2u+/LoDalAiu3ZjByKtV2lT7hJtqUyqqQpOe/+E44aZtsAUAQyKJomsSjUVBeyraj
bGI9Sbrn4ipQoSMMLaq2FXFKw+zERDTiOuKcBz821QAAGcWOU2hQlMqpEXLtafOKabF+vOUlgc6B
AbJ/uapxSTUuOK9P/IzQP+Sf8YZfPo6ErY55KreKmNI8Alg5weJPybHkPCybcJ199WqhBH8ws+Kt
+5nIkFbiGr6uW2grZ6jrmfRukOfjOTgAHG/ypIb3FAajCzt441rhU9JqliVCp4nJmektOB2WlRU5
5FKRdTTfNES3Iel5dw2P/ZstHka0nRIERdVaPLDp7AnxoXZSD06cMaqumjlrCMdjec+rlbYBJ33s
1aZqj5SflBMC9Km8T/8TQUjR3bFQed6E+G50tqfKQneQzZ5e1RJzn14XJ2SJkn9GN+mp8pokbfhC
7t8OQMk/numLW4abFhAHgoqmv4fFdWW74z/oEp5sNBKmLtrzbYTePC94hanJdIjDz03XG+p7UuZW
/hFRQihys3E52tZJ41x3J3spO4YDq4G49KEy+phRDlnjvNG2OZBGbHDMX5n279vEeSFV6ik7sfR/
eL0MIAuSkpAv3mrpmg1xbLtljz5FYeT/SImfmx9XbR38DJ0P/QGpt5RkLH57pBq0llmLQkphscVh
ZEA0uzWPzfKL6uWfgWk0XrW4LT8Nt+sI8B350qjQNyzEg+cu6eTzx2Ju/HGeUjCslwUX5Y7RQrwt
lhJMifVxsI1E+OKGr5lIh7uIB/tqdO+rThYzcpkVMZH5xwrMVN051lkns2ri0W5oqV22IcB5UH13
QGFPwpnCoIDGJ4igkED4cQ/UZWRPeYUQVhYIp+O3FriDhC0oQnN5HBDPLir5vUN6qj0QJL2sK2TE
84JJWClNXJbBoo4Rwl6a6Kz40DvOFLGl31zaW2WifkJOUjVLsL22dBnifHV/1QuhUfHjvub5qJbu
zCBlDGFLXkRbpaIYiZXPA7ywKSskTx/Kl8wr+y0IPHVlOBIuoF90ZttZqN+0+mrCwBHIETg+46pF
ssr8vEfZRkcg6ma/EZ4ilO+epgstLCgDj6rtV3hjbASu8mf/GBqp6kF4WvBbp1Qzc/pZjlJU5OiA
EnUfBTnpaKhiJVR2BieXNs6M2K+eGxEq2mnHkemfSw8u9r+Vc9BBfmwXiTrOmCMK8xQeQosaPS0Q
ZIVtSHvZY5W315nLugrw76IjVMTagKPYoV2Iegsthlb9l1HrnoqgBKV2a5d+snUp+vz7YxfpvjVu
hvU6fes6NEK84QmTR+f9QemrttLf1GNH6B3zY9ff7LZZDqbQiOvODrG0HPrIDv0Bu1+eg8wfQ1b7
no4Qt+kf2mpv6VxGcUbrZD1zf1yEP6Zz0qEmDoNbReSnBdaGXiK9wOPgy6SR07qLOo7uPC0yHfVq
DGy2LrPKx+1od+ORcKVroou/IfqzMrPGN7RSFhlKXYBg8xQeGrej5H1XzgWawGDnlMw5rgYmBNe9
BJVv4lFnq0cNhaWpi1lWmSnvVoybpWuM7VoKv8OZDQqGyPTUuGwQfr+f8mingfoQB+uY30bR+zAi
XhSk5itKvdaLE+GlLYJWXeCv2SGdWCrBS2LDy+5hYqE0lSaW6vu8wdmyiTlguI8sqrfjlgCfX8sT
lCZbMjDCym8mh8+YYRKACh2WnJtV93C5vFevRPYvxQ4G6e8IBBcrwxb2KyS8yEdxAm4FohgJiRtx
oef1aLkAoGiwKstF/fmJDOciz838HpJiIxfIDdWMINRTlnCn6VsZ+5bu/vv5mWEGI5MV9tfY/Wf/
JppW8nxLrFQcGa0Dg3A3kUjx7R3fIAE73VR3z+pZT8AVMdtY8kjXVm09u6etvS+M+iexIEQQ7KLM
7pEBz9wSSwbP/gpUFpcI23BlDHqGdiba/97ngl4MJTx9Y2vjkh8jgeTFFkdKwCC0OGCzrVRygUAo
Z/pDg267wv225jGBTM3QYuSY+hKbkMn6/U2BfvIpfDsQvq8rQGF3nlWj9K//IcA7DZOxKLcVf5wy
8CK9PCGGKDYjt66S/zXAUojJILF9CRZEvKBMtnbMfvcb64sgSXIu2eCUUGIXaNwmVGXCtVNlVAIo
CZN0li82AFXFPxuNW6x93Z1SPyiz6Jv6zEXSjJeFZ9Gcu1KQqnl/E3sm0r44LhfY1zs+LXDdAN7n
a7WFGC/Y0nlz4mHYD0GYfzG9xChwQWENpqMIf7UiNRVJb+TRAQdkTGKH1NPnkPtuo2dokW1QFpis
WcC0k62Yn8ZAhECH/LdDdsoTfOSEdKeAx798YiGU/jHjPBHb8U1OKwSdIVfzyFeNWelAxKC/524h
pNm1Uh4naOfvZtYt8oIWVbBtXEB5JTaVq5alzVJkxs9R/4BbFmVFLoKZyZVZRj7ofPPtwfy0sJ6t
2G0YFfn4vZ59OLUyTut0wJxkwJiVLIO7QwVcwdJLFC4LH3Y0F2Q1Zr1+zHwb4Sv0pX0HR5UdLt8y
ZLMrvFmr0dteM+pMUVQYaKS1EAN0GFe967KDrQiVjfDOCNxA1i7MZwJXDlbUx/jAcD5ElsdMGf0s
Tt3t8MVCc0JJw4Za6f/9EkA00af+x6owiZOsc8s1+8SkCcaFPYF3R06bB7eMmdDHNsKhtg7riyGB
NeGfbDQZfMfyfcS4efb9SnNjBFhyC6oqQW9+Q7p/G1f8Xr4H47uuGrOp8xXGukEc0PXF8WImo0kv
HgQr/UDtTBwJrYBrAseI9NI9bCVLJFgtUlxYngNtZEQAbyjWltPv1VH9EuvOQ39F4gd3+E0RZA7M
kehltlRrpgpk7Ke4hsrkEwQZXcrCwh45tIixus5m1GiBk008JaQRuejjZzpn4fR2exQc8sBmk6ht
19GUHHQ0e+B8K1HUA4kJ2hoKv/gPfwDRBdA6MWA+0K7RibITVUM0uKDkx05jRsGeNSujLdmsbJir
4fxPgPw4TkOSuXwu9TVSDrYl0s9KkpziysUnk//x79qsQP82ZSw7ICdtyqbR3FIOIfRvuvWM0ccs
Yg19HYNcwYB0TtjXiKjx6Ekp4+H7Qb6NFFRJTBLAT1NhnVYtnXzck2AmSejyeck9m8kiZPkkn5/B
Tim6q+KBQ2hVH7Fz30VoZ0Zkv3sUJM0wStyLrnaJtQi7mxJNsw28o886nQToAdrcFg9mFyx5Z2vN
KiuBF+yQkgxXpxUgCWE6YI9vIp32G9E/y0EtKrzhA7ZeEx7LBsmFsSeR859yZ62Au7vGno5Ivmtj
r1smgy4gBPP07Lh2Pn2b44GwQcx2olfa/truNYILOQE1c+eHEwdVcjhjwWSWurJhrbXmLTGdc5Gk
UiTkxG/KaWftWo8M0F1xcJepFGC1l+aq9bEuMz4Nied+vW4adQdvHt0zdKmwPc3EBZXak9/r3gIv
BHj+ritulPE99EF0WBjplu/KtyGJTtV7Mhecfnkb2YyCHLaXpIgbxTc7xL3koHM/2Gwrm0/QLbjY
lfl95ZJvw8IwVEaw7TvNduxULirgaqPNjd//VlFZSbFrCWRMGQbSFwFCy+9w25bgVmnEjrFiUIgM
ZaH2PzJPPthhrTPhmu6OUCSBDLSfZQaEEJ4W40YRkeapc/DHhP89wnUMqBJaLbRbZaIVRIR/EByZ
op1A4DicT7dY0KgzEckvGknEVGd6kWbHSk5Kfeczuca1/MmhOMXhlmFwX2h1TTTrLqHPG8mjOnjf
Wmz/sMs6FDkLz9gAapU6Vi83Q7sUe5iLGhNnWwWAxowDJT7QndCalZ+N4l8DxpfTmwP21Gcb5889
q+PeKVg1FZE71o+YAnSQCCE94s9wzW/PyocklhYsISd0ZlmktgJQUNnf6QhZQbR8mekajFf+yNiI
KMboHJWAk/ZA+UDPe8Q8LWCLNgW2UvVj8OQqKV2q9utSirgAJ+kxaBTA2cKKBpUEscW57fggK2O+
AvwjVVN1r8D2wynsmTy7uq9uC/QoBaGHkLGFxr6WXthttAOOnRsFCgeRgO3xYdUUKUseT2u7V9sG
fGQBmYOQb0IYbsngGqN4pQLCEAJWDuM8ayoBy5ulKE+4rvMhLwL8tlsUF1cgmjlXoeG8UGUygOXs
+lLJIqWkObQ23yORwWvdAmPBa+/Kdt5Hh3p7RqDzhxlo4DESoaqqKBcuS+pCRHatdMfu7LN3GlEH
+xqyrliaakvOebaW82LiZDFTzm+HnYXR4oddYWUGuOHBb2+Fbi/kPNPpaekFsibbu2Kw5oA2eNLG
/f6VjtGqSfm7lrJG31PvfkoI/nEEYBuucQjKJfw2LKVosMpI8cIgY4y06LSNtShklbFd2A+IzTty
k0q2InpO5Ug7fWm+SjKnDhXacrTj02a+pBWBHb4XQzE1gMf583l/AW7IbYpCM0URrkNVaG0yQ3ql
BNDOIpk2+blXQ48Py4rHnfY/J5RVHgDlkkUoOM2WLsDfQqRyngmZuS7lrcPzPaawXxcEYdDGGbQf
QyhDcDPDnb+gL1OEz0iZI7Zi1e/GAPxbKrCnTBInjShSsy6Slu7d89AG9gkaLbdiRaO7oX+zzz1b
I/0SReI8fh8bKu1OYbPs2/oyROtg6i1/Lk+MgzYWXkXkL8EHJFU2U/l4x5zDqVLdA0ueeovG8Ikj
SDLqCrw8oal+NAKxBlCmoP2/STzczj7TodX+yjw/fnG3JBEJiUScDsbWJpqtXhiwnnxuBzT3drPt
W5/T5pYv6RJwATIhVc6ZIx7NkchEQ3MX06zAfX7Mw0ToHN41z2DQBhMtdC+tIKA9i9k1NPzfXq8h
9hJj/CJzktiizPsgqgst18Xv+O0CBqTsDbfxZcjb5Gyd4V7PxSrstOs4MqaAJDIHoede0eyEAeOU
o/iP1QL5g1SqsSrfF99dC4VSUtnBz4fU6Xm3ClpOt6XO8e9/W2aa6ryUCxzNCn5lBEgXC6Kgn8so
kym86ApRjDvXnMR7KWUKrixvYWkf1m1B8URvbK7qc062LfMdbdzqVpJgtvN2a5+ph+ngEMYGF3iz
pbV61gxLv1hOeVTGwXgHD5gVen1adyBRcSQC6qUXIG2C3vYnBVUNjiwRDUwaMhcavOznGH7VsyNv
b4SfZUPywI4otm77mVGN6Mojc0roAulhnDSXsTHEXuzcJBaAnsibub/pA7+Zt47rR/oj8u+++RMG
DlAw8jnI8E4XqieksHvIajaDS/8G1LlxQ6ehydn3Ay/DFDuX1YgVDKOSPjP46pGw/MinSN4wBV7P
9Ntu3MGYA3oNeyjuoWWjKGjfnO116CHV0ekkL+1AYYjeZeiedwonP7+h/IKufNGM9+Kmvl8pEYzB
yQySoC5VU2jRDriMYuVNVzWWyRYlLvmOHklvibGkBr/KBwu7UmGhHy+G7ObXUokRL4QuN3KRbD7O
Pzkc4U62owkACQ87jfhG9g/ET5SryLc5NwGRFsY79QMkGicKeXlp5xUFdbsYQqgx3PNs85LU0tHx
wiojVjM6kQMafIWyshDlv9uuu1dHqUDJMEVXVFT2m4JSJM5OHaD6LxogV4o0Gd1/3MQNmIKUcsVv
3EzU9/sERxH9RNIYmMZmB8gJR+70wvWV+xbCQ73CA6TsaO2SIAc0b42wmkE617wn96IpsJGOZGgj
LRBfXZ5YUbe3FaaDq+H1VHqUfM6OCnlanCjcrHrQrl0/6468haYGt/rZ8KtOu5r0wOPQ5Cx0QgBA
21m+cz9Cwgjp446voI1gtcdQasKrWdEIzaT3asyjKtYegZc9vUKGZnlK/ThRyfL05MuswV1OIdHG
GG/Ir8bCR8OLcGZUUELWP4fOq5SuTcc0RUXpu10j0eAN26iFs0bblNiSlrw5yciqnVp+6/kLsDks
lYx1tsdG9x6w552oTkd2WGDHULB7b00NT5lwa/gZmooko6cuyp4H2v64bCUjdtOpttgb5+k1gsZf
IGXqrp//rObCihVkj2YtbupCNVdv51zLw/F6LmIZrRShGUkLZgacPQckR9hOzOUgE96hC0lxwpFj
jBnrDvGvp4ZsJUC4pD/ivmLEz/lrXjxJVILxAe2cq/uoQ1qolLLVhLRKnkwJwgtJ+FAlRjqXrtie
gp6qvArwEn6n62vJg4c/9BPkEz9f7SHUeEwWjIndPvehkLSEW9mfclMMtt6jlP7FY/uPL1HIpZtq
Wvs0WPKw8fVnwidx/YmM+3yTsK2qXoKefq9fz1u2OzMh+a//qQL/5GSYpoHEFIqBUgIk6ktOdDB9
fpNlIoLvOLDmsfEVrPA0PNvOOmMZOddDCed84xteuOgytWfKCsPA6pN8RhK1WZqrDEBSSwA5Wd4l
z1XejY2PnAwFexAMALuCesjhS+83ZKfZX8K5ssc1I3jA5zSfrJQpIKSQfQ6ssl7X6OwXXAkwX6/p
9ks3KhAor3t1W6D0Jptaf5XPe/9nZrYlOw64mzSVw/pmhn87jLShLQvybQf9WQ1n7m7+u2egbI3d
UR7POhw8o16DMn2nORR5wsmqxaUZxIRZmlrai1nGVuMFLM0yTT8Iu3cZ3rrQLPah0PdRhtcNszMS
L4wuv8NrmtcgttW7KNEcRhLX91xlYaQfMvbj9WaeWZ7kiJJcgfZ4o5YeYlQQqlJ8DCdtCWpT0euj
/SbkdagfAJmhAk1uiVd7h8os4m8D2v39WofpNBTPJJLzZ+ChROm9oDMpokf8VDv8GpkP5ncC9kx4
nEYtlcu4Fmy/B0ncL1aK/7TtNh6iJMQ4L4d0k1UykIMHcXi00Gsq52J6HbXewLJIxrNw6/4XhyEi
LdEuxg8k8O00eIkWIA9gjnZCXIkebJqimqEP0/aVoFmzgA95dSz+lMoh7Z8v3ObP8yjA6xzIgFpf
lPB3VFvfvvO5s2tX1gms7lJifiEEGKXBnHyJPYJIeFU71tLHXvK/7f7ZZEUZh5y3Pl2Np6cZi6e5
Lhor3CSIAv2RYjCxc13N4ZrP4tdRttH6f/7BaOad8KRuKbzebIO0gevnCj6pScCzNA0WssHlS2H9
gT53D8cZO3hZUoOBya1ffzakUNygkrcc7Bhlw6OqI9iCYlDsgdb8RCqyLqTu9f4vWsyqXZRC9JeX
uX1LP6kbnOi7DOJmkY9C634ZYuSYOc3qyLuYWVo0ItL/lxns+B9ow+8IH1JzdGlQ3EV3v4emOffh
wC2PA19E/PJfBuMhb0AcykuKKk77jkD9T2ofJq6k9pEV0m8YuRPob1BOoNbNQd5/m9yyCOTjqyU3
GJMgnaMP2oCj+IW6Y0mEonKw5FycKtYFH31Tmg2gvvYhcYhxg2/7LGZFv3kMlHGl3yeGl+fMfN+u
6NmtuI4ZGrEgIRIOhRlubHAXEw3XyY62LTkJfS74ovmbyDv7PxAuGTqLO/bgl5zbCtDNTejha4rw
onW+gakhwbRvfVrgmlCM7KH8ag97KOp/tFX8aOHr4AfpOm4wnpK7wmp2jqj5NKpNgK1qNaW8sZHz
gH/41dw0SBhLw+zcniaRXzD3CqPffG7zgRwu18goPpnKS1cHABM5QweEbi+vtrAOQh+5hiutOt6t
jXzweopufR2UfyDMsEvdl0Qkp51UfKHtW27+qpU6NXL+DQpaTOX7/l4nIP2461U7kmIUyVSRUZ86
fizFkDXAXA8dUSYicqQaLUlRvgV7KcUJl8TQwOTpkD5dVfvJsQ2vH6RMG4tm+bDywZw6uQxg4b3J
MOubAoo42RysSQf5QUCDwody8raFZ13M9IOOBbZIIbkqrX5ppdfgo0D3uw1FH2nMPchEgbTKStxp
M+cqFwP4av49PWJkgZfzqyFqW5R9CmiC/5M6R1psCprekjUj3oYTH5mOS8maiU6BsDZCwG9fdPLe
yMnfL8uMIC+rEj4oq2i24xUlFZ0iFl8SFS1qRPSXFnjDYTb0SpdotZzYs7bCcsi7XWbIIH5Q7Mdm
Op0dde/BsGR4nh20JMR2CEqBHOBjLW7ViHOUBtcfHbxU2vkr1jyMw1DL2hbzlDFPzJkBXesAA1Xs
9gg6ZKy8NMuVWHgzSBm6W8Yvj13AevwPKFOYSH0+TCvwEpd2G+QcaPjfHos0SiSDVsgRviDdwqIK
6VsgpmzgCW5hk3Y/wbFOD5dcWGV+CY5mgHh6+3NSYhgoh5FQAthvVr0gqWrrit4vvzSYvkoUISi2
dE5mHCwYVCZA90zanN0e223yvVAj4VLzvfYdSIRUAJpYLwHSAmqw967qz0pQq9EgRE4sV9//yxJC
w4wouQ8avM7Opr/Bcr34CC3KfX+XFY2BhAPkQnUEe/4bKxqw5NoMq3HomO+TGx1xoLD7ChJjijSt
a9oFsow6WMZXUBQQ1IwFmFG0jAXvaN4J/hGT93fU4dy6UxPg3ilIsieQKyeR8m9j7IJuNJm7ImdH
PUFHkHSElQZ4I+/YGq6BaLDj28h8c1cqzqRU69qKm1fgfj+vgKvENfhAi/2vSptytMD1yj1qPLZK
LorpPO5luFcN/yIzONKFs5wCFOVsx661jE5Q0nfAFwQLR0wUBpJAxQdYXcT2MH8lc6iLkTMsz/K6
r9n9gMoK3q1muD1T/hPH9fm9Km0i0Yh6phLWYyWkEqgOcmcr1TRbAdmUhtQpZ0PPZ4tOvxyAYXII
rrkORZzoxXrZpzzZ5Uy+QSJ/qCrDJq+jsjG31cNorh1Jw7rU81Ng6/gkU3Ppc1kNkkVzvIW64oP/
ewZMkBgrsczGlLmVIyynlYmAFmQsla7/eYsOehhtexuMbFTVOkA2Q2pYtp7nTs4l+9zQJWJ2ozTB
PZmjGp0lgAf+8fzTcJtMypX1A3KTmbeIQjZp0HpREkgM+lTEa2ySN9d+ftDII+vA0mTrrSqRMjFG
/9xyAlQy7bUcgYYNcTKGN0i8gNt0yU/yJj34l4cYfPe/bDouxL6ewmCRHhVvv1q+IrfoHGfjcH12
OAk8jhYSxNZRqgNdcHO0aenbUYZJjBqLgyOICRi2FsVyPO+Z7qhdTuJjwhrnFuya2Fm2sU5tXqRE
aqi4uer2WyEJBzaSyUxRH36/YWF5B/fF50i56lLc1anZI35Uc9hiofWc1Gewhmth+jwAl7WhiZ9e
/T1VLqtUNMS9w6w9gt8Osn+ftFcVcGneXEJxnyxkn6OB5Nl/7QAYxJmWmqxYJycwpCaDYCDFV6He
RZ5c5p0Rs4bpJ5Id2ReUNrbKdH1hIeCKLqFgPh2A27/U6z9nCBO4osK4ljsN4i/fMYjvseP0nC0d
KpQvOFfUcYD4Xn6MTzqF2EkJwhFIcoa8/O50PQoIePo3k/S+AATglAwkHZ6uFjCPagGV+FMH+W5X
tILzHZjV/h6ddTkBAu5RImyj/xhe91XoEml5obqNo6B0Zeq6P0qw1J9afUH9fSUeOm3YXe3Uff5N
z95Vf0sknPt/P2fkk2Do1Vn3ke/QmZ9pseUM9/ZebyFynSpJOLnwv96PyxgiQYpnM+CjQcvCwi3v
d2k6PrKgI8wylsZW5zJ/0zaAtfoxe0AfY0gBYbESlTAkFTGZTrwoWAHQ5Xcg8jCOkOOOOTJI8ItX
DNTlhPOYoP66ZqNxzTGBSDwoSJ1eM3WC3wtOWxph6W7LOI2Ps4vwiC+AvjQUqkUM5m6cwKtquu6/
yINjlzLJXoIrFozpI1Eq2qjVDZHOJgQt2i+umTqB1lrjSBLEygRGf/pEEp+/Hr7G4tmAvsuiVpvI
z6RV/VHihS0x/6FyKTK56Lm7+pQyMWyHErrPjbzSXltFLCffDo7odZuCbhd8koIinae0WJsSakLn
fx4sCXTtQDjzX7bBXhz0oNCeDenBtdlaYXZf+pkz9P5d8cF7aA61r7lKVAWefbryijYG7FrkmeIN
lgLLO6PiJ9hyK2M1dsfBCUVL9H/KIUOdbhmNvEN1HqWbNP81i8w/ulmz3ZIECOIK0wL2yfKy/AYn
YqlQxWzcZIunWvZjY9hGtJV64KuA1FzRfXAQ4U1TyIoN/dBCNfksbK7JX2CHa94/mbaLXfJEjhu6
c2ag2fnW+BdEJT/TR8qyHX9DSL8nIHYudZHZF13R22QyU12k/vMlZxxwnAWsb2cSLVNbcWC58NgE
4czstXF847StpoUpCf7yq/WWaVyKyD56qbcGqkNnT4R4SL+gb0tqTFDLbKanHcIfxJyz23FGroy4
sKbpo0kW+dNIqRyprNspLryuAtWAmW40m4cOYO9B0XHHQXiHSaO8lEshiCRWhQY2B9YhljtndON4
A3nTKe7ghY+vng5SwNLRchl8oIdgujoyspfM1teY4Jn0G2kb68Llnkj1gZrj1suO2mgicjZK8Wn/
opGp2ibcsVdB+a3PMq9BZnlS80B+manc3hbCx43xKWqoTRTHeaCcC4mXHAqk7lyTlwQXNJDMk4bA
ynPSywvBTe88/L5Ajvnz10c9vHqezujyI+j6V2ux1Zk4CRO3Lrv34X+3lneqsdHvFYoB+dx7SVoV
pT3JTOzf2H+JuH5NMgsycv7ewelBdDMRCXTs1KIMLLIgPCP+LcBp48iFgGDVHPDdmPCFvaq9f2XC
xnfslwgOwDLDUnKrabhqiiHNOJtsTpbDRg2gKUslRbo51p9q0ir5V1IBLfwERynaZviJ6nWygO2c
FQS1n0ntI9BqGrsYJk9dlg8IRgF/VkRV3DnmY3iDCe916wVWhgWxpmHBCp2srpNu1QjOCbPFMLZq
iAa3PM+fQZ1iMKUjWii3iJRsbSQp8fA0RGTv6neDH/AwGVZZPG6UtVt+HvHc0pGB7suYRRw7H+Zb
SNGHqUJ0lRIz+BzwrL6XjRjHXxqUV9/fyvi0i6sf+pSFRRBz7xn6Qf3MNT7/XtkILPFGaDC32fJJ
2WPz2lpbyjkkAmLOBH6RfbRMV4mmfz+42Ly86UtPTsRsOnWl1SXfPKZ7j7ml+Vip8cft/EtXiXkg
olvjCRJFZTy9j2e0CTJaU5WzciUd1RYazcEZBPZirmfRqnysDG1o/5RZalV3pTA1lthcey61Q9PJ
kVFl9iX0VFe/qPjtTO9iqsY5bu4++GCalyHrV3i2NhzWkrPlXE0Wlmdw2aQNclcWeI8oS0SLo5EA
NsgSiWZ5Gt8R9EVZM9mH7T3Jb+pAQPO8HG81KnbeM8pWQ7d3MWIpkAF11RE1mDJgD7X5cnQxuhJU
td8ZPrKYCqGoSc36rbEnHO097jeeqGIRuP5FUWuRi7lMrjpQsVczbPqE3XZ422Sitvmf1XOmC4Os
cwjmvgrys+kYQ7zAi62jVFqpvFiuMy7qSlc10MBIvn3rv7GltLevMd9AO5l14cMBT91Q7KyOAhZ9
/ni6+UYdaocTFb7tQOZnzUSX91TyTLsiQhGz/Il+HObiMGNGYgduLazdkSAVjOMNUQAjrxJsKbCn
oCB52zIt5YtaXvxFa5YvwVUvwlvEmwgaGM6x6gfWJGRVo3pcoiMfNkLvwfPTChcVzvIi5asnkel2
ud8xFTVYO+LfjUzfqMpgtGzyUYCHKu0F1QqQorve/3FRwNGEoXKOf1Lm6R30X35Qu+k4C3nPilwf
YXnSxy02NiSRICI05gdOWd8vAmtkGCmxoP6mP1WcxFtkVbxkRreWUDO2sMFgVGOarYFInYgXrpET
ciy2e3RupE7fMh+x9FCMOiMU9O5whyZ06lwJ1r3NllhySx7KEDcZvHVvRdga5+OV1cpAE08kbgbX
n03w2p6o1c1xgNCCxASNFiINypaBUCCUDX1hXgp7xf6XEBG5DNzY50CJR7TFOr/yt4zo1qK8bbOX
UTgl8jFlFxdNKbHycZyHY5uT/fomMrL0qbvhJ1r28Ez2AjT3NG+2VW7vpFbkNfvTPMydB9OtuPP/
8eWZUvUtObTU8U/7huPJfnzGJVjtM6tlT09xHXTVUdsWloITDrmP759WAJNP1u40k1sAH/KQI+kK
YOOW+/bB0CWkyZM3IOhFjulnNTdtB4DG8zKJICAHCQ9eSvWjSr76uOVkz0nj+MRtzuW+taEoraDT
UmaNsHRpxm1d2GTpCEJvwCnVWtR+D/TV0sannFcgUm7yCQbEbDQ+hPNbEUnsXj15ZgoKERj0ndsH
xVwNlomJQRCdm9Q2wU+MFOT8C1ALy/jdcdYfxlBrfWQMMgCiGbcayuSoEQ3NMFZsFD7a++/qb+dI
R79VBgonJKhBoAypBXQRMWtRfI+WNhYsXwI+WyBSDZQbtU/kHuK5B8PM/cUyU58AjkuXeumnrZlY
RHNQjNi7ow9hob3Z1xu9lGn4ui1qyC4mAHpJxkbOPc17TJJHUtwaaLWLf9wqyCelSRpnRZX6JqJp
fWH8IbBX1xNXSMBfAZOik+Cimg8aMd5oYK7betQ2sediPDvBOBbJqHCLcwH9YrnueeMqsnAYr/3m
THoY/UGWLj7bYUQqpqYuH+Vc1B2cJc2FXZrI8ksvy8XkzObafeyRmegw0vDPeV4bMz4YoONXa60h
o3OVNCjbJ1bZowJviUplwXXnPAiQZcNvAME55KCF4xfvDdRnFNoB8DdvC58nLhwc6pLx9V8PNhYW
iN+0gsWarf6EvwmngNn9+HpdzbWaJfHqzE2m0gt761NFEZux83FOzKPq0CMvrhUdL6DC583qyHwK
kEdlWydlYKEWTtfuBGcCfcNg1r/8gWG0JGV3pXf1CULJA7D5eMFwvZLTkGvSO5MuOhZ/8hnw4l+b
ESwFM1a00l+q+htVb2FWXO3o34lbKCifLsh5QNzBI7RceC0soKy8lkNaZ/NvKH2N5OxvA8mD17uR
soIQ/wGpY4n8/JhWQVacCK90jjUixiVqs+1YPO9ZwrbBg6gfyuZLcESA+0UOFKX9aR5yZtXDtlYL
bMQ7lLNt40GBGghCUlyM79N+kprE5bpiVLtdzZJ9NIg0rFjl/sBuMU/soVH9kkMV56JJxvSxYfYp
zC0n4By5AMTCOgsV5zWkmZDQ16iKn1Pn4q8SzqrgTDCW1594cKvogD7ols36Tlf4ODSQRT+BLDX5
ANfTawleefnvDTk7jVdeAzDqLzmUoao14HWfQY4ZVzSFKxCG4Mc31toOazpIOJaERvRW02WyEmeP
G+U4C5uYv5tgrVx18tvEfbUnLb6ghb6kcK4TtB+Z+JnmiwFrG/Fs3IoSmph3HR3uEO3nTzlOQrY3
wzWbwUn5HTd3wtX2056EDp0BgsFSGtO+T+Kw+Vd56VrXLYUNdUVWi1o5RutjrAR4pb18CD4dna5E
RzgzoEO8V/AYGtXk+YSjtty/dAFVtyJFyZIROLzc0vJlu1m6pSdGx26xVmPBwqP4/yjFd2i9t8Wt
yFT+B0dwrJ3ShlXHleKgoTLm09omkjWq6Ox5GgmBHk/Scku2NF4zW0nFatRAP83tD1JrKQcC/lZL
/rH0Lr33PrTABWHJrRZ2uak6b8ZB8RC52BEJ3M/k6pa7nvf4m8kp23KfLYO90WvJn7LWNP++8OMp
uf4g1BLtoxM5b6W5oPazIyV0cyVFVzgARvBk563B9ar8FLpp9VcESxLQnqpRPgRaZggKDgcXuChp
zuCtUCDag+NjA8HjOevqe+jGtAwD5VrtdgHm/vtgiL/JgWUUgxjrS8exNvD5ZhuoEejwlF4x3v7I
XT6Smt/lfLpexW4n1mLO/wj8lIFF9X1UD9HR0dldaHApOKGpM70AWO28IdXG+6mEYZcPDv6iTe74
MIQyZHzX+VhIbDC/21K/EW6hCo1k6D3ZRyoDoI96yR7QvosngAyxHAqI+ntSGP+zpSbqYXm5TGLr
bqEldaYUfBa8MWWZDzOYBDy4Eh26D7kG3DlZMR7finjBuZxhL//cFUHeXYQ4xXjr4+/oeoOBwEVb
a/5i/7mNbiY/FiIwn84tbmujWWKzxjvczu/6xcRl8z084lIgG3VV0kA0tfcn/XgZCbsKD//y40Gj
Q0BEvwZWvNiSBLwZ6P7WzLU9t1jRCLGjGP+qSdHjUwI48hntbcrb39biydiv7rJFaHR8CMBw4cSf
YIHx31NW5/y9pZZcYWuZabnfn4TtN85gr8FBMfdFUUPAOkP8Gez/5MBBHq/Uf7UxaVmR3647xpLc
q2eP9QkWqMJirMX16ihvSFAu+Zvlej84AX5NoN/AMfCNhAlOiiOesNH2Msqyav8ANmJ9zEXfy7J3
w6ysVS5zZ7nVkEs+Ztbz/hYY5nh/m2UFXAv24SbU+FXS9bvGNYHhR1gJUT6mMkiREiFsI4YWJ3+T
b7wysuFmOm0vuVWcIgJVem44a4MRk3o2JLH27B5vjBIxG6h9mDcif+YiyNWZYjl/TGttaY+ASRf8
1YBodV+UIVgz2nK59KK3EQrL2UWZ1sSHWwpWQQLnNF6wO7xFTjTz2Yo7Ij5b3M3xhnxG/cs4VjA0
fZDzrK+YMFaJWY5HHMieXfddvxrXJK4uQi2zJ1ONz6EX7+7uOjcNUYtyV9NNfdB0DksoDe9VLfHc
CYDgKffpjqg53yGj/R7QZmPR4Hi7h5pkryqVxcte4hPD8DKzXX/ftnbEUIZQBNm1E+qt3mFiGnb7
caCN8RjkoenGYaEG4pcydVPRLnME6Lk9Gvj1D1jwxYyBlS9RFfecUChxKq7Ge5xZD8zmZaJnQ0Yu
5saw+NdY5QHvVJrImIFSisznUksVD1j9vNQL9G4MaxKNy6IrndE3cPvn/pe6EV3VF04X5dZxwx5I
SRQnTgqzGeEPyFFnHKWYSHk0iOLziUCq/bVez0Hbl6dKLjFTLkjeuaJlX/gdDgWC/gbdbAgSyfs5
rGnV5nQkr8F3DK4X0tehgT9vMEYe+i1LbdV2mmVsOmZ7D0ry89lT6q6LGpO/cqE96iJOWMiCA2Pb
+XD+ec1g//xM1YHlntkJQa/Ix466yXtUrroj2mBo2aKpwWGKS5gEpJ5n0v10CXozTAPe6sSIvnYQ
GHrz+GQFO8T0nTs6McISZ21fawbImDzrYIQ84V+y7lvobOOpSGlERm1iaBW1wi22VOVkhn4aC0k6
ezz9LmFFi6x7+oBg7SG1DmcNn/VJM/fBXG4cbPdQ2qFrFg+GqgTyiIEPLu+kB1GAcERMyombhhMZ
NJbYEDm1Q1MJT6wNzaMAHiGE7DMlKcOqI51kDtVqM5KLCBpAN9P/jvh/tYu2DefrmtxgGLRS59x4
fYLswJmW9wEglgW9nEmqg9ka+fnEWJv0amEF97A6f40xOARvLvuYSkwxoBz9hMKlNW8mjvINXRdC
vwMtvxdXcW68uu0LElN9esi70NqyMOmTqvSC+4FPN3Lc0PZWKNdtq98zYrCCQj8z4cdN7yRr6FH8
DNvDeZh1rwfAiY77pe2U8xt6RRiNCX25VZx/u3ztcoSHCHWAVuvuLzoeMnnvIUE993v64YBVWjYT
+aAi/NlsNO1k3Uq1DL+xaNP9Ry1wuaJlJ5Px9avV1in3/xrxTZKTCVLvKvdLuyob3C7MpXrahxPG
/rzXxMx8R5K+kwx57ndTr8Dd/jqEcI/9b1/n3e7WGaE/+s9fPg+ZL5aJuyd7Q+iPNL61g7jvVBnm
ZxbFBqUQPyASUt9OFsupxP26reoUmMco5DsH5LcE9u1QRq6P2ItaOghejRLJ2HVgi+wK/knIXN9f
7plKcfBOKa0D69wWLnUtaVNa7IuD3y18PgHS4VZXvItcX3Rg8ySyxsVGPp4VueEQ/6zdAqvyeUtx
ruiyHibgXxqBFdWVKmk4Z7ZdPGDG1utJBnGZNB40rIk+PHvhWPPBD932YFdbidLBRP2v1Vv4r6yX
A/9XFeGIWdgqN0nM+qRw8OTobRGg5o5fLiPXCrquXTw+tcQMUQ9BMSHyHDkLeC8s1jbMkFrYUaPe
+r8BhyBsnr62JLmRphQ/XR4o5Pzt0TMTc7HdiXMxxUSMJZ7E6azD1fR4+Yp0ZVMVKMTx6oeQKHbE
gL1w3lkuqqiGlTStD4T1eQOF1mqK//5c4oB9bPFymVffHN2LRR99ECDHsylP6qMH1W1UD9MJfsHp
FRM4SJAHw1BiE7HM9svqOf2uwKQFE6ux5EAz53OPWurNegpakWwNDCqfGULoPt66U8YMqgb6zMvP
tSaswSHMMck0v1QvCabL9hRNbner9/qZ8XBLAe39ylWtU+2wckAFPe7Zz47Ga3jgBhyNmW1Jw3c3
e8gX7FgolXIvRkYiAHD7jEp/oDn2ynKAMZB03HQ+bg+bh6uCeMkMNFikJHwR3EC91hJzM/dIteSh
BzHK1A3vprJ8yVQnUDvSBTArW3T6wO7X8hXn4A4Ne5JTDfx/2OLcxW6wZ7otPlQQQlUpZYWsOzbr
9vUUVHMNJ5iVUn3eVSQaHOaMT/EsminiHjeMLP0TkK2HQRzU++7sQAIFsKRfb7RpHeFhay/ADi3/
iwxs7mQt/u5lQRE0MwpoBfdX5pPxZGrs6zS3GorUbR9wz96qXwdVnb9DhUfco/GYabrfOWcET3fQ
EIEsk1WvHJBYwf5yG8OKLn10r7GulEYghaQ0l2l8HmBSHzxUo/WXEMgxxQqHvR61rasQ3pGltWny
p00aWmDB/wD+WTZlXpLYYzPrzQbrMoCaqgbk8Tej+nO7zy9q3+/vWFq+wQDQYHakkrOvCV6W51nV
Qc0wzlMy7VxQNy1LyQ/sGNYgOuYfhaOn6yzji/NRGL053oOTYymIrUa89ePMXm17UbGPnDkD/4Ju
o2EyCravfP9LFZNayG3E3xrN0GyOmrWWuiQzC5x9UEv5TsRyVzZWZM7QVQGl4QgVip3Ys5AtFHnG
6AvG5jo2LLmnOVLJmigZln9D/fCzRaIbmiDLqlSSnN5A/J1/jG1V6RX9HY8VldYinhjiisWNWGI8
wivrl1u9ea955+d98TOZjOIyraGqd34H7kltozY6noLozkjw5Nps7CtkTp92eRm4u4PkZk0iwyDm
yNVYbxOu9G2DcAyLJp0/KHjoIy0PSJdCKPllnKIdRs4Vg34QND/HyrGX/1A18CZDs3siQIpS9vYw
1oPWtDcitSWUx/dhIRDTty2WTV2fN7/wPGAPiKCA/v8n0afBqyOYzKoYVkyQXd/qSXfsmDUR/asE
vC6tVEZBoN7qnWF3+O+tGRbAnDTwGEcId922aJIpM0tcRC4GHkpHXt+b4YrGXquASfM9Zqi9UbNM
4pns3rn/mqf5NM9aWmTXPhQXDhFO9z5QCRmWjxECHHUuNg1Wy7058F7iDEeO9RYIIXFm7krVq5V4
HY+NRsD0ibRxVZEaCwpGi5x1PpglZjLBqqEPgWqAXEHTSqIxflHiMo1a/ZvlOZ5TRkkIJJJsEjhL
fODzGSU4fC8Ds8aR9NSK45CEBd2wGQGMxdEAJdQVyOj0nSur7hxpZwK5uynUdBx0WA78Ym7Ulakr
WzRxwdYVkZpG8wy0eCRqVqME8C2Fekup4wIH5T5zFFmjgMac81wp+0nusbOvvhAvZzFe+l+r68pM
V7xz9Br7gNiV5pvDeCpxb+Ze+tYZitm6wxGImcRJhsBX0/gheeMPJI1xP5jI2JQA1d6bu12m6Tdv
omKQLuEnZm2VGlV0ohb0Ih4I0fefMqeMfHLtI2BMjE1gUxu1v0Kb/ssFBEikrU7o9UpM/XxCJH8+
e1qX76o1hvLx9/UA8gUdcqoeU9qlZuQ90IMrmKA7MFtPd0L0mm/t3Fdh60KbZb/5VIAwCxl7wzf4
vgcB9BjOUU8AkMsnJwSqanxjWkDcILrmD1/FzNSxOG5oTC4Ldi2q6GHE+yy8siU6t/pXeeQWyRWH
Ng2eAo9CL4xOCihGg6Q/E4TBCccrzWPiZ3TCK8tz+gnNbBUK3reDsWoXWDoZSvCfbI6s+mJmj910
aYEALENWohdSMcdaWVjnh+h7gw6/Ctabb2erWyLBm/beWNREw8VwHMwrueHrtRUjqn+IY+v1Gxdc
mD9X+piI4q5TMnjtk7xxhjhvN8FlSlsOJLo6lZHMIMw/h79LPpg/TD825v9x93esAJDEXM9ZOB4F
6cGD7s1/6/QhGZrbaO3JyHZzPyWuqLRRyJ58UmnUgHf3r85lpRRjxxydXpXPmQkmRMKTe3vLHEDo
cvZq3ACjH4/IDUN1MOHb+zaVR8yaMVyPeCiC/OA4BCTiz9BgTHPBxlmxFPdJorrtBbld/L9ME5Ca
10/vH7Cqw9ACUhft3gzuQbQg60JpSnMzATwJaELYaCmGSqrWQFqlEyhr4CllC7Zwgw1POju3/Gox
FTWHKg+ExL6mGb1Ceb2P7C2MW4Tz4SUIrvktwV6NQ4Aj+Utzq5IUBGeOJObDVKOfxZHSdIghQ8nM
Vl+kjpOu3nIVZ8AWVoOB6Mewzj9g/JNCAGahp1VMFnvOHN5mbabwXQy3319DzgclMnPK52Ky2WQZ
I5Xnvkdf9SKl26bGcooTIdcBHyJAITO0McCw8qh1aUb1IbZsWvbbnjlQ6sVVfQoj9FgRfOI5N4DY
N4tK25lYi+SVgcsq+ZttVUQhXfpLwkrUnAgOQQ6fewXWnVKlEFlUfXDTPNkgOLB5QaWbUjjdzryi
VuMGdzKGRL5w682HvMQhllfUJP6vbtjSSEn3IPl9TdlAM3epyEOtJa7YoPxN6INKP1VtjgUd6ii+
qZt4BeyZLLXOKLNLtnhPkSirWRAUK8qWEqS43nV3QyP5+cb+TBANO4SOnPZ4M/4hAoceSn9Dj1eg
R3JSt2ycpCMrFjqGJobUkmw07u1WgVfu+1CIPQVB5S8+nTBeW0FuUqhC06cG+7AUj2FWSv8JWRJt
b/LnL8OSNFJhmeUYE3G0uv5oMfMC81xJTqdZRnpTUYkIJCqO+qyiluRIfK1ghUgWZs8NPA+LlYdn
RafRoe1wAsp8ivfQlNG8O6DSJu8z+lpHHwTFa7IH7XVc1Q06NJ6bNHXfRLRmTAqOLmR0S2ciDR+Z
ruCHExi1j8d1qskKvFGcvMf5msdMT2wbqXBwCxyAdJEiDRdZ2F/FgOJRLIw5BCLFh93fKirLIbF1
Odj1F17W+8o8HKo5QnF1Ue7IXpUVHlOxlHqS5/pBoOlXTm2YgociiIBAHpVbbeiY57ywaiZIcdW/
UIlHINmtMOwwB6K/Drc1erGWLCT+eCQ6VArWuCfGuBdiw3n22mbBvYpESiCFoV6WTNv3LbXTp74P
WnrrKlnygE5qSC6Uil4IrQVlJM7hDpEh13XDX0w9jELhKau311+hp1TV9hth9DeA8zwrscgPGNvW
zUXub76fKOUljPSLLhB4zKjb9fjFdn0y/LOyM/vMwjheTh2xRtLfrzBPo+damsAQm95LuhRDfhYO
q3myN8UA13VL0B58EreFjNjLYpEQhdVbcdZuqRcUyVQaVdhKD0lwkxCnAYNv+FzP9Qeh0Opld7vX
snIRmj3xf4urlWSl+8RgkP3dmsPka2oCENaZaC/BWo8ElZBo6BN7H+4c8ml6XXRzCUTDQPsyDQFT
1u5WOc8Umb9YxjtD25NvOIV3llGm0MXYR+s9iGBBXZYUpKX3MdG2yC6Zygky8oKWqA/qPT6urGMN
3+B09YhD7TsLidsUIe1aOQxCFfet/NLR8bt1oFPtxHfeS34wfbPvrrxB4hn1BdgqhD92wsPRyigN
OnX4kr2sn8QSVwHqobgrVq9sX8q0Sv3rQofTW7Xb6p1BybhNIs+ImohtvrubyLyavzNYa3v7A5BQ
a6vfLeItA5kORtYppTbxdvB0tW+fDa6kaavCyXkjmef1WbMrz56uN8c7PO8AJ0l9AlXptYtWNmZf
/Iy+/IUk+ejrJkT5oiDkQs0QXBLGJF9xHeObJxTMQ4YJzRT0jT44uNxDnnvNvgOOaMn+fqC/lCPl
GVCmlfhi080P2yc/IykSzgsyYy8+nljsfTkZzVDrPltt18ovzIoRUk5hagWFsB/PVlkHTJxOuWpv
L4eAVK514gX6m+u1G/30ttbIskRXJd2kGe/CYr8cJYMkyM+EUI9DgaAYSG2Bip8SMyBXswR7yqXM
gbQd7fsO9viI3Y2OyYnDQ3K75TU+ekXyu511yVKoakURanP6z7GqenNwaTANLeGupW5aijiC3J5i
peIjiH3lYfdO6+fmFhm9M6HZTK+r1/BvwPoLszY5TQ7Jf7P6aPTZZ/zKoHlOVBEya3C3k9nyT4Qg
yBLbo3QusNAcdb5ca3jcBOrmzUlvaQoZF3rewgyeJEV2Lm6VC8ls4cFhxXH/XDB4veNeWH9lpCEN
R0TFTqYcKW07GArAaT2SSsdb0RcfJlucYAcp/BSgjN7uR7wyT4dc9yBByxlfiPiFX+RrbjFH2PFp
gh81kLHG0hsshUXOsQi+jmosW7sAL8vFEiFLMIcQERKt+vb5LxGgI9ifyUFuHvxeBxHgHViayf9p
9OgWNKzNtrRHA9XzZvkYSYVdzPugjZu5fWc3wMG8pQhtypZR0RUDm6lnGpNvxlBYI5yEJcLE7XmO
DfamNy4v1g+x9u+8HzhWYWhlbchzxpCUrJgRg2k/mlLCx1WIZCPjPuz+1kSDlnixnNijYb5CvTqE
WAVWJ6GE/Zvr5ZlgbooPhTBQIuHNHIh1m+n7ZoEnyA8AvrExaZOm7bX1IwG/ZKml/SRsvKSB0YjE
gzr/cLpjj9XjDwA72G9mtMSnyfByEKkUZCmIiRe2q1XixELJIej+BIpdbZ677Ej2mLsT4xJDDAbQ
m6adGV5OCfM+9XEQh1HASP6KH+fs/j6jbZgzTmKdwPOrhar6ie6/w1gFZc/CrwjRZM6EecvUvu3m
J2vvrn1lw9E5MYHOfdYdKRaLcgE667wEsvBWYEgjjqBR3kzJZlsmBvVZC9txpKH9YlixJ8QXYwXz
iZqwbJBwmyxLrDlerogcqB89frDetnygbE1e1Ddn/wYve+/rugSmSC6NLFJ/0TtRx6WZoS1oMQJT
VnS/rCxHTDVur/Pqa7mO/M+DoawbpTI5bv2JlCggBDq1Q3jOzwiJ1gklvGfzNGTO7qf8KXp3YQqd
rzevgYCDCTYqg9xVWCPfIBpWZYtVSDPTBNDpIEYm9UBQX+QowDMl6UKo2dhOXNv8N0rNc9HKVYqM
nIth1mwDvYJkz34l/2s3BEy0PJroeP1f77pMQSX1N/fbalinGfVByY0D1lN++ZcY/BFOfXAVKDqV
isV3NPF03Gv7KMaoizsFuy6/SaQvOaqJ1qzH9Isej7JcFmgCAwVqykTPsGFjhBp2lhQPNdY84yVn
DwJIGbsGvq6SfuEF3BF6vTDNXyI93/6TmmhTPfKp+f6Zv3Jyqye1/JqpFwFF8fjC3ZxD0OuHPloJ
JSzXBshkNzUHJXaTra4GlixAFwlcmPMrXuxbqeg6Zb4a4il0AIl/2rWJG+rxfRRVADD15ljDvIGG
4TUFu1zRK2olz0+VySjL0SvE58A7dmz5ej2Zcs3YSjYVRTysdGJY8rWjooC0CVlw6Czi5mwr/iAu
RzI5JysgU/MRYT1apA5wKdWyaZLj4c5qFKwUQQfbR763udzMXinyAwvRTN1X5CCy6XKwZQKizARh
GFv9XcbVeWsWsphaIsx7A+jEnWSli7JYOf8fKcBRMg1Cx6uqbXLYv6bHGNm5w1Zqgq+fulWC508q
NQ4sRXDsQef3nKaLQdDIV6l9Mf9lL+fcrVIZOmokFnmabtEyU7asTo6JwviWWGLVfdiyZjMpWBam
/1P4z1f6CwvGoXBun4c8mi0Td3bdiWr6VnnZ/4ylkiKXs64MoqYCr1xzmRVuotL2hLz2gPHiCMdX
hHnT3ucvwc9L32GXQSJe1wWnVm2GULkfUtb5SVAWKHI9zMPEJdzmuWLXmE3jXR63BFPXB1UCpDg3
qH4Tp5TiQCsxUoQIVWajfT9loy26bV/Q6GXylcfPe2fX0VJ40FJ+dFsKqKqDWZXeVbidMMnf2yrn
0Uet1Yo8N0CWw6sHaSspz9gg73cRuiXi5YT4zVjG2ntj/ciw3RfFu+PUb0LtZWxRaPg94vu6vUUc
5j+BIXlaN3BHG03cpaBjvlXQT5YuS5lULthU82XdGEaqkiAoCLCQBaKwY15usxGOVkBlXMJKyIyZ
ii+a0xGh73WAhWYftNr4NbztkeYQUG1hPkdKG1ApOaWSI1MQm8b6sIrUUt4KXp36xd7a+WlnLTn7
ONYQN1eVhi4ZH8aKQKjuuEiOSzRgpjJli31r0Itqr+LyHiSr1ehDkjjuSKLLuIkLHZsL6hzgJ7JV
cKyHFW5iNvTbXankR2Jqeh2S4FeibuJWxqR5CfA3Cd2g98IV1tksI+pyJ7jhqMKnEgRkUFI8R8Z6
AhvIdles3tt33WSkgMDs/pJ2z8SHs1vcuzbycCIoRKqbXjWEstX8xf0NC7yVJE4pZPaRUOZn3+LC
ib919sLbuh4w1gmwCggCyPDDrwVmCybGeJzlbdVMIRvSv6yoDP5KfT3yJyxE5LKMsXSm1tS2GBrP
0s/ImWG4bidjs1/ydif8oRIGlOQ5mlIUYP64SAYsM9+880v0y93CtooWsGgxwuGeLmiYRKxTi9Ti
CjtianVs9UwizjIiSxcObumOJu2vdKKUIMU2KCkFoQl7PdBfBFWNXknG24wVQYRGMwXPixHSyjmh
nnilD1jxgpUpKGNZz0Q4VZc9wZLCfZNsuCDviFpossquEi1VTogZ5GJIwCDz5m0VG2Mbu+YXAauu
VRS6UXiiuW8GTT0Je0duC5StdIhQuhPivXYOoC+NT8MH5DKuwERSgErrhPR1hCBSAFBuI8/ewB0+
9AvC/b6bI6g9ka14zk4TylFIrC1DbTWONOP6/AQHIVaM8+LfwtgJHGwAmbd6NPlNgcCuXmVcWUAZ
Q5xaOwMiiTNxajZMO+g2IBuV0vJ8081sXUpcV1ZI691lsSKlUq52f/Yyu9kB0qPvCmTRElXtJMp2
McIbyMZO6ku4bDfJ1CD4bcgi0lMgqMTvYDA/t/Cputwh6un3Q1dq2kIycFybpmrlLeaC54OGEk9Q
tb9uC4z3A8+kMjwKz6QiHJbVI4JvxGc6VkvvH9C4rhWGMuUqQqWfVSwQRwDCcFFP4/xbY5Sdx839
JK4Ttu1Nvca5HwoJordtaTfDEbJ0MQwlXteoH3lFmfRYPMZUvgnE02la5rx6zbL/U6sirmOvu6ot
+CEzA4oyZXnu8A2Y2hPiEmpIQdnstGFuLdTjAWIzx0rnMOnKD3KrcREfE5B+BNWI75aPml99Ik5Y
ndHMLNLX/O5YTbOiOgGC6ovvoVEDHyCe+HbvPOMzARI6IPp51u8PHNVbm6XkEOSXS8jYQMWtry+D
SR0QSRPfrcx7/shKzidwUar8giRgouyBb1ZWbNZa+us1Xs3TeqzyInkvRNs9r55BUfhlICMu48tz
IpM/Li8PnCvBHVVXoHkQR/qlrsyOAeJFijKHfjHjGRWgWMQ+OfeL/iMeweoqXlxZKjcHGcAafCgH
0JEK01VOaVzK9uCdXghmThSRJ8lmyWWN1YVbC7kPSKnSLmohEfBkR6mBQ2fhVW0knwx7tdcft4AN
qE7MbVAN0OYS1xAjCNB8pXG9PMHF6I4IC3P0vFQSJG3mj103rQIPanbNqGvUf5/pAPUkDlDfS9Km
u+ZQJsW7OuC4iOmrNTitVL0CTPjIKNTbvHB/towgdebiDQLQR1GMqISs87fPkFBSORi4q9Zbqpp3
aBzFwB32PsKMBOkA8zbfctRfRxyIrHDBVx4xc6QYLh4RpQQXmlkyQuX4hntAaXoMU+W5zEPBiWAz
PWqpk37xePnMlyyeEyXeOzZchw2aYdyuoPqbL5qgn7d9KtTlIojhzVXTSRiELZOS1uinRPHGuTqR
ZWSJ6qDqRkUk5DbvgRxAMbKdhHL5c/2QJPVdSucKhrklchRL5KzctmbJiZ86O9i5RjjXr46/iJd0
SwfM8WC4om8nwJqwyPbtRqg603V/0E69YBMafLkQcqpM+eHzr3muDP4Za4ZgxEGN3YdpaexvuRdi
pXYEudoNBQRW99lI3jnitU6swBje5hVALvg16bsAMzy8yrPcxAibLZ6sLRrB3jjBuv3zPSW77tyX
MBboUIXciXKGDltuFLHrDuKX+gfUDQvaONApOXGo5/dTochccrfXPpghO2898W9OyrK9NbA/E+4H
Khcl/YaVlfFV90IY9eNEZ3LFJ9z57lS/1974zKZHwtAG2q1Ehl9Ffc6hJj8AnpOGmn66rQn5fqyQ
2EFLJEarqGdZMG6XVJYTYax7rbvfONaOnSOpsBh5yktxvMdq7X0ZGo34csxG8xRA8Mzhe0qmkXsz
EjnOp3ZcjKvapvBIOboDaBLTDJQjup/TRCllRbfslOhkF8UpMU3DXsBz+ulKUqqYs/1S37GckxNi
MCESYpATmE8+dBuWEOcl332NuhRRWmDTxLenRP3ulpNbM6PEEWZwaRKgPdmlWXtOrPcWffOGLYSy
exUL17u/aojYpnWnawic+88mvAVcmvVcHGpUpU2buEOvU0/zgyy6IGksUPyyHPRNhIxyhyOxFXzI
31gNXC1RPiV1K+lozfgcagcEm20Ijxb7KcS7pcNR3rjq7YwwU561sEZDnvyWlPGWAJX6nQ+S3J9J
DutRIlkmpuZbWUpKV1SLOpAPmtVrM/UGdvs11qyuS/SmQd/UzfBhalWHquP98xJq6x8+0Tx3bn1f
b0gWa/lW04Rh5cAc+eocMUpaeVots9DRKL6wCaELwoNqLKE3jUGArlrCBWG6TYnX+FHuwWjz76X9
hHq2ZJW3Y7ZY2/0ECAkgNNlBu3rWyaBv8G5lO3uG+SabtKis9QhgZDvO4tjxCIbvH8U/G/obRMXc
ZCaD2+ZrdA/tARO2ij+yvxfEUtjQZ5W2+CZ2gaLcXZXWpWonALSZH+//4vuo+Fb7mxIpVpfY3kTb
9nMIBtEAi4eEfsKBY4HbHhnBDvDGRaPplrt45vjuzpmNZz9+7fVytnJlcA0Jks/P4R9k0YEmA6EV
DXNjePXJGDsT969LhI5oCqvMbQP8wdTLoP8y4gyxiNthBNCpd4sjLsXlDc/50oagJpQ4hbO3EltX
XVHXy+N/sr47fF7En9Mm1w75axagFaNfFDvltbl2Pd4sbN/XbeFhYwvZS60IjDrwsbP4/Zshr+Nb
VeyKM0rIyhGVTeWFvZmDVT3mYhuYvGY07I9HmRgbGxUBGXe+Eza4S1BWaiuRVcuKCtHX00ceqUO3
WeoHAesDNi3jV/ujoKRLrdKSfL8NTtzaOZVwtnvgYQu4ieM/lxrmznVoSHLZ0jD3OIUXSkdx7RZD
G0lu9w/5uiWXObW71Y+pXdPpL3fOaW7Fn/PkGkjz3Mmtnph2WQnvuy8oz/rUGfsdyus58/zpt/tr
Lg7jKNlu5TA2xrZP8VgKgiBHOJm/Jval6jHan5f3SZnXiNCwpRX2iDatHvTS6SNlJQnJpH0+/Im9
M9iAxpSYUKrVN+Guy0XMVgJ0rc55xawkj7U4/qnpalMFJyyHBhoxiVyRSIpzP4d/gKg5tJUzIBiC
yNK8vjkVknzlpLIJ8F/D9cdRfNy+vM4YhFShzFY224UfGz0xuRie+BXABVgms6z9W6lSPmRUxRNo
DX/hIjhvAQGNDf9HhXifdgOe3CtCJBwCsU9m+r337LhvfKS2DztrF6NUOTmzH/5q2raBl3uDxIbL
htZpoz4ai1sag/sER3xfGjv31fhDN1v/yzBzKCFF4NC8jEUkniexFbPyG9YInPr9Cx+upkP5RN/O
ZZlLju3O7KydXrGC9z/QUuP/DNAmsYn/SGYpISYOeaquytiaWokgzfFIlniLhH4pNpdqAV+pCBRq
9vhKNqpPgNSxYGxIeVWwq9+1sLUlRfc1p/BqAklznqS6xuSd/NrM7hEwJhn8hVHxISQXUypFl3rg
x0uhFSCKh9+TSDhBPE+QPzU3fbBwuZtqGGB4xBT7IO8Sraakti8yDvWuO5zQfYOyM1/S89NTAr/h
1ZRve9I5kDHm//p2zZeDHkdKkd/e+YJ4CCLyypXRlrT1jswVdS+rFz8/daJIfooRFnfnwCXzeSt0
2t1KwettFVmHLixWKJpWEDGqNYVzUj68SqtpRIXmyyG4khSXMd2dlZM1vrQvZ2jSGwsBFNbEoscm
A4CdDzZJqnGZUDd3hmRgUrMa+drAfm5J97DCw51SoZehdroinGArHf50gSZmc+kduxZA08MCYI/r
Z25F+HeyFT8eSR9jLdZIvl8n5H3bJ88c7N+0RSVTwRYE83baWLYT0dv47NE1RjSIiLrIQ8LZ6HNY
puVL8+XHzIVzF/bisgKxR/6NHEPPnWd0ChQwTJvIPsvE/z143edkdUQYtqG7zTP5nxwrCJmGw8Ei
194Jxz6GuoqLo+8/39iDCF9xerlC7kTuI2n6kh+8y/tW5XOGZLf/iHkx+nvRR7O1Vq7Jjkj2Kybc
jrIqkqiao1T/wCqNAJk1t3wRFkVF4XyvjhS+4JJ/wCRs/gXidL/2XvEbUVBRCABUA+CigQcyJKj1
Y63yedeRF6T8iMDBcDw3VGpqnw5MHy0fyoUf5m9Zx2t9Sa8Pes4ycn3EOoJS6XIYGcK7EZhcHIun
zr1BrpmQkIEDN77jtT6N8BEJMoHfHGh9C903y2b5r9td6Mm3INk2tu931ZUr4iMD97VJHJ1vu2YH
obAV+YXiqeTy3nYjXEj/WhFs2ZtfytS4gzvbhYVWnvhvQhFr9/TXj7sFxmiEU36QB8LpJ3Xtr78U
RlpQTEfT2P+0SmAYx9ubZsGQ9IM3Ga4iw76p3H5PV2QMHm+i6/3vwmLd8y1d3pSB32/7IivwRT0U
DRak6o3WkA9HM2BuywAuIqwD4003gAWVDBqD0JQt2PSmsCtAcxLt2KQxftL1eacnrIBK6AOe0fi7
HdUJ34JcnG3JjSJm1hpW7r0Oxz4GqiqetR6MEdzYbBprkXZcA6GHPE71O53wPDHRGp5kzHqT+T7N
9jrigQN20u+qyN9BNnLGCfML3cgRYm6Bb/yfpaEEhCC9vu9uW2xcMezW6ivUqMwO4nScdwOkXqBN
c0rP+ukknKK99kOPd6BZzxGtE0AQGtjrTRneWhsCFCwepQ6asNEGA1fWlD73zaeBCG6g0T93XxR5
toBgHBjp//N7rK7nSPSzUPC/LHBLSq0nE54FVec2oubAEZSWSKWtowy/zwCNZlrHAp45wZepfO2q
4oWth60HNqbdKJGSM0yf5jpGAppEEGLZZRIdZL4EESmtp7G158+oN5PMHMN8BuBg71qvwmOdWBGL
17Cb1y5OwdgBSl4efzUskTir0sRWZP4s7l7zMYLmsZpBe6xVNgzr84ffuN868gTxPJvTW1RpUjnV
0CFwD8i9t7wGcMf8UGA9vTkOEVwrUaX4oMuv7A07vk665F5NjNevmH0G4i4N800wc1yuqwBaqTe4
QTKd5QyDYjKcW7j1wL5jdzdWubTi9S7KuENPgf0HCx6KQiuehsN7p1xPBr3hMFP5079DmjuI5brF
dTOtjhDSA/pLP8TvSBAjKnokFEU8IMQ0azQUdzPNoy7MRmyUwS9XMCQiuZr4Ql6p3HclzNiqveZh
nfGN9gwEyyTcljYbLM3DS+/Kn2iEwqYs0U4CKolQ0xVaB2Ej3vtK6xwxsEMMOicmiBY8s5OIRtWZ
VAT1QGUdvbwwu6go5KGgMQzshKr+n50Lyb6NGH98Hen4EzPX/E4DlJRwj203kgl4mx4G2PSAMB5Y
TUnXm5FWYU4/X/0GF0XgFkB0zTCuc2VerSWKAkz7ZX85K3VPpXlAksiGDGY3JcvoRKprzD6n7oqq
hSmVlIegTgVlKdlG+yCf+ChaPeTEns8KXlayqRimaNZktGYEZvXTbk65D+teKbYPgqAtCocLLjav
ReAFA8vvcWfz3TBPbm8w/8YS+fGa/scp5xe4JIVVNsXLD1mjcwcqHwe/oij5mu1uA39ow3aSoKGv
GFtToL9bnKyS62pf8TZEGBPNzuo9pYczCJdLKDl81CXq/oSWKJlfm5TuXbRqkJlI/oVzmXrIoHOJ
SDWSeyC2Y5otOcq6/NAvy4K4TiDyV5jKK+cnYD0GDIkHR4ODz+CD8ki9RnqsZUv3cyp3fTwLrQFa
0d5ADRu+iYGKLqMUdFIvz9gWwnlt4z6rCrqVy9aZwh421IiMFj0CKABuwq6pMNUbJetlELcCHoWD
O08CVzlMXJXLjEW56K5vygzPf/XzXfST36PrAZfWcLyhKhedNOvQ6dyWKU1WWVogyHMnFSQvLFIC
+Ywmr6NeKmwfoTFMKXHP0HAP4gqzGtJ/yHqZVtDTjAaHnyRKEUVCU7t61dzMJyBJ27WkMIIlyon/
Z33KYNeFwBt93mfRSg9PGb1C8eXsQAJ1ZEu37cxk40XnrbM905hRhv5/VRErwdR9P8IRu6YSPbRH
ONraVdYZ2tGuGGcl6XRxg56pNfhox6UvXlBmllVi/g43ZDEOEPoNaB+yOo7NGHZzU/kbKujiX4zp
XKDbcukmOak3emoKtNA/wWmQibN7mtY9nwxoXI+IODMIInV40aKBH/AvFSsDE5wX+sSqkeekTQX3
Q7mypQqUkSg8hHveYO9Yr4dw5X0Tc74ivyM3LLV25igPVN7U/1dOPFpnnDGD13wTSF7JVUI/695a
+SbQAeeh85Qmx+wNCrJvrjfIrI2v4kCdhy0TTV+Jvt9WmudldaAz2rR/0n78W4/1mVUdB5CpQ7KX
cvPrxPnwA/FiTkQ+yvNJbX+ZJqg5KpJ71pOfyw91Eh04us+6YuNmQZQaaEGX4X6yTWgCpt9M7pjh
rXzYOHzDwLITrBPs4IYSK3MbZh0VGZTxIdg6f+mjSQnrLMAr8I4PFvTdutng9BMZf0QABTqHlFnk
XHR6Cn1Xxk/lllvCwA0NcixIf7RL2ge77J5mXl6jQ3RzxmxaoMXw5AyvcIDtg0Io40g6DH/Y0LkU
CfDauXtFFZMoCLG0HacYMWEiHKtpueZd5jj85tkDDWzsSSSZEqZHWTFTdJ6fZt2PMs0q3yJ3lwSb
Gs/YCWhc8RXbFQdEvYjQLjEPe7nvwwbxGH9UkxQki/DGtUCk4s8y7RrcTjJVswnQtWRi/BNzj/Zm
gZ9kZ72yBsVIFdSHxY2EsQnBRLR2BoYKnKgGabzrDfX4uECwK2MeqEw2NEK402nGp+3h+S/IWSN1
CV3e3c5o8to2FZQIFkrwZNJKO+i7BrOJhOHJvUHGMVMEbez4heoIY15j9G0oLjR45UOiJGnOgqPF
Yo/poJ7ASTOMYEMMl815Wh0RFbKkBOyzd9V2cdGzbXI39kIMUFFoPVTBnpCCm6A1gO9Sr7xBLaZj
iGTa+U+TTEDOsD2b1mZua7/K8wZpgIrQDBEwkz0OFUI5KNDh0vns5LWXcC6npJqXiKKAwKdQeUox
mIVm2ZgvRhDTbzUZUW/Kg6hOTssk4ge8jR4fYDAxz67NwBSYM5nx7QzekLg+dnV8jYYRPNC/FPsq
cnM+pX/nfV1cmO0uexoYdFjFHTbLT38vuCQh2QurCItMqasE/LfnDN2+keRskCZyQEC58Xq/JBpE
XJSLvTD7ipfIPyfxgMSVxaHtebqXvimx5jNQWlvJXOCvEzdDMh9fLHfrq49mP4O7wQJHsHk77WmP
L3ch7hNeKo50rfIx4KOFnWJYsDFPCmEXaOiHsUk1NnzlM9YNmBgL+ryFzFGMGWE0iH1joW0Kn8Vv
vF3GsVHHbuFB4P0jZYnq9qevkO8V9ViTkT/720UZdP6MjDMwt695i+bvFNh6Sbp979qtU6zY4rMY
xYnvnmjPrCoDNIYgV5M6ZHI94tlh9EJoyAtiKKGRwa28OtIZ5g0WKf2J4X4HzKLffvasSMmn9RfF
jE7Jkc1N/jd4sz/UPSqeP3BCXG/jyNEtt+wpv+JnPXfts35CyRpYk+sxEFUjpRz4uARwG1NSObIq
gUnyRHCHCErJucfJrVjjpXCqmGLoQZw2OJiZEd79V83slSSvmpkSGoT3/EPvddT0RwlAHqhmrbx6
o7I01KJC3J51J40Rn/kygdwcjPdxginyNahbpx0xLm+CREnwknCFYsGT6YFILJMpAo/X8l2MItBx
ArfS6OL8CcB+7cfIK2MqjJsw0g0flqiW4jII1I0lEx00Q1IXtOOtWo3/JFhEcHGeTqJ9N0nHPdnu
OqxvftsLyfZhkx6Q9uVTvPOwjnAPKOu1ue/B0fXFSqAhzdkUxtPKHDc4h1w9yXKTvgeJvESOc9Sm
DkqOgcQW50OZEJxKEX4RR5JFLYxVYy3wMIEgfA3Whm32DBaY+V6W9INt6fwBJpl8aeKaCRF2yy08
f7uyALBPgtzPRf3iSWrvTAA/BugD52ee6tjF7G6iq3mzlMoK5CBf+Tum0ZZHujqfRrZqBLsiJv8w
wzqOM6fSk3V3HjRxUYMZMZ2RQR56r8SK46exfKViZ2cMxCcCovV1Y5Uo+3L1pscF3j+AuQkpWlZI
v/HnhrCEdYbHTDTqs3TEZZQOWoCBxwa7URqkj9+NZxm7LT2suLgfcYXo4ctsAkjUVNxTsQGElgqD
KJrwqfXHnpIdcUTkhzzDscl5nUhKq6Zo0732jeVNJaWWkheYIHvYFsREU+iaZ/Ul3DwLXec3f9/x
rxGwnCO4PcdegGqZhMMIVt+i5eCcxY+iIyC0JGc/mqhThlpb3UDLgQhN5Dr88pRFG3rRguNq9iVc
TPJf4Hznj9sgTE6dVDNtCXgF2Och0gWrR5Jg8EwGXq9Y884Z0WIpWWZ/kFOTUxsCxwqibpoY5tWy
nTcG8MZyOF03axOuD/xPVbzdeT/0TDnJjgqUkRV/wIeDRi0UJAAD9N05JpxHU6XGrdPbBt3JvI58
GjnE+SYVl0zMu6lLo6eJKksskioXz/II7IKZfvsJJ18KYSTtwO1uxqQTs5qOWbe0WunX7fGxCmWQ
7uvx09oHZR16q9Scqn7efm++bi5CuTmrwuDvlQgjHMlA4tsgg/h+DZmRL2q5cOmKIfGKtobzloEz
q6v60UqKJrTz54sNZnBw2EGn7ZeLRGykix/FaJM0pTyMIQbkIrYgdj5V3KDLGCnFOzIAaLlaOERf
meG3P/Sq4wIpUxkpKr4idzkRnko4eVdsiT7TiKSNHjo1cXu/25CJ+2J5MO6WxrsJkLeXV5bbQSbm
s6GYGaiVeSlBOYIpyuNgY5Pc9wTCzvWi0KRZhJQM+w/Wf0WC8YnfxHfiedcuwRZzjkME1d6Meqlg
fBNz1bsKd0A8hD2FGcAIoQvIOqEREV/CbTKtywUQuTzZz7JQN8uTyXaICd4K5pupvcsafIADfeOd
uOVOjo5BRB+vytdrAt/7T7n6wqY2XsUREUBSCUCF5a/XFAsahw9qDlGo8a9S4XZjzvBySLWZ7y9I
Nl/ZThmqkcP/GW/8bbWDa6qifQXyYxTdJ9GwfqrSI8JSK8kQLL+sGdGD3MDdtsOzG1i3Y382fCBf
mWOpt/sKt5in8/oGbEpHxkWwtTjmtnlKwZZusfM4E+KXg1/BVO67Z+c/iDFF+5+411KA6VSCQq/E
fAh5GMiVLzYIQmbblYSgdjaZXWkWaHLHQZtL+rk7vVbqHCLvSFG1QDKYrfvcpqwnfVmsmihfgbW0
zsFthLLd+Wl3IL/0AVyNprl7l5Q7hgOB/f+/RyM8UAcavG0dOI86dXFpJKGTjUhPaXeBamEkn/5K
yh4hHoOOKXptJVeLaQHI5CMUD/8fVmnj60JYKc10iaRvWI4MKERjVsDwJhZ4wBDWfxsEr3R94hyM
5UQHAI7gcByMQ3oKJUx3kNoXVEMJfzsLHtLDbHIS63d8DJzWHuJyBJUM/T9qz89V66iWFv2/A5pi
2skM6zZC/rrv/QTFaGSGKfd9RZrVBWr64XALDqlQvhFpWEwKqltpgkMbrwG8rfD+zcGqTXoqLVkQ
2UbhDOX9lObmPU/ePvESwEaUyHhBg/hJ+b6R+APmyUOz/fZNBMUJJ1qxkYN1V3Z5/JyYHn+rfqLB
pNLoulCkB3tnzQyVvu7DTTw3FMXE0z2ay46Hix3zqgb/jeOJYIJn8+WjwqphaghhRux3Ye6TPHyI
+Tpg88OfUlvPhkqjpumeBQboJyRVT4usOf2Exw7qL7T+BzcD280Ybn1eL7AHAeMbg8YXkGHfOYIN
JzADPrZ60cskMwYtbndfp/AhPzl/pv4OYyFjQQprwLZG3eN+Cyr638jT7iVXYhfa3Z0KWQ/sM98Q
MkIqUtjUVJAB87vEPSd0Tqpng9F7mxU9sTr0u0C7uAIhT4ODXIJpcdAUqlld51Bo0mJd/bqpQhhQ
4KDrZPyQJvzA9DFzHcDb0g7FI/IVQ0OEqpBiAUfT75SxoDRftHtHoJQ9yGZiOg4/IgYCaqTvnzmz
kHOPqpgU+7ZozSaUdqOsO9orRjc7GpXswHtG5f8VESZW2hB45lQOg10qz4mOJjQ+jMJUkdcMzSDr
/19xPuaUaeqUAVp0Bu4175k38Zspwi3D6AnhJDDWJtxTmRul0mUj1yLk2ExE1ZpiE3GHN64OI6h3
Yfu78nF8pIV3YY/xCE+QrjZZv/fw8VfnMxFMy5MqEuoSfqpvNYU7PyaPo80IpLUyH/+j+EreVerT
yuTGVgtHWvTR2bs/t6wfCR+JO3SroPpMIekH/ZvSwucLd5dnLYAjrOB8xoO1eELByeG7qHhIYSLn
c/7Uq5sRnwQ3j0U/g5JSPxwU7j/ymqFTNg1XfG794UHTS+CA7EY5XO5VHkWtcA2wNs85E22RtXhr
3z2P3TXTd9Q9pNIpV0HEBINN7s+0JAFED5KcfroenkydoUNd8IUIrJ/uz87pHRe3+85bZpl/gOY8
4/84RfY0W388eK4htqmwGfW33WLMQVSc/s2Eyo1PR0hMOd3+1AB2Yb1UlN/NYwyujWD3yCzoXJ9y
4mFw7xNOT6sCpBJAIWKD/RpnbMvZcYCx0xq8KP+krqTyfknPN//d7QhSRiRk8RjqQehxbj0tuLAs
4ra5PoN5cnvQ5CGozDY5XvpMCzG6zwzVjHpUOFdu5Wg7jeNdETeZcYVFHRhEyF8GVqE1tQr3Akna
PPl1S4KilWMM1iHrgTgdCiD8A5yZy1khSFMGrb3u/4E9nZ+MboxfGX69ScjBYETMhqnMeT0gQ+ov
3ywqVfeZAKa2C3/inuOot9ZPzX8rRCSqMR5Y3RFQUiPieawzVrkFUk2s5EMs8TRY/at73kwhohF4
dPE5W+3O+AgnGiGrEbopU5kCNFFtyOD/38AdgiCgPdhXEyTcudIsxDt3ldeF4VOSO6RxCDU3O2G2
4tfP39aSpID6NcTpF06dWKwUcp8wi8FVG6bYQGTzSqBSwjszfag9pJ7UrphqfN1+kHus0/rGWm+O
+DKy3SlqNAErO4Z7gnvGL7rXxM6AvQkwJoC0cducL9jxyFGMlTp2KbjKNm0VtF67L4DOZ9XSYpR8
B3JCCXTBHqF8cyjr/czh7BLkLPtGpvnWi9AvQxbhui6ZpMhmyej5YMT3VDjBTv0hNaGDsJW2IeGS
m0SnT+CRO026HYb/QYhR8877G+BO/YrzPp01o0FSLHxGKEj4P0DchBe4Bd+ffz/aH+4CKvE/3Q1+
51yD15LTGe/JXq7mQRGYCCkmuigfc77PfJ16YrMOPH9yytWJxMZhRS5M7uQhBfjX/O9nJiK0cuJZ
dgZ6jBcRLppVnVFQCVktqMIvHAwed9gq9NEMRTv/1XmmIEMb5TBmzGBZlErAFPSehqgjKTOkRz/8
0gan5BUgtKe9DGoVsskawYlrhnS0TYikCpmoM7Yt0TTLXe+7geFQ5L/E3+SyOW9qeNLEYHxW/hff
UPgEmGsvTDMVZt3cafxNP2HURbQkuhAvA0C+FBqw64tgnrZ5S/0pEYQST1O82CeZDVyqBpHob4HN
+ZJZzlzYZESUUWz0l+WOKmQ+wBc55REzPzTuKWOr1oalnMyc0n5Nl5yvqIawWuElT3kL/pCfzKkx
ddt8HwUZ+7NL9uSCnIAdr+S0xJXShbM7zSuFDsJ4kj6hn/LgfQAZti6Z+nKXdDzCPLzCil72bDT/
KiA69dOxcly6dlvEd5OCzXvLpMPhCRkv8lF7lbgXYR4cBpcgqyylN9MEiVu4+Ci+JTIUv8hDfdtA
jIw11sYO26UI53eZl/B4NDarEY3rMydQdxhO+nz4TLt4JVekWj4uf1aggYEMNNMMVrV+PG+ORSa2
3mI1IeLKifqcKPebkgGcThKVBywbY7NBOXFbNCKcB43IFwm77h9hflCY+FAlG91x8BEia4Txt7Ya
vG4zL8Mw9T//X9Nbvr9HP2rnAbK82x/iECnbDNDoJ8WSABZXcGtH+z4M37zgQdc2pxXlPiPse0wz
9B13k42oClx5IUEamBxSAKxARNWrs87g/xvZpzlrD7fyVtCFWhM2sE37pL/rTeEWrQSsunLyPyN/
2V9S2xXDD0ePpmXKenb+Ra5Dp7LzhSfPVl39cuMIskvcdSrBK8fA1muzk+4MuAmI4AswY5Jl6GQU
7ZYKGaQlfv6aTHnHk8bJrlJuqb6yPTZ5KgNwbOI98rwIo/TOf775mLcBSw5oV2lQ/KTieUzKhcRQ
9snW7OvDrdSdXWSVXuWOVaxq9QX4w/WkbdzFB0GILoPld7Fki5pUytjdLtcOijX22YSjQcoNBU3n
EThFA70WIOo+k038YLMue4OpXHP5kxgTBns0QU6MTFjBaLSnjcbZUaZ/ac6nTSYVD5SRmBB0KUfK
o63s69anfq5Q76ah3ObHcsK8Kq2bnPdGz9dhpkzljBfBTpTL/AHpuPj1s0VjLwuNf/g029kVKCjK
msU0IaD1OHqgRc8/NQwJXiUgHlwqw2B4rVre4pzvlePz7NPfPyy4g0I1QdDmxnE3kjg4jjV0fXDw
aIAvVAucsH0+aczC8bYJ23c5i41Wmk3qEYq4okDSS+WW/VbYcS9tNG5dIftDtNW5VIyOPbuuTqm9
M++sgMmeuRjlkRM/oMtxYd15HNHW3llZpVgKrt31N7JFXv9qTt5FSGvP/eqUVIrCREL23GgeuZOy
eRQHZa/O1xCrU+A4/roWpt/TNiLAAVWLJN6role85WUTriqwM8azqkGs5rj0i/RuNEYK9ATCMIsV
MOzrnC2yWDS9kj9mLA2QVvc+YFF/k2+FpcrzkJYUdBQXKesFE3XGbYkMmrvLBFg9KNDIh7cCbuf3
HbaqpBH7Sa0UbYk3oD2v09hPWoyCnBmw1naozk9xBIDg49bgosCI4Xcw8jtOwKthAFJOFYGU9gEV
X2o0PZ+qq+c4dRx3azdUGixMHg4tdEq8vldo8fzdof/DAPanvRxppAWNFsFZOMmi/NMcXlsiahJQ
jGkskEPc4DakOFViROfwF7MSsXiYhG7zGX7zG4pV/sfJFhjXqcf9xiJLBsC/q4D+V2OcLpySixv8
zJVguVhszAx6BT4oJg2HgOsVez4v4pXFn5XFl10pBQ1gxCwqog9xNxsebSBZ3nzRRj30u+qvTOHw
9O26XdM7zmHK14c+uFJaUC475YWis1fsSTGo+gEdCl+R6+XAvqVFj8hHUYc0VG8vLa4orjSyroBx
PrFLoku0NY6oVscJgKD57Va3J/MRSh+kzqFVcLniW5Ws9vqEnNhCM8iPyFjvs2C4562vRkJafACy
w89IM9lRT4HSeINzIKQlIdyicuQ4EeRGBnB55F2gz4yO5WSHZQuAAze1i9SCsKhT0KMBGlMcue0r
ZhSkGFD/cgu7XSa2M7INzMZr92Icv1BBzVK+xFOICqWDv+p+vubjJjEGypcpvXyRLtKffg2oiI9H
jF1oXtshmdKzn6QHMrJUsgsYZDUMoZ4x1pGLJ9g0zq43AERuFzUza5zEpWyWAMKYlpiCfpcW5GiU
wD5jIoeZKA/bT87ROC8VKNLqeq8wp2k5BRQoLN49g4Qr2ickx5mfnnCzyukaOrnuIFI8ZaosKCfh
aRhJPiEzE/Q/kRCk6ulA+qg4CiNVDuzKmxq6IgAlapr/sepyMIkTAtUG76ND0ytRmc/EBXMav9M7
QZQjuUk7yQbrQUgp9A8gOV60uoLiAcISTl92gjkATuepDn7J+TH2lnDlT8YUWqz7M7XnOI3QJQ5h
dd2fYFW2xsMwi0t5frtdQWNfGfA+S/eAQzLPL1aSLGiNLEsDWskTJIBvUXsnkTk8s6XDVhJBd8Pj
ZqCRGQQQGDGA1RRTvdIf1H12USj7x5RB0jYgZHc3sAwSoE+KOwDFvzCTPkcO5p5YOhUbszhVIkzl
mUPfiGPOB9m60ElR5dgs8ei0PyRMqa+YKUUHRLnJVj3kimOCQwWMrwgNW7gCGI0kJ4LCAz/j2xOk
9g5IUzNK4lc8CdB/3ejd4CmqmQkP4BgYvFqzxy+vzvSx0YG1YGfeK2o9FVdG9bWAsIJpV8t6ysxG
LBsxIsoJuc0naUOHQeWfXtXumKX+nlHvifGXUGsghkPE7LpD6QZsvjgag8+N/ATaXLxhH35bP3yP
Zc3lhFxmm8g6rgEajFbP1PMSWR3nhJo0gDncBAy6dDAX9k/u2IO1lyWUL7zeb/b2U75LojuOVI+j
/hNppr8UI5hDipRCXkAQK1Jq+n5+HDwOc+SSY0fCspchfSL+LuweGyAJ8hDiJm6PU4GsUXsL9e0e
z6cKGgPxep7B4WQWkRnUYHRQZRB5IABnhWauxfG3ks5nbofzh8W11LTEVF32p+zHzgHNBvyouyvV
XA6wQxrG52yjOtkJ1ReUl6lU+eSHenDp/MjUonwzJg50z++4soVYVeNoLzK+rXJGx+M6rpToGadY
cH6C3x8Vq+p7g/0Nt0+vY1xSkAQOcXEK3VrSouz+2lQislI6/21agho4Y1PjjgODH3iH2OR8r0wH
rE2rlqDXLKAKP2qc53mvwfpMPYEyOyvOZddvwOtzqaS6Quv40813dIg8GUVStjIJH+JH43EcGq98
qPCL7LcgCLYN0VqenvP7+0/tphdWEOz8ylKBrofkXLUWIYVUy9PlL2XrMYTeu7KweleWwrVfE8zX
FEmO0rjN/H7s5rhMNnZ5i8nTrOf5DofmPz5+Q4dXd7+t4/KWl8btqZ+9Hygt3wpJVrQDfSHmHnPR
ooC0cctGn79B03Y8TDFHD0yxh5sRZAXTFcQV8/dJxEDJvWhlmMnktFzVTo1Uy2xCU8wClJ+BVwRY
gcp4Ah43DNhFpWc9IF9vj2SZ9lgre+tnhozi7wvKj5+eEeGwHmDUtFHqzCQ6ldd1dH5E4UNLdhAH
byjvZy5sOeG2Q8AXIGAYt3XNEHnuAcVsz1dDqjmqal8moMXHU1RH5HGEZ0l6fzzXkIMdlZC9KbWO
YpfPA+ArB+3TgDSWU2hNHgc1sjA/9GdC9GkpEvZlD3WhCEDDekRWd442X1gaPirUMetMhTjS4NTl
CXRziebZiBHzcoTmPl4ZIB55Njvn2VgvNhGiosOehnxR+P2MQxAgur545b/5FB4rKB0XkSmQFRG6
IqQ9m9+x+oF1w42ZhXWRofv0PQfdRu6Bz/FAvKkgjJAqOCM6O67c1L7Oo9kqe0F+8if51RjZDWb4
6A1f//XGHNOsEeCrQ982EFZ22+6XcHFY1E5Kp1Fy/oUvrA8fiIXqXFvwV4uoZqEKzMaFPS4VTdwk
1waK8Bps57akWQt6WkoLuAqyNToRAWaq4/dgWEeYwzb1wFHMUA00Gt6VVYBavCJgz33zfLRYn0fv
RK+XRpsWflUVtBY9jL/I8fSa8asDAsVSRu+LsfVHBz7E2vejBSbS49p72Lyt9q9HHLdjxP6PDUZg
Hskn/qdd/ZWXW3ye1bDm2Zs/RMtQQyWOjBPs6RsBt7JlEseshwf/q/+IT95DcC4H6XIiBy6yy2EO
PWTC+BKC8434qX9Cu2ufoGfGr0We6lHcVGgQnHzpMZ7mE8qP5vTED81k3L1NyDgRZVJHfj3caqUC
PTSU44ZyiZdITSzMUSEzZW63N/tph//UeXL0094wZcCkLlk4KwhdnY/Beh+ZLfnWRXd7tExX8Yd0
gcgw/Di3wvQgJZjT9N21O99KFkCLgW1X6NT0lEXkJLgvB1oN2H7FOVlzWmBWLOQMYp1BZk2tcBEV
HGeRtf+Ack0zVCrZwKwP3jbVMkDdZSyUI4hzg/rUMf3Ce+gTj6175YBED7ZL1MltJ/XniMdHUMyH
BPX3t09swwF6c7l3v2E07HOsauZlUn72WF6vElic/jg+pEJK5Q/ZXCZjyh5bSixv+kvWI6a7tr74
cJUZUbZ1plFN6d6zlrhvrknV16vkSMt7ZPzn7hgT+knBFbXIiDJNNUEeSQMYi5iQFjZM15+rxWoc
DIqm1gpHp7ecPhDCyGy2/+jKJwLCLyKMAzm50pQIp7kIa5EFS+7NjZNYzoH9xtNoGKquubiadVsJ
DgxdGt1A4GPYxliPiMM4AdfYkWrMNuV4K5c23M2Izo/pP39hCJC0QPQu3NqLH1tJCp0JzQpfb72/
fSulYyp9DBosPtrFSgOq3cNHcYhJy0VmsIs4aZC6lESC8j236iJ9PViWeAimQSrgwa9W/UrdgszI
iNZYs41nMSaESaPA/vfd/c2oDn7F5ZMCMTTdnao3bGNK9l45fYk8qcgjxxyaria6AGZLX2QXUI2M
OXpPU+N0xN/jXiG5g8XD8orIKaVp8dSpy+Qk+eORwgtLvyg4/fFmiO8U/nEKIVEM1qPkIsbA/1CV
0+abqv7RYe0yJ0h94hAeceeAh0fOSA0j1YnKk9ot5eGLuEU2Hsr125D2RfEi8HVwkVZ2A7s+kRHo
ahIbQr3uC6Y/7MeMd4+l2ICwbQp8aZPm44ZIxsYencd6Uc5SX2QBFX+lplr2LyJYyaA5AQBtD245
AkF5qNN03CnWDAexQRdlll3XfA8V6MBD6QF6wB6XB82ysI3IHkIVV+kX5Ce93nqkjm0ctuXB257b
CjWwS1aLKCgGqn/yMV/eHBWGiGHUDBjI+rBNOXDsuDh7HuXulWaRGvxCKG2BO1W1O3oNZXg+2oNR
hP8OWBnWAgYUA19HCGLgYYHvyhMuSO13cPhA0QM76TgZQIobHHjb4fcrXvoehq3NN0pwqbYttAfT
sf9CPn1704t6q6/CWpzP8Ho5WWAgz+Mw0ih2GcBoVF6ojbECX4ba0XnsUVAyMAdsqaQwfTD5bkCI
2bR2bQuUlndFOHVs2WOPhTdvpGmzENqRcVy6vlC42bmt/kQHUI4+gee+uiYsqVI9XxAc5aatQ8PW
WM8uebBsa5KMJzuzT6XzT/suuELnY7NYndcY2RHyiSe3VBhnxVL8B+Bbua0BFv0k0nPRqwWrq8nJ
WrXnT3R2lj2XOStJIGvpdp0rsamqCiG/MT2WwQVdLCejTk0TrhkSIpy8hyvN3yjtrQxNfDfoqyNt
6bTZo4tAVDGMCwX+zByrJEz6Bh+5AcQiGWb+tpMaWKB/8kbbAEPFceligkKTllLrxbWbmzz+c76f
5auU65DCF+tprGDdCcv2fdJwk9j0igkAl8OpLEYbyUM4UECmOalALqKv/FJ0xloQ36sOub7QulKI
vviQsSK1WsBx8hpMz+kWa25KGseMvSVG657BIrrS5iVNHGzti5djm6w2+v82xM9AcYR+q1qYU2tS
4y9jksoI64JbLIW00YS6udmTDAr2AAtVB7uqj0PxoyIE+QA75r3igtb+iZs4zyJkoEI7aLI+RuHh
WM3jhjtJ6lOozkfqL+7DfkL5CudsfjGzHJL4PYpmpFtm7ePRsRS5XFLLUgmN54wd2V+dF/9hK1yC
6r0KLahpjvOShNi2PixaY52L8BeWLXFccxFMKNBLX6IU5/I1y/g6LNYFi8GJH2bqYuov4S5kPZ/r
I0rMJO+KBmMRtaaRVi4XxDaR1uCBhPQAs0yyCBwcgH0VqlJPxNpIsM9UhIiSri2QECwsWC/uq3XO
CRI1Ce3E9e53uvgEL7hJXRinA9NNSzt2TLAiLOVoK6QPhHWrnvJnp6BL4HZidXdck3uoTBqo2Mxe
DATdipCiAhoYUgHZtqQ+Kstlv1TNTLDFVmo+zFbjKl369P7BEMRz6I4FBsw8Fd5zjbgOp2fayRFO
s7kcoyX50jVCQX3D99PnramIqsCZeIfbWZR5CUy190fNbIthO1y/oE3SArQ/vMMpXPVd3yyLLHAz
WLbi3Uo7/9Twmq+gqd0arJboMq+IkZZr+7LcZ7sc+wX8v7yNOcMhV9bPKSqt7PRqI0mpI47Rzeca
1PO9jc9RM4aqMaWu9O4T+DcFvXacmfvIGgsGtz74Aep2K8SlXoqqm4I6XXPLj8zYusjUQ+9VQRLN
ojHDTN6DpJvm8D+AzqItQxG+ox3d+TGQHdv97NvsRpAtlSHLHAmoN6RvnRo9A6yfT2bR16KKFcK5
DK3rBWzwTkaWw9PO7vMYifLTQGVBjAqdgv3afRN+KGsLNzMG5iP/DsdIcyUsZRBFuxIicfYFcMeS
dCfxll/4E8B05NyXOZoBFC4NJ6/43mbKqxWxUF1N7PNhJ5UNpjuy+bsJwS434qFml/wrg2hsDw2j
IiLEtIVgkSPZ9swZhJBC97lZiya1L9RtuoL2H9db0IHrZmV45uAd2HxRzObh2t75wyyukVC1dAzc
lQu2tthIeqnEhdZr6LYtfVCIOP0f3EnVlyiLcRdq3FZgoxw1JkGasIJ0ZGWrQv4k5L1HcrBip6n+
WKe9CxfBw1CC06s8O8sBVjTo2wo0RdAgsmnfWPkuwYal2Vd8HVZBdIJS2dCMdMvLo3HYkyjPSlpn
QIB61NUIkRUisT97OKLvm1ao6MZyHm9x9azXfissxCSNaionB+w883NynMfcSEou+tDk+p9GGIjL
ihEUr4N6FApX7keGq4nbHnqvTJ1jVCQiAGi/8FPRLJQf9IlF4qwfZ8vhtTe0rkx21565rxV92CKb
Ykl6XZZ3LuKqzZmZSV6KPjzmDKc1lAdnMBXYERb7/w9WMTyx+C5LE6b4ZXz1lmdBka4dPBWG4TpZ
PuZ4fvth+7bFUiDiFL5Duh2QBK47LX2Az5BCwHrm8t2syF/BDA3uNhKQulH3Z9lHqXfrglSqsFRT
S0K80bAhDtIj9J0GRwjJr4C4HLHefPmGtPLYxhAKfovYHV6k6T5HR6WjUfr5phthRDI7bB02gzD4
xbxL/XTJrGcvqcychE1KQCA2oE+Ir8OAhhROC9jANRTlW+SB62nbmEP42TSdV6s2hd8lXjbPJPo2
QqqPmdJYl9dZXRqYqUeD3xMhE7g4CcA6im8tLvE/1BbpHk+DX+gbyRWzr6OX/mbyfkAgj8F9jOpR
Uu9DMrMwwXZPk0ynkoSJlocNIwkhQCAa+n3NPMsuDDJRD77mSMOByqXxHhX5uG8NC0fpTO4ai2zz
RsXAY5rdvkTjCoKYtgihxX6CuJ4H3tfmZKj7EUMLKeYxLyUxlmxHBX2JUNhKmIJum/qXxzmJHjlF
a/1FtjLAOVBp6lJFNPi9Jo3g2W/cIXWjzg9iDBlVOBYQUVUEjNgBpDGsPp+Px1br4ofgYHFfqU2M
VAPTuOgMYdRtaRg09UDb7pVenVW9aCysfn/vRWkIX4xw9G05BV++pUzAhigygP88Higile1zALPs
neSA0PufYxfyG4PZ2ppv9yEw8oh4ckLT0Uir7OK7KJqj3VMP0ZrgTL2wrfojSSopvZHFxbwwutSt
WSAZFRgh1+RvxfNRsIHzeGx68J6uflPmUJ8XRSPxLdCyJ+e4kYox7EVwTcaqJkyaZGls20xjZ9M1
gRtqO0jEvoNv3dCEytwDC5vQkujNa+8Q7wddO5k+tMSscpYVKPaSLsbOfCOQOmBv7ms9ZPn2f1+u
fkPFv8IqjY8NireS7uP32GjuW0aF/HP0h4WAg2+reTawU8N88F7/fbPVbooDqR/l+W3OD6crpebG
4+DlCbt9Yy9yPMHR0JlMXr3RaGgMrDl1+Kb6Fbal31DCVCoZQEYPTAktlhn/3WVgK3fuCOIlO2hN
XM6QREsJ8sdrVUKYtR/Wsmb3sKJebIOJnDF2KQC4VK6KYtOvtGcyfD/vjILUkrUPBTmNocwMrQCu
LIEcEAyYjALD96GKwK6NCeWwJhzYoMOtPtY+WSTxTWyOfL/F/pz94XBuAuxdIZBy4dIPgJSDpWh1
WqHGdud4V7itGmIM7Kbick7fdWgYQT6+aBHSNr37VFAkopvzycKSs7lcj5T9tqxKbd+oVTLaX45k
LBBMQ5HBXGPCNH2ll4ix/j82LKlbuZf7eCwyhT9oOLuivugi3rsE0xlks1byZHZJTxd6pVM1ttmB
3C9RLcc5QHFMQEumsal5hu8NxT+mTmgB3XQbmP6GQILJ7D8ctxvXSAhXEm7AV9RkXFkJuyYxaq3+
+HvVHkDcx2Z0KythZ4QewCBN6kFW9arQMFT8v8pvhwiJkns97407HAi598o+OsUYZ0AfMH4dqgI2
Czdj/mHp0S+YpRTVj9ZDGg4N+uOjtkPJEYPobLEtOTnR9aMejYGRDuHBjg7WkDqbakhcgNvPm+u0
7mxrVpUyWfBPLtmIoY/9cwXi6yJmXFIyEibCWbhSu8ERi4nv075rt3WjfIBgL+Vsk3RCMDHbqEi5
5rz3lCmcAKQUV47p/GaRoSVKG5WlkV5bIzU329IHTQzkM625rau+pj+oRk1P7/v3Zju6/FOeOIxU
z888CB4VF5ZP0L5x9gimbNd03Q8LXZvDPsbCUW0JBUM++OWsuR6kHhG5VcXQha/deoYac864Y+e4
Lbi08yQ8ZK7Y5NERbtM/OBz5xqJOBEhCAyHF7UYzG5VeGTYUFmzpGBXFrbK+A/8KCCaFzYfkGv+u
aQMPjTErnmIE3dym87GtjkjI1x0xxLjbQZER+f5mDpTGqqUvjFy4JQqbemaR77v3clf9NjW1B7QY
yIlkU5SUozoBUp7MrXBZlZPdwEO8fJn91OGkbpguV6doscMkKVH7ZaBcqiZAPJBMltGj/sqVAjdu
1yO19r2g4wLTYlsvxVfBgmJAIHTEHkgdValPNLDK+kO0+wI0Z25ZXIEk63ZHrutCiOPRvpV43bMG
iOEkXEX6MBnyoKWMtDGhc4gTZDy7AK8kpgSOKWhJdLZ8RnTDlL+JigG2WB+AKglXBc1vwYcUluFC
rOltOrZiuLQ+Vk1lIG9z9X7Uw/HdzfzCcinMkCgqgUfKap6lOUYD7fA5CVL9mDfLmkO13BX2Halw
k2YfECXR88YuJb0+Luu9dZqako69ENhhxteBdLwvD65hhx9ES6u8Z8b7gjm1BmoJq7VgVdT6HRnM
V6uU0NiAfKO+fXqEvPLmhMa4bYUKoh1Z0xa19nnldWkCsW37A+ttc+OFF+pXAcQPEpHaXsztt506
etl+aXC6Zh77AhV+JCHPCo1S2R8XCylMxbQhL8exst9QdS4fHbe+1T73c+uYUGUMV8YiyVWuqsj6
mcdnTxkxG41C7Ed0o85Vaz1OtH/grlXsMnEdMD2pkJfmAf4At3TNIR5DyhpJe8b83XTczV5WT6nO
BIBrM8uui18hmejsTOtsZQMHvtYtuu4jeST2n64v8l1uqAE58NJmorVzHmaShC9xXLONAlZAgt9d
RZQdXBqcOlXHO1vB+88XiNuVMb3K7Dh4EY/0Qg2YidHI+BEjds4PMYBZbajZDo4UG6SOVMrbWFuo
e7FLIgqsiVIYYEinJYFZhZLw44tonOUREGcUemvV1GWouoTX9iT06lufXeoJjG2BKD2Zuzh5/qLR
ddvp4R4NzNJ6lap4Loi9TQJMV04YZkTxQk9yxU8LmgIvn46eWKvGHgn0qqSqPFJzGhO1BR2t5p7P
GWye2TsCMZtrpsD//GY+C6Xucgj+gQdc85fQBuxcri2gEulGO1sh3j+aTgjGnm1rUiUZKlVs9hKc
hUUoqpj0ETuNvhcruySBqSf8r27YN1CrZQqFVnPLPKRg2OqIxAG8iAbSbdvVx0HSr/NW3+IPjpdH
wPX2DZl45cGeGid09lBdif+vW9Rb9ZF0GQABOSAg7ae9+8W8+GRkp6BPrIOLjVmOMM9PuET3vLyW
DP6st0dbG9KzEDHh3nOaVb65BC0GXnmeeptcRJ146YokeXeu6wdaPFxn7z00NWEn2bdrasPtE9U3
JqidTHw7Ds8Eu8VLiJBU5gAQhboUQA4wCMHL5xm1ogXqvnL8N2/6+jDSzUMzPk7DgRYgSMeO5V4R
ue99iIWr82FoFr8warH1MTVpadDKG1wt366YzD6Xx8yOxMiUxJneTJbSayviT9Cy7hupwHb+z7db
3ShVDA8eK7rj6poouhNuCS7IGd0iRA6iL7E7PFeellagmq5ZELeWpkVmdn57xU/l5+mS0br0wYLG
TcsEwXNKD2DCs0UV5vLx9V6/Qkt/n/f+goWxBAKkrm4Q/6ibayWb+Z86nlSN0Ci2xUDz3f7r0Kji
Jbv7ENGfrQ2J/L8lKEV9CG8JlMJvIrxbz3nMgW2Ihzh9quc01MBXJJgUrfDQGNQE21sUU8upyBce
AJDXZnPTxyS7lHei9BNHJq91PNcm+o/oRknPHfHQULG9LdRUodjwJl+BiaSsu5/u6D0Cj9hftfLm
MuNF9BvUSzGdfi31KeyzQXHgqbVSM1ANgYUGNczVQIIj1DfMnrwXZEHa/6g/Yhna0qDUyoK7/xgJ
1reKTuoDT9UKNYJ2/jdC/07YgdwwAI1zadQtDa2+qRh05ImX2dsuSMu2pa9ghKHV1qfbCrP7BtdJ
coMiAdl4Num91XMwSzZGohZDMFkXUvSDa0VMWRwMjeL3VUK1dkA6W34fKqzvsZQTpciuoLo1kYZX
9wMB4AyY+oYSVCZ93SGRbnsWRNsUNLfMi4mX7ukhFap0VcAXCgORIBDFh/n1+yfcaCtRVY1aSvcS
v4nzcZSwF6Guuagj3ykQmsxZaI9ZL6MzHXSul7niVBNHQL1HEvrmAjO6zpWW2QX2Y7uVL2hxK6yP
Gy/p3Ag8NeLk7s0hxuTKt224W2inT/Y6YY7ihQLwhH6mP9qOYv57TZuSIKUbdiE2OVhCiwlCiHNV
Ayd+5CsvPUmsLHe38m1lnmsLQcdRFlDw6fK15usl2Ia2LTavrZPCe5uJ+Tgg9PfqG+2JR6lhVdY8
tJXYorusZ+BCMr5L2xux42+5AS3osB/nTNr43r5f41AUnzjCC3NwUiWUIqof3R/IMK8uJnNKpSSk
YlQELIitJntWFfrOydLXsWCl/LobRJUoBMe8Y+fg60MUxYvs6f2HzlkmNxZSGGDaj4XFrTTnW1ZK
kWYGJz2J33q7p/0LXMapjz+trQNjJjCzjJ+OsQocXMo1pR4NgKUQN+oW34BJl2ymyJmyQc+ocBu7
F3MsENB+yx0NF0AdFL0ySh705B7uUS4QY7gr9BGyXEk3s5tWCWlWqgipIWKNzPobb0iKyXWCCdoN
V2eaLfdLjluUxJWE8nLZPJjK4vgrXgygfyckkKtwJ8vSMRUTO8Ic+hCovjlGchOGEj5PSGqo4ZE+
FSUE8HvbBKOeNqpLEbx0HwI4bVeuT+iWcWWMuYutO/MSRY61RrCk6Oyeb5Oiuo5HELuCYi9KPlop
GWM3PiJDFzeuJXJvCOuq5hWceQGM3lpBE9bN6PSRe0MHaPmbLh08NVLWSQaaGKupHm7UT6+nbrJz
p2ccaxo5wYBX42rTxAM75VuMw2XDsx4dvnMyUnbVVBaanNk7rnNJSMLF2UyZUSI2Nbb67Iuz/2u3
t4o6Uym8t747cecwB10YA5jcaHKqY3JsTw1HGm++W+JTaMFerWRLCp0wvCHDjXKlCTf+6h0sXRom
iDEl1caKvp/RTO2Bw/pSavxRRYHiTyuoUOS0EdoSCrGeYJjC5TofTBvX9cckdjyGWB1XatHo7S31
YbuxTWAsdLCjLLcaLYHEjZwHSdVy7gwobCH+amidb+cKsIV30xIuEbyXrkf/c+6U6rJtcv3gCbkZ
/B3x87Qiwjx2WWyE3yyDW/cBKwljBup6pVRqshYApemGZoeuhqslMz7+ywqsLpjOiAqu+Db5JhW/
NRl1qOEodr4bQgupDWUTVMdIHsYUqIRlXGfNYY18Pd0YnjuqXztfNdQqe8m/OtwGbwdjKBepZ56C
DrRKynLTQ/Kf4iZX4B1aS8CHV040+XhCIGiwwpgmW3fk2MGIchbcu2/bHC/1NGXm5t627bgWzHot
9upBLbQuUN2bS1AcdbKsEU7O8GoPCXl1OyFeEAMQj/lXEq1GFRM10Wx1uPi/J39lYGxxRDU7Kjkp
h3ObWUIXtl27GyAF3u9ZplRX6kZPjKpeKS2YUR0RRF/Q4UX9EiwONyQhjD+qshTa4lPy3si8Q7N6
AAKmvR/VbHu0mEuXEWq7RGh9X+pIBBB8lu3GQ/cnvzZkGbOo2jQ+nL33oi0pj11aDKu4hDQmfEop
nbz36sBZiKKueAsNscF85zHgI/E98TfLigDMzOC+MMTEd1H2gwk7yu4ro7b6IDRt/SCsCjfPX5rz
x348r7sqNn3XBd7RuQIPrepl8fpPirc5I9D9KNtUpoShmtzQ2/Ob2TVtXrX5QkJJaPUV4hKOps6A
5NB9PGWhl8UGRbi/rMq3ICipYFWvYR6EVTMPj4imsZMn3zS4sLPErz2+eDMB/3PfnYgy9FuQLU0u
6962lc4u+Gx/xO/+dXsXN1NvTz/xtof2vTx/I7ue5HudPpfwHokYwO5E73GolL5aaRYR+NafYCY2
zQlZYdEuoZolSOchQD22iuiHnsOPgL/zvNOKq6G5jkZm2kufG2sVrmKher5eK3LHcGl/H+BiH/Lg
/Zlcb7jEOwYdJUjOCpRiBnEVnikqLuGJtMuF4BSTE0yOUeeZNGrrCtWTld/0q9qMjwwz7pbruahx
5bdo7iabnkjXou2Csmdjyv6UkXQV1zhI5RxcKn6H+lUJz4On7J57O/B9HtLUQB3DK3iBX4Jxi8Su
WgzsSnaZFjFYJpaXXeg5WJBuHiyngW2H20Dl3fEUox2wFsqpSD/xjgUPMWGnq/2wGEeEeqWXtHb+
hz1q9112BaNIFMnsi56Wl5J8hk8kMrOABsYf3AFhP0CjFSEMTjm62QVM3WODH65u9L+hphc4aZR2
NjO8auLo3GbDXSNyz7rg5IOejqGwBvKt47xsjFIvmg9rnB+QiYSzb0gax3IDxvYaNP90IMMrkgUp
zfW/Lt93q3t8/a1RGuKuEKHhD+P/i7Zvs+1NNKd6PCdp4B5u40WenYjMp18ekvtoNC1FcFzmauzB
2WEHj2GKQxv3k6h43hu5+Qk+iKeZwVAHjG6Zgw80k0675UZ25VzaBkcAECgzaiS7dgsDahoPGaWY
Mw6yZvmRAJk+NX5e23eoClmfu0A7QHLsvCSoOxBA202M+ndYnekIE5YpuF/c5m1ivCZ9kFZDF5DI
6uJN5Qto93h2N76SVuVkRElKoJYdjHmGRIlIZYUu6DeqFOBkJBPGYiV7bC7r4dMoSIMmIoErBf6b
C5oN1xpUdn6hTG+e6xkIh5/pY6c4Nwxg/6Goe48KdYXuqXXifFyRiMTDfgCET7IK8fA7NsyRtgSt
920URHsJYah8LhlX0tL85C0v5ozZOG9P7lUHRSO6V29LqD/iqrr9fxxxH0tHiT1OM+VPlb093cZj
kb5CPlt/Q8RB1Li9GtlH3qu486VqeypAAj8goVWfjWTFCfIGQy5G42M64EC5ylBWzIi4XptnsclJ
j0fbkfGyVhnfsB3b8oht7O0AlqqIMXYpO7rskf0lrql4tJK/8t9AKoKMD3NQT1jS9MQXmqUOe6IC
+UB2n/RRCOCBQic6xjrfeMrX26248F93D8AKXzNlM121z5H51KoSmdHQZ4Wvj6SgVwqLxEbIHqiO
6j/IUXYpRUSWgvzuVs9hRihnPu9SEwQDqLoLSayA2xeEval8Tfe3Npm+sXkVLFe3/vcZvuANemPJ
okRROb/0gCRQd7E/2wDxVVyL9+GheU44qt6lWBPAIlF7yw6scLxrkMTs99O4Cng3v8Y2ns8mRmPU
eFXG3vOLVhhLqxzE0kDdV5m2mWiioqtstIYtnnlD+3YAaXWKtuP5dS9g7vklBkWpq8ZD7HbhNYc5
f1tTU7aVZopTxa30Cv8i/TrOGJhsjDrQErcdKE0I/hmqjGSwprXZVyfhOTfYCGjXcxXAc2EU40qA
gxU60MX/y8opLb3TsVkES1frU9G0zQnTX6fkHjpFKKDHGj9so7trQAOBaqLRK+KzlMd8YHho/CcI
zvJMabpqzinuCB4/AqXMQ/7pe2hrqOtSwlQ9xcWz0YiJ7zhWTVEP0FvbrudnpBUGFGyjc6wMDBsD
wbnrcyofptee3hCwUUF4cHaEWOb0vOAmJZLmTzTVMTlpRlvztk19NpcI9uvuxlMr7RkZYEzyW/eI
8D+fXqYPqxUgMpVd0xIRZCDI4bK8RinGspUODmr0cvvsCZ63E4RpgLU9aGCgfXvMp71uoj2iP0lq
5f7TuDPdAPqK3xwdrCYpIFTx39c3dhb52beuZhxAJFpz9eaUSMCgFTxx+7Rg3U23F8aHk3SAmi+1
5suzwqNA/lT9JTapyFIfo6KBAbmJ61oFtLUZCNsRYGiaKdtTHW0zxSUhSOyyCQWZGpI/QS0PMENN
3+pdKxW0G7/OTt3ILurBIqjvykQFpGLdBixf/pdGjqoBZzN0FwPcMYNkZ54wieL1hkgCMi+eV747
A25yrqto0ehRiVvhBcjiqBYKnoH43bHIqbKt9cJyIWYaQBUA3N54osxWz85Mldbnkjfv64vpjkZe
wF+CPZvcUjhi4+vN11286y0HcxzU+joRXJW36CaUcZQdF4Dyr5VwJcJANcKT/Tiqd0VvXvBUn9at
62/qlxLfXir42c8O5v7RJ65rHSM63uW53LkShk5CjS68/Ar1hDw4qpqb/wJKBBnqfkIEQYVjrHJy
u0K32VFTLhyRkRU1dUHeAU6lISFfkppjL7yMF9rL/DpmHMkh7KfTorqbJ1o7UkVT5k1ffNc28iyR
ICNGorBKWUUZATRGqA2JmG5bLqBpPMa/4WzQ5arj+8eXfIqRzTvB2VXWArz4/r2FwiY3RxPrhZIj
IICBE+4iMOwHm+8Eju1xruLMtjCeLGI2nMoNf2GlvdHvpuTCB1Q0LzUZB7PfvQbzOWgFpxWNv9YN
vRmOQBEx/Eh4hlXwqQ0BwYATSFyhZIZ3quiNA/bPlujt91HGGnXE3oalpC08kaEam/gfWDtzkFyx
LaPAPiEp4QA1PXx3EHBPgEClZVwLZ2//kjESzNyMrKqksrSQNqWgFFWmPg8zUq9GQVDTWM93MpCe
tKbCcdvH8Q2RXg64SDkD9tK1JOjFidYJhBvzsF7ChRkQ8fvdfJi6/kZMi7kvacKmOPnEv+ZvUtsa
urVOUg0vU7nPLOTMHlTdeB0bmMNAZlMYENFgVcwVvtud2djqdStekYYMABpleanbwXZJfomVPVR7
tzMI+WQq3NcXYB7a+f2CqehxvolmD5mTjepMuKlL9nmL6V5Tnjh7iqgKvYnIAwOUBjMPwCublHXy
CmgsnkNSMxlSIZGQWM/41eGtbxfDtURqKb0RGOecmng31lrXY4btx7zN9Z/Hsh6Ytl5GPlWl7Fxu
HZOZ5iG/CLeWiY1HPQ67HB3TWCXfvyWZpOhLxbfMJA03uofnkfE+PLBxnRHRfjuwP82Dsy9Qptmd
vH6M72/+xA6bQTJnvnunDzBDtxnlB360jjR0xR5T1EXfYvMTNYIWJBtgQAR0FAI55F1M223PoDvW
3P2JFba4CejGtIvxuRX5+SWPz4AYtxM8+BTB3odjMsE6RlQYmlRgYIw85ferbsHmJ9ABFSdvPyXy
ZBFj6Bs1r0007ewZijCDVCu7zaOFFYIiVTTe4O3e6gYiV82gXhvmxgKbF4gmLSsiwb6z81eGcRPN
PYhwki0twFTqFiVBf3W49gjaWvDBXj+Enoa068eMIz4m0OTZ9B3yvC8tWSbiXxyTHIe2IGeDiajx
yP3WQHvcItyu0Ga3v/KFTDz/1KzYiTJSbrZloM8msNjHUjBG6kZ4+1XqxfnDtUubE9CnWMIA0P9b
kTFh89qSbKAxoLp95Fi/cJXK+hkf90lyOJv+dKsDEFAXYYGgbG1+iSNPuEAPTts6+H7x2ssWbZMh
gYHZkPP3N0RG3jjd/RKVBpgsU686ad3yEysO6MkZWsdeZA6Svj/lwr8uPmV2D17AAix86mL4HzrY
ZVREz615WIVL/EegHlZJr1rtTepXr/1XcH7z4UAahxHd8FKdszlIRMq/OLR/wSXhpV9XBunlInmT
c5H9J8vrps9ok3xKSngcSlelOhbrO58FFNXYHiKHIb3E0KSahmvSMw2pxywS2+ETAFDJMHVD3TDm
OuQuhYVfFjCGTtnYaeoPeg2conx6HSHQhxK1riJ0hmmplsmxwLllI6Am0nfAXpa2o+rdr2EEbvGc
8Ypyxrk6Tmiq6r9amLuopOUtcawLNUg5lvfiYc1ec92RvDsHuVkyWVYEu0uShYvtyOKJGUAkyOgp
8C1ZlIDG+fiDRmIK3r79sBRZifSuCb8O0klRYkdL3Vb6Jbkui39PIavEwQpSJg8Y+wvpI2SGIaZ0
iiyyWdJEi5ICVU9C1xfTcQ1dHqzGpelpRlI194R2KUOigIhqB1XH9b7C+oPxv8XF2GuqFPY/RV/f
rxG5q/a8x08lvf4bLvfsWrvqOB/+ZXb6EFh1R7cVVQ0ddFYD9RynU0wKRo/7fzo06onnROym+N8a
dJV2nZsXmCY3EsnxXM1EyucZqylsgWeAmJFcYXYAkeMmV2/uYasucPhcQbre+gpSg9Tf43M7xCsP
TFMXSLsMSo65iWgPZ94mozN+XihejltIh4+Ao/UiLEIRgoipQULi9C0pELkOQUd3U1cUcZNWnAUe
6EDdmYKML29s2efEoESVX+7y0v+z0zdJo9zy0Oqb5UelDnqPSVZ6T9R2D6xNm76QJA1QczDJu0Lg
fHQKQ89VWAoXQ0X4UfbCTN6ahbP4AQJ7zmMhe/4Eulm1j3KsAJEzkyobb46iQSxwCAkAfWGdKuR8
H9dBRYyGgH/ngLD0eneQafvbWmB0kv04d1JPGsDOpaCsJ7EB/YtTN5HAbnZqceQByxMUY1kb2xAL
IeSSMrnnAMB5UiCkJ0YnFQSZ/6/uoY3QQ/r8uqmeCD9xWPA//Y2riRNPIczrr14cTtySxdgDbEW1
Lzwluaa7Sy6quP2LIgm3PtKsnb3/t7xAFjdu777fmLRFWOtuPL4/PL+c9ICiQh1ltxI29biJpbrX
cnnoygl9JParvecujZ0vFFy+AQiaKEl+NTCh49zWTtxPPcZTNS6SjNY0DmnuTM/w1q+r4OWD/mKH
WOa//R8VdTvcx/AmQYfym2Z7Uou983/29hQZdVcMPkTnTeCSYkc2dyht2T4AkxsbGu1y5SadCLJr
OUOgGADxRkH44s88mggVIl0GB1Na5KQAGGQbuTxrhfzezzelTJ8iuwsyaTVv3cV+lYpH62Splj9G
sbeLdEQ7XeDqagIuA+d63fTwTobd6TZ9VzYn4S762u0kJX155uuFJtaMR8YM23dM7pMJOKR+E9hB
AA7CHtS4BzD0m6GP8Cqq0mvDGzr1Sm/AP3iz1KxKVTINOwXOPa1jFFB57OsuJWVs/o+O40r+J+M9
AJ7fux9AzPdOsq5A/R4BlsKZHSLTojTSMhyROwRmJp93bTv8ZlKPqnnBaUjlxyEffGf1Xo963Ay7
sxk+nzKqpGMq7DQ/6oINYZDiIwQC+qzC4gMXtNtIVcVatERvHmxYjP8a1iBEd+O5PO7H8k0Godri
+CqCQEPutACzuRCJsIMEpW53/y9nKmArED55kzLBp5Pesh5Wa/NEmLAOwuEzObuxQrH+cRXqjvow
ljEga4pi9QbYcp/bnPsQ9QJet985NfQfgNUt/WS3PWGr9S2qBb+G8X5EfmatpKrVvEA7L9LvXTZn
8sNc7JIgzVxpGJJjz8/2hxmEIKfEfAPXUpkKxb28Nb8v2w5+rdcsnu4sjq5n8alREkzjwQ5OOxGe
TlN23elWjo1reXGxqMUhNu84kECTCRO0FaZVUdWu4akumVhnPKMsgAB6nwj6dMUxKxR7rGyHndJV
O+FiOexoPaIerqHqepCRH/CVg0Z1eupa6oi4OkFO1bzYFV9IKOJShE6UpAE94rfEMdf7H1T2wvIO
plClsiBUx2qFsK7jh0ETJ4htQl6ZtdSHSW5wkDvozFkkWDrOnbSdttpYH1ygJztKMU3LZzoM0U2+
xWOpla/yVlvHJa7yCZw1Zw9584gu6BGEVs6OXXrDvxuaq8CAyU4umH9tNBlMJOtxBsYx1CYYo3AB
CQTOIkmZLxT6OnKrk9FdALvTRT2K96JzprtmB6A0xU+3kB3ngDCyPyMxGX9gjIs/UYuFrBGReWfS
PyLLwf52m7fG8e5BvSfkErIBvtYDhbLoQKgQCU8YzxbXqC4MtAPOsP4jyzwhH0Q1Y4X6CFAu6zpR
BTT2G/dU7iEjaUahjB5rlgtPW9ayeMyEzS3s55t3+B3qCdPiUgax/Z4Z+4Fw+LEWKhyHjN5gt3xN
aFrdrLnrSSvvFkGs0k4LdUxU9GBsKnzEz7w02OIb9IfbD9bMQBBNLRFXC8BWh6F1T2wl4s2v/gYy
cMQJJLcHZEiEWvH4sOusGTkB1Cnqf7mlrd1X4QYqszmtxJZVRuQYXa4NoncxoqBjWdmz1v5HroNl
aGgAH5uTpP59NhcGS6tvOl5sX309tOKyMydTVuXDexYVigzewdNDAmEO3vFiJls9oBi5M0Gf+7Fw
m8HFeGYUgNqCckwrTchciEDfXCV7yIUf8qkMUNtF7yfGLfIqu1oedD35HOL7nVPQ/G7tQlwo78XH
Xc+ePmp6MSeiOfqM7OiNPJj2wy2DNsbnKHEUxrrYtj/me8k1s9Z4IhPGy/BKsk/HBmh0Ep8+1+R+
dddE5yq8OMqy3DOZHkKYOG5uJYGjMt85Xq14gVTM2e60+a0B3hx9XfRIikFXF8xZ79xQKOCKF2/z
aJ3yYVU6y8n4ITIbiHIRT9XF1WAKQcp7HJWresB+vAceZYnxUUKO6ahrd3uzZ4vLrKVrWxHzMiR1
Vy7Rw0X1duSAejll1sd8KmHI95BiHAqSeDtvV6/r/umgwwrjyq5z3Ut20L0uA00KBawimzqh+Hq3
ML2uM0ko31nTHdgZJnYYwrf0E9mSOmwOLxrR0ULtioAAE7p8RlaK4Al5IfwzG57tBjEEwVPuBwmA
p5lbW5VWfuCOJNlAjdbUinq0eTzt83iCndS4s8EyLEzQn/uEm0N8zoGQUXwtpMzG0p4O5rEirrgE
4LjzAyQBP7yAMx+66fIWS05RfFrnbO8+Ctu3BEG2TRd46T1AeGNfLBTeSgNV+v34vjm3LFTQXMQS
DQej1uoIW1ybc/6zlFrwPvQxeqsQyGULSey6sMu/QuBxIAowIl1FXejNm8ipWTTqdsgepikhkYjz
JuX93KMkM6YLYjuT7K3QGVeSkEgk/tWYZXzd4QhoLLqFfFg3G3gBBl19VMA6wapREpuLFYeH/EMJ
93hggY6iQTMI4jAeNQOl6T9IEhZMWoRyrlXAA9UfoEc0Q2aCHvmpBJuHlhEnKtcwHEL4jliaS6ep
rTer+uXEt9MVvtSx1RJI1FR9F6TDI5h8JBX8RHiennZ9Z6vdEVEsN5GiCfQTeRpMPvh/zdRreAcK
32Sn+GJ1SiuL+9YObz+MYYO35vgWJazM6H5D687RkMMeSnfbZVV3Xm7zK6XKZ6qeXMnfSmu1/nbT
4DbuJJNytakPjdqvl15Nsb+T1LIIuGIWiqdT6P6PKxPVtYH9PmoOILu1N/I7AQePq9+wWYQgqZOI
Oap/T2/MofME8U3DcJmUku32fdSr0YIaObUIgELju1DMVvu6rLNauI8bnOw7Ks7thlbSR89ZErwL
SdLvptL4/xxNSjm7NvtGL26waxriMLvWGX3VYPeqg5P7yccJIsT3wcqlWn+kc0UXkS8yyTN/Eojo
qd+y93ze2j/DCWPGJjPstKj/F54AC3qW+Gq+BnPZdtW4jhLTYVnwwM95/Wz+B4aMjn1EFIIagWwY
1vOFgKbXdm18AWl+vLxqO77kKUznuVQ0hPdcbHQUwhYrMPSVvADfPKgbesjkk1Mw3ywLj/j/gJ08
41ml2ZBXtpvMZZGcN4vl/aILZbYZgmKiOTdYhcCyjcH3HmQkOp7AQj29DrLGSo+eMbl/VaWTyvCs
gXdJROqVz92PhrNuLZ12wX/FJ4NxZon6gD760dWRLd1JpGZX1fs1vGBG8ThGtCA4bVPxRa3m+NQ5
fO+LtT4daxObYEbnw+QALWZFdNp5gVQdGC2j5l0IaZPMn+MpKbUiOKF5ZTVoyU/Y8xOzelfpNu7h
/lR9KfJxYp9gFEpbkxT0QWizA6PwR84YFbS4IS/GLi93vNd/b5ICvCtYygVn7rhfj7mRqeirJA1I
637u1qJw8qCUG3AL9fdmE0a8cLClAavONQNLxMYNtFqnikfANazDNWKUIHWkIOtEDRwm8RWseMIJ
CP2js4LxC81lTW78D6h920PtS/J2agj1gwIWEErN6mKuHCiY98QNdaupoHh/vbzCH+8Lz0Sju7Sm
CHPbfTD+RQhpefxDSK2rniEtprJUrijAXDRr2Hsu6g/DlQ4aAd4bubO+9jMlXfwlaFlpi7d69Yj2
nQuJdPicC6rzF5NWQqDQYd0QhvO11+/KAgNEDO2/AVMATDM4mDSM3jsqClfglcJdmTSFS++uwNCO
nXM06+ZvdQFx52vYZY9ajmKWcGe73qVmJ44d/vjYBdfyqVwTBvrOdp8AsWZlPi2JJkSkcABH2thf
OjkFzZzAd2S04HetUNuRO5yrC5jiFXDxkbra7IuqUliDKoWLvFOCLBX0+AMphqLB22tUESu1JT0j
zCFB7NxOL7vjZaGV/hFej/fk2c1iWIbhv33mxO26VGS/jRSsYPZCL9Ns+OhB9eTQsHjbwTx8U40x
ke+VUjrsZvxDC05b+zAenQQPWiI+4cTOgwQU5K7P6db6Sav4Wk2CrtTlgqdDMJDWys798PHAH8Wp
2+bFiA5d6BPPz8JBky5cUqfIMSwazb8ydjZ8m+2GBITHmhxEd3qZBYkDAGztzrigWAnckZOjw6s6
E5bXLREVyT/c5GvUQZmYlAoTuSy9dZxKqZj8O4cS+I7HnPnzv+n8ODS6bhuXL8JepU6yGrQRdI8A
iTnuO2pYBJ9eu2oPWJ+wFFYoiAa9Z4SgDMtG1OBB4vrZ3cmMdPxglHAtiwziow0bK7nI7/7TS4gC
ugayL8JooJ4VrJDCxqXcjiN598AdpEb/Sc7a01vqd1rqZP9nHnXLfprEj/XXyKJAPMhlEuVRnkR/
HJydG48Ih4oosnrnxaTRaGGXU3jURNipByGrA0b/xcQIPcjUgFGPYEEol2sPzSpClQ8LZAoP9WB5
MIBnsFkxbss/PqvjclwdyMTANl9QtpcnevnKtkCknwXMKlrC6YVhto3nn7KWHkLbCys0mIFbxtja
z6q1pHGG6fFFPEbitHN5cfhkEYCkUzcMU3bA/KegqkvA2YMMUKvLfDoWYX8l/VbaEZXrSQUU27MM
Qm/FHjyXxnpHNjEJhPPPYPxUvgGDH/m6H+2H7YJFKyp2nQVPiEAbwK2HAu4YKcrDGFkhngewqMaF
oIi8cL+X8hj84GPvY8Twl6bQRyaj20vNP+2Lvlhly8vAcPMJA2C/OIwrVzd+vcoXaPcU/zzAVTjH
VwMREyzhoIpCSMQm4hZv4vPeVGtYxvxCud7yaX8CHGhfYikPFffYN1Nzee06v2OcNjOZKRDAmfrE
Y2Kl5TYk2XG3/87N/wHT3aQN6VL4CIKt2ZlN8w0O+HvLXozgEsurBvkIYSfRY1yuyRs9yLAZjdo7
By7RE4TE3+N8TbGldHYxMx/SzLGm4Abb179y2zSRdQ5jVdtZNGwLylTmK1rTv92MCiW8Uo2RpTw7
sgeALjmi4LE6A6vajqnReT00/YkE8pk1y21GAyA7JZ/gvtGi+j/LpmiW1NRsisb21s0KNE0louOi
fCi0utlfcCVPUT/Ueh/xsqrCsEMx7Zf/ToMLbQRWAW6JGRPqoU3dRdN/I/HkFWNG4TTrIxDjK2Re
lDdkW/6MysVKxtEbi3l+tg5B/cI3nXhZeGwckZtF6P34kUbpkBoNs0MbJMM8dlpZza+2UezdebOB
rdhPo6GMZrtxda82+xSrie/1GNzzPVXwwJD5fT7DvmOEwr67P5CnR9spW2+8vEMle15o6Z96s4oz
T3eZq6nKsvq8M3l0nEX5aN1Dm7hRjWPUT/8d6ue0IZ5c5EnWh7vUOR0Y7sTZLVz3JjE5LXvQw3Mn
s+Ai315nkWQhnbeM58p2sreQRRplOMSofiA8hcEiCt//C8w6SvwwL0m/jU4nOkh6qQJiy6/IQ1vT
M9/n9Gyr4j5J2eJmIi23JrbacsKGE0h7E7jCS5DlqXUzr+5CmlsQtDZ1sfOh9nu0H4VxIErKzqLm
LvNAnViO5yC4Atn/n6XUqbFfY7RUctBDe+ywCFR3ly8q/LCTeL6Gb2iOP0LTuinoJoDcfIxRqM9a
37wRZvBtFxAC5rNJBFwdclx8OdF1eAanagNffxPV+QzOEXBH6Lals9ep559w/jGg+TQpgVyl7GkU
lRo8dkKTUMFbb7zu35OSqsZLQWhaGmIdZAA+MYfS2CXIYy/FzAH8zGsayvaLls+sKVoZLdI35DqM
2XgZqqTQAbRCB9DmDWlRHXGf1s+YLnofR3bFLAM+/XH457ar/YVf7c9m2eAdTe7Mi0CCvWFOEvEj
gDFzy3LBBynRW5HX3duMQMmbsTps5Xlw3FRfNTB1gqNxfHAqdC8r2TF45uGVT4zwrGTLSVtU/sgl
pgdxqhyuxGs0Rcwiy0yDfCsWS0WW1McgA2f59JnlAeO9CsbIGwSvqRtVdo+AmeZD1pao86O+0k2F
CshpHgCS7ZHQa1HGmWJ/9ww2HbQs74zs+DEwNVjBsXuZXViDIZHxY5hhW2LtmkU1cE/MbochN9ab
aGEwGjxkgwoOyDKzMGnf/8S4Vkt2MZ/jf5Hk4TXqAc/SJppEhCteIZykju8N0AOtGjJ15G54JfSR
tH8jeW6UHGKHs/l4oJQdlJZg2ldLovL4jJQbgW+WBzCXEAETGSxNH2O376lP92aiLNFt1ZvWn81w
57RoqwFQhwmAP+95IgXiImlONw2gPMxWR4E4mToEWF6ejckMcBcNBiMAsyHMxuNMVQSs2TN/uUKF
tk9pTThp+I+1eum0EbrT1GUJA4RZWkaKoNpPPJCdH9caZSq27nVLnKDFsoNYaRAIUzOT/SpBNGsj
TMmoDDGCnzORCiVt63zVTu/NlZOqjOHVjSGaat+9zPnAXShrxt/7E39N8Nk6TzM/ICei3D9pUCQb
fxOfQ+i5Uxj5GdItAjBkO8sXJQf6SB00LPCp6uWOjQqGbsvLV96ch1h9eCamTDRFqpOd/QWaqGxe
TeL8xf//pQ9z9VlG1G414wK8BO/LNDaGL8IzeXf6BD202kimb9VkKI2aM35i0JsqXNcNqiYArWgt
scV2gMHEv1QJgtB22zkavKbdnyOzEpqArrPlFJJO+6fWzD28Uh7bt2Wau2Ug1ieSeyUKX1QmnHLR
ebGcJEnhbVGlXhF8/pDDH0Feb35uSn9mJEPuByx3tWiP8gtF+MdnVJJX9kex51s9o6BrfsmgbVYU
2ff/5qgya+nYtvVz2YGCh74GwU91wW0V510Qn7YYsZbkEN6n4oAlc8SR+aZNgVJPMatFeLnTPDga
erF1+OynM+ZfIdjueJnWSSoVm92YYRiQH2ZUbgCBnW5QSkwafyhdttD9ZXGXu2K2X/iFZkgu01Ih
YfHAmK1Sh4t0ams8JpFlnSUAtUCwIPb1V9lSOE2WrtAzQy3O04jsm43ZuoTcFomZBRrGkotxFmVd
boSsyO1uzZWA2ID1OAw8QBksTuBDyfLy9PAax7MhcjPWIUweYMxt/K3VMuQNyf2fphxUHDz0yH5o
+812F2F3jtoN2x80nC62eW3meVP9AU2YLu0XuNNWEOtWekb6/f0sO+N+WyyawDsWq+vMn5DmjcK9
jVz8si9RLWNirwgFPrcS19iyY2TK+K6uIvg+bMaDKhO9E33uuaaF5nlryqEdg14wtdS+JtfJDwY5
pcrMykFd3RavkVLG3scjKhmHH4/j+PBgLUSVzNrwNqCJdn5ni3qKKcAEfD7ChjB+bAQriHQcJfii
EnYKSvzWVBwf0opokjou1a1793Dp+kTlPzFJ/TEScwiLLIdtB53gC+1rbtA1tNtYHD1U8lck4voa
qpr6vLJ4PFCAhiHy9LaL4QKp7BLUU+xq68ItXVkeSUy4v8ncTgRvs3GmNPr4A14Ta+8ZOJVVNoSH
p4wejDnQ8en908PIIcM/mHcddGiF/7PJIs95ZgIfATb6z0g21dJi1ktEf6it7fxmhbm7DcLYzv09
Q4Eg3zftHBS8dGgPg4AuDg3ELkvqYxoLcW0tZsnVJBL4AVBhS3tOCsbUDjmlRDiEN4mFylxNktId
KJDmleY3oxUWHZVA0m4039jKtbmLHSCs9l2BBntZYng8jGWlrNrYQjHvSthAl+KrgyW9yKzenR42
2Dpaxk3XbnbOJDNng5+jHJtMeUViTEwLpIo6JjANVCegc5ANFntKIw/pSyHjH5sNZodqoNafw165
CmEXy1dqPI3jSj5ieW1eko9aDrwE2KYnbqp/uapmEuEvpcaaGk/8KYFOwDMxUkJaGwc09d5b2O04
CDNLqwRB1cSEnmze3eQoyYK4KOVfKdfR/jjY+L+tYRtOawH5WFFAJDf3vSSPMqwSJNuaz1oTDSTA
W1ZVA8YTtcJIcogaBUBkMidVIzefBQ/c1uqqIQtumDF9H+oHrYi+ByEe25ySUTjL5qlHbD4FuItZ
6Wlj1jSgYCpB1TNqRp2feIiQVl2anI3uE0SjIBM/jgjWaKqK5shnsyx0YGV1d280Jz59JomK4ruy
Qmjk/Juttu1kC8YbzakbuuCV2WhX5JVQDTt+pEVSGdhb0MPCerNW781TNQC6VKTGIr93CMAMFyC1
yU1PAVOacoaQ0AWjaelLHvnsZQMzrYk9gegDap9fRHWEaU6KZSoQr0OOP3I6XeCunR7ENTkiY85G
hKcQ/dGUIjILCRjshYEpcYe3FygyU6bjyxm94zMYdg3+Ts7HNJpn6fH0AHMN5xcN0Bd2BJR+CTdM
j4zTLrydcM6FPW7K3JLMP/JwEcFQqGYjcxHKT8FWuEHw6mkxdzTyoW8nrHkAS5MxHfa/GK849zMb
tPNmm/qi/9Wudfi2xosnoo0ABRWgxel6y37AQtBYxYomVF/Hsc6vLMN7d2m6z6MXF4yneCCAcK0z
IseoF/EaplSLKjObWCLHgOQjU8PZiFoFobePsjDc8U0zKDytlbFBhePzyd73t95jYMjWsXbN++qC
6G4OYrPcgKhq9dvP4l7XUYQTp4w94267M5po2iXPi0ZMSJJ8OYZP7DqPEX8G2sslyoUfU5gi4Wgo
d1Kn/XdzO9ZGvSbKQ+USmJq2bYVasMhAeLHrjoqNRhqHTFzRfesM2bVQQD0tNdmyD4qbEsLmKNFX
+vh7B51thorbB08sW/2dvr1gfsK0ONEEHWqh2XN3IuNFr2Q+NuYg4yyOv23qlButg6Nu3qghUCmW
yKWV99X0UePd8R0sTdehQdjXw/lhyZcW6owBBAxSXpwGRXpMf1bgQV1o2NCapTj8jVdBvp2hcus4
KF2OFEu2hyEHMPfG1J07a5i3acr0UDfNBjiI3bWogaPUeRfh/2BsKK9nNMk6rbhx11gBG82Lj8XC
X8la0GRivZivtV0MmT3cCZqCbRQP9Aa+wBJq1PK7W7kJH9SFFnDZ86CTaYhfWnMWklISYj4BSiIT
dPFA0j5enj7ooVTaNx4A7LpSuXoJXQKbLr6ZsYa97uveVbh4Jzf7hVRvDzn/VPDqpiPjcL43Yz2c
kJrGoXLuTW357TyFxixHkGCducVKSUt5sxPMrNN3O/yEHzdgeVhE3UsSYQkYiF+D42lUL42D4PdM
3zT+6zjgZSXl+UjQUuDtQJOfgP9B+/7+fOYURPIeYk0gqJJioX/AtIncDJ/DIAkRCiF69YG/vlzj
ONKC42tWJhy0NNvjjrNKuYVoCvnS56K1n0dpjp0nk1Mb7aPETGla4EnURzFOW4VyMjOhXUYHKlQJ
EwW0Pkyh85JIDZ9qHcBBmAsG9Ty3dtWdGVLkgMsri47Wa1IYf6JRbk1qMkJtRP36tUHit7TnBPKz
fyxqfAtS/lPFaRmuQWeNCaJdtDGW1JQvkdYSBJqRQymbz3u/6vm0YaUUT+2jtOgD2sxyNOX4u4Vh
smNFGFrYt21ldY9j31h8zKBSlDJKTFY1ODlig6v3GAMUOVMyB9UeETYhx7QMYmLgrxsxKf/4SgwP
8tlpj3LaYnP6dM+3myLdx9VQPWZ1HTPn+FZQvNxa+SLgoWzwXCfivr8ghysAAEDOcOBOtq81v+pl
0tfrCtzunS8C2B0y3jenfDgxn0bJou+9PARNIWnQf7ON0xiBXbGyRlTDXO9/c4KRGTuthmg5yblY
t91O+c9cUq8tOPh4lPlKNna4UwHzO1hWuNAtHJSQehN/62P/qyN9lsng8CIkPjAULrfi+H1mRKQb
qrulFf/Jig/xhHIz2Nujlg6OrOsVUnVcbvzjb+sGKmQvgg0eH2QNwaeId8tTI94+1UPlOv+yRk7a
q689hEyTn3XlPjIi74ozl1tLR9DoWj0OmpDaqv01aAehU+wjsOzwvwwQo9EDsZGBFknUTjdbN4TW
lxV6cfB48gWaVT3zyJru+xF/Fuqug5C764jC1zNemM4A7RxAHCds3wHBe7bDf3bvWg4H6ihfDHCB
rWcQYnDY81gOZPMbj3fkCHWzLaEVfcOaBJa1K9JJiCTy6GCvmhg1w1JBCAHwk62hIksX6FNwJUsd
BKhKF/VXUBvUPIXAgeBWF01Js28tmI5XqNLW3/Wf2OssQUnyc2hdkTavlUvoWWA63GVfKlMFDNGZ
PlMfm3yvcfSZgLwdm2EiVnoaQmkGc+ZMxmNDPQe3LSzZUXGuMLQMwJd3VB9zZgEySIqWYdIUKLUS
5cFlpr3nwJ0szBN+4QayrTrZJAwMl+7un2X5Uso7M50PfRTJ8lOEojS9dZL39O9rtPHKA6Lwa7Dt
+hSloHCLzXLT6t3O/64RMrRAU/zttyWlEJ5eYFX5Idze8cScpO889NFjRMRlgAT7ICr+MwM4YRDp
HvfgSzIu76TIldzj0CDALIh1LumngdUnLXrRiOx5IxjrA0KZspNOx7V3bNkpxzn3+OJym8W+szj/
VKAalPDFx9MaEqRO475scDvLjUnjkjqzXQbuOAmfWJPHwUPxw+hn/MO4Qw9GhCimHy3fo31ThNza
0We2kOz5ofdnxb0TRG6XyKuiYmIMQ9EKOacMXNSFhM7ip/GKu9JcsURKRE0Wa3Mir+4EICKUGJHH
erguL5DCXaXX4huqCQWJqH8jVV7p4+lpODBE/AhyZKNDzfRT/TkiBYBdHi3GK7BUrsKMxyPUfrme
/HqM5CYwDmt4poocyPuge0bELz9T2cZIbGctKt4q5pEOrxhpcR/KoVf2U6iKjsKrOdVrfYiZj15z
4IqSdr+vMjvjvpDdnsRcVukHPg+WPMsf3KLpWmvTTS6fqQ1PSuD2vRl4/1c4mzcMbUuTq2Iz6Lr3
wy8H/N6AtYXlrteFoSuOnABQmVVDnUaSLYOWt6c9SfeDEKttU6XP9Gn/j6L+vvkRv3aoGyHpKTHe
ZQUKvpuuBwe3b7BtEL08hAE8MBW3Kh8s3qkodyOFbO86JxpWE1KtLlOayUMJs+jEFKJnJgXBfulo
EFZGwd8LgzdHnOTKYlhwN641VyMOOxesnizvNCZfZo9ZRZgioTMRjSt+sLKHIxrqbgldiB947eiM
dMPCchqZRvLo+Dlvfd2ayilvPRpnnhTkBvPk5Ndsa5HNHE9eqp4sR1uCJDAD9Muwg3LItWp8YMsZ
CRdjXNRbe5p2X1Xij/nD0uMFdMig1cNqwNsU9ZFK37EkN96pd7VdDv6MbvpQxhueYHEmclcTR6vx
eToGzDJS+w0yDCp19JBqcWwUM1zSNHUc6zznm5QXT44KuS68lz/o3j57il+whTCwajFlUMuzxWPs
+ixkB+wlodbM9nepmdPGBDqlC2aV/NjHpSEwm6BqWTcp2jXvVh0t1ESXbxZ2jrEgs3XO83tljm6h
25nw3vpUAQjZRrbwWqcK0X+78eC/W6YwPxwJh0jksrbddlCr6+f2pA7JFEq2udMdV24XTVKgvZOK
NuG9DcmLJ3LQm/zd0R/BXu4/emqkUG+KF9v/Y5x7lamBOZxTSDjN/m7p9EbUXKq5czNiELEcuM3a
DMguoab45DcbAzW0VwGnSHOf5iy2qGSPBKQWEh18OoKgf7dg3dKf7yCj+QPJzIpFlwUZQUItIghH
+iP/xFIKLIogN+MEm1I0hIuCPtScEXQQbf+HspEhmymMn2gISazc4/acNMJyHr9G34THSa2NqBKt
FAWX6Jp7dnQcFvz7KpENMvmZeCWFCJFV/DqrmHVsbanOpLJK/7eLpngjx413rzNzAf3SX+rm9ALN
iH4aS/0dN8Vh1sA8Ktk273NcBF0FLtkcBWeAAR/CgkUtBU2k2aOUMqwlxV0SN/v1a8201Q13HWzR
XW27bEYBFz2alW4Af5/KL3fDGaxYXYhOIqI7Q73VHJ1QPqfW1z/teq1IRZyAprapTkJ5fq3ZMEuT
NhNvznGKyxm9atFrdKGPO69leUkb0gemdWxStIR92zZsrlfeZus9tw0pft6x6nAjc4NW7LiecCMJ
eMF0n6N36VOdqd62SbMClacqwuMfsIpUVg+bt/wn5OuJk304MHeXuWf2vEZ7f412if+fDJPwpwTx
+CdCdj249J5IIlVIdesgBZT6ZS5uWn1zBYrRnERV2MQt2/OVg2lGIYCrbuKzwznPNU1R93eUpv2g
E6vgOJuaBIr/i3eFtkVPzb38zmYEd1RT35G9GrxiE763lNOtRAEzLyfOOh1f+Jb4PGoziGPiSqtx
ZBCxCIoH//asmOImX3Nho4ahQ4NVl+g2tevMnr57mL00WD/2iHzQMlq92Fuu11/0TVCH8glc9c0F
C7NWoj5sr9XxqDN/xd0iEgcHQ27qDSRNycdbN13RmE8Wu1X555isXn8JP7iNDdmgSdXYW+l+mKe3
Q76teixgM82ySHp4PouccuMXNGCS8NtvMETLbGydONkYWhNB21nGmkJe8tGgAYAZe+iiyAQLFXwV
T7mRG/jAevr7PTP0SgNOVgkiFUPvIqszfNO/jRI1Wgu/GP85svjk4R9+03E8SW6Rn+jNUeCoZD6T
vxH8Bk0L64YalQ3Z85wz1pH0w7kEvTRiqUYNb5yq+mGQv2qhSDJGmGBfqzpPFXVWe3dk4JwuPmhG
Ux3fnF/OyTS+2JJDf8Yh/9uYgw32HymLabc858OXqCUw5dW3La/BPX9k+xLcojcRo5ZQR8j66lbJ
VTxsdd4aJvP6uK2xj+tQ5Qpq6W4eS0NtsAQesLqZ0eo65XWIs9YmB4Y5JJ+RSns0jXGWhECDxqRL
3gf+Ckey6311z7ESxN5EvU9DQAfRRzAalcmGAKL4yHz9eXWFvoBpWRt94UtRyhgqzj+6O6fbI79p
Mz33F4SkNRkYbVT4q1Lk0cVThNGPbdZwks9SPFTqYcSl3ynf9Kt+jzRzX9p8NJ6OHrg8LDHcAIKA
6Iwg8ioMaTIXncQuWjz2Ubjh8DqAM+mdcum9XcHbDVvUGfV4ToYdW+6ALDRrbDcsEqgFfEfJy+4B
IQd4a+RmliYpXUNo9R/1kVGHd4v9Gcpzb3S8vy5czn1t9QUJbaDTgZ6ihZiPMtjdE3yce8RIz9iN
EFXyTLyOZPZmEAJMqShz/OEMoKFpBO+DWP88oue+82nPItu2Oghvhrlrg4rM/quDDsALNBdkPsBG
tHX68jYXjnrDRsCTZW39CLqz10gvGMkdDzmHRYx3c4upYKbRvi/NW0DZaD9eHjfPysPdeg+iUxcF
4sEl7LQAXnNV5grrMe3DM6mhcFxV68Gd+CmQ1ug5/nxG5HPbWM6se9303gs9TK1OWOoRKMAy2m/J
sUGSAOtGLBOdxf17nxz6pDH0VGl6XAp+8wBF+TZ9KfYhzClyu6j6hx7BW8PVeGI6EPqIblP+1RqT
qyqsTxWBRsDbUoQ8zZiVyvIyI+8hjm1LMgdiia/C4IfCH/7oibjL9C04q7MThUebr5PQaEbf2BK7
YcsKNFukseWXzvxmiAif5xNoomce3xDoTX+/0zNkTtDF6Idx9lCAuNBW7dWTE1R5TlsD4h5/tXeg
1sQJyfyAV7vO+Qhh2vmlVL3S8ylC7AhxHNiHjDipYbdVrZqpgez9xfvv9fyy1OKIUbRcm/IzDxKk
LH6EGx3ItmvZa1TjpvPq9bOjdgcsFvYdMb3MT//yGrmtcmb8pXq0fTnP0xt2jJuygTYNquojKTkx
sNdMxm6KDgfFHwnJrkkMxDh/t4s89qb5QEAr0VBxYSFoKhNpzjZGONOEJFZpYOs+x69rxJkHg4Ts
pB8IrxwGrbcZwqn7t7LELV3VYWcM8AJaUvcXXE0Og7t8EOYTSNRnqyC3sTnVoRlsEzw4TD959wEK
kvhMftHlDhEsIKPP7RJ2eAwW1DwSxkaEz516uZw9MwU4Nai6fyKb0grtzG9qD5aBoz1GqM6D5HER
4y8ORvTOnmuGV4kxQBkE0a3WlFSOURH0lmT/48irWssCZL5pviDY0+MHIuzcS2IclPEfmfOm78F0
woUJuLNafuakMRuwPBsh7EDlh6wMts9yqSplN2uUm39ArEOrxcNXxSNygVf1QH1Eat809BcZjYI5
FrZ2C1ONIW8lDDAztcx45E6UazUiSWAZhtYT41Q3W15jJ6e7g09OrS0FcxSZ52okuaw7Pd9Zyqh5
jdqsovZS9QPRkyMAAUaIGfL9u14ThtJG4Zj9w/OT0ZUR6CmZiC1LdWXYXTYV9lt6L+4NDNx3zca6
yHAN3Jv+k5aPXx1q1ywuqcgIvwD9ETEiCnbvOZdRXilIN3oykKJ8nnGAc96ZZ0QHcsY/Ml8eVKRI
b/HIR1aopwAnF7ineO5XRJua0KjWwMkOgPgJzchrAwtyaGbaTFYsxdGlK4digRQ0xVkzYTtxTP8/
+j9jKQ2NYDebtlLUaQ31EgPNiFPEoj3dnxPL/qaS1SiWogXQlXb/yfk1iuh743TptTax92GzO4We
aUf3MOpe/sTvQQbrKXYltmAsbVTmi1+YdaVgx9XeY7HhuG+3CmKQrp4C12gi/9xluScsZrVBu6L3
VpXS89d6DVfgrAOdlIz+iwwu0nieNdZiO9lFu/SMiYXqMG1iyVAEQPLhKm2r7wnWKf5NGbfSouty
IY73TPTnK9hch1jRPfB8a/eYMhjualoNISYGtAT4jupiPSbDjh1ENdtIc+TPSylgrGmke6jT46L7
5C/xLHhpboX7K+229kWnwV4a4Dt53Qrf6zDHyc0vKLuUeEIbmpw6tSIfCEbTScE298aeuA8+AObR
KWuw2hCeAH6+ThoIkHgcTe+1k+/7ucPnHbLRz9DfMn3tG1V3fr8MK7LmQBM9gSV7T+UZjfllBV90
MdTVMx8siIuEijbRFbYQK/KA2bXxPA4DFoe3LFPaipTITyauDPi0sPVASJW/FWtrRvaJshZHOSuF
eryAuSOx2HZuf0t2K4ynEGrWCXeygV9EAFxmZvfIxGJhRVuu22pvjS4Doppy21JHbvCeyRkgSxzc
fW8TeGeJid2ia/WATIbryuxXu/h5VgNY3vR26gqvMBcRhBShq2euyI9vEtnQZgh1Qm2VQ+hJyN/L
8GCfn0qriV2B4XpEiFxHjjlbN0wctYAMDoywGfeskNrvZwJ+oGDtFvwyZwewsp7a025i2nWA79aG
lVKc7B41tiDaCON0dqf9nmfMwegTHw6BTbAc0A4Od/US4Gw7CS5QqMNdWrnIMjlahtAgdsbmN7+v
VLZCyjhenvsIz252p9ZQ1/mt+hMLwjmjPUF0qAD9zp/4yDQxjYQo7SUQrGbQy2D3ZHJx17Ojc3fD
nFTRY7AUoza7igP8BesbXmQT+DEJrzXvze/rgMJE1eShrzCBYeZAtLWuAY7ET2WAqPlyASU0b4Ew
RGlDTTVpJ9wVirBWmbWy84pJuzDhHIAmLPhUoLo+WdCFD+LRrdFd0+YCja3uVQlwB8iY7OBT6gx2
aJvVprUvl0zryklJ9BaMLPwyqxsjW7HhT9wGkFSaqtgugFcOVHb/TMqp6k2qls9/Km+TJGaXh6fw
gTvn4BhUtN/QF5XWjS6ERkeGyGV04AAX5Yy8kkihQCcsEu6h4Zu9mf7SGDLckzEBp1k4StwaJq2g
Wt56Ho50V72uNHkuSlOlVLrurkLLeF/NTUVAnqiBnfK4VPto+J8bCxcfLza+AIeqB+jV0NMT80sj
HFL5c6AENe76czqxBZp9EJsbFf/bWxVePFHVqK8CjBH5JHYGDdHrknkv9o9S96JIdmDEgZJtJQJj
7ScZ+95r/jbn6aBttrleGjtrNupYYeyRQwpoQijNYvvoWgWUQ8BSdrlsXhV7po715kGbZSjAkmqs
p3za9YhMW1UI4Fa4NDihLYS0UgYBrLCwkffYWzfHdgxVRjeScbrFRkyTQc1Dt8X51dDjziCCv/d8
zjXyeraAbqWPgMQJHh/wogtT7KqVLltsQsHQxF4kjGHzfsHFuRS4mXM2SejVHKPy/jtn+vLhdHQB
NsyXVIBKLNlwggLIkt4X+I+kKVnf9VoiO+5bCnWj7+U2y/jlRcsi4C7N0i5AQV73E57o6HUHAFcZ
mDiySXqqo6QOmMDES/jr57mC4YLjdg2vu0T3r4JCEcQN6cowuWhNgLG9jbk3BsnEA0mYd/68t/gd
+ygUN6+wjv32ihmRtXdvtXDyfEILXRXSZcpzOkQ1Hdm9rp6t5GDaZkVGPwvE8qIHzvbXrQEDzvFy
mlKhL3tcV6QoCaXeLBWavkelNktJnh3RrvGpNZoBgjBUKvW3YcZzb2PoiHAEdoNFninGL5cbIz73
1P2aswWV+u/9GdlRvkVV7x4YPDUD29Qi7RiRaDw357kcG29fka/gNNayYXIkmGaX2fjCEvbOnjXc
GwLHzp+9S0gK2AhRTlgCQSdorvSEzOsR4PMtfY8+QJX2ehHO9+0P7U5ohjjqMuTsY3hAY33+dUgL
12+0AgwOq/lmrFdorpUV9pRK0pc1yPwqBMPmb7LTWZsoN2oJb/6sHmC1RUd7KN0orHQiEG54Yozg
ByyxWKVlOXp9YMYjq6lLvXkbgQRJJr9GMnh98ymQsHSCBgMI0tv4md9pjajJYfIQ21gHviK9E7DA
0XjLBMtePCZmalMe9uYDANzquk3/OWxEdPCDHkDp2i5gTqb3M7Y2hGKlTtU7QSYq2AG78DBXI4KC
J5lSAxBtPSuKZ7Ou9JWb6VRBP8F5W0R0xeuTbXgHUIueelSBVc9m6zg8oNCsZu7eUULyMfXBxuB3
o7IJ/MwH5DIHJTnWx3wOVGan3HOjtxaEkOH9aWnlsuuO4GsRThTFvKhHp0+LPNqMUxxeoA9hCfyu
3sVE4Q9ah773NVJ84AVL387guJMqHfb80czTMbpc21WzZcU3pGVRPnlEzy9gIF5FiH0H+lEpYHFj
zWgPEZBdB6sEzjPxFieGP2D6rJcFkzIcyWLD4PSQfc52nZC6H06zlBMaD7RIEcch2NUTJ8MC4jJJ
KLRMnaOwEV4CNABrAJa+1feF+UBsvy17DPo6f3SM//w+oOYIbqMEQXX6qIbF4EdOdUtOUYOqg+tC
6nne0IEmJIXgJI9dRVJRgn/jO0YB75x0UM11HKDSM/itLlQgraFGKyI4xsLgbZLpSYdJ3QxPtmcm
8AM8LIIs8HiJVPxeho3Dso1rhf67YTu+p5S8sm+YbcBq4fUzqMPxbfu8MO5Vcxm6xyJ0HGdJ4FYQ
caWAdDIzBI5GzRTYYPmHuYG1Blg+9wVRZ2OF67/JWL+N4PFq/UmbmbKC0B/7hlq1gzEgdFncDrdZ
36DQHYRwVISIpx7ow//rLqGgeo0KvDAtelwnd7EY3UiyT2P+7Osb6CNBxApOFldjjKiXxP/uWRZA
nTUc1BbMmYq/YmlJ3mGP/bBEL2X21mliC0qyIzuH/HhpHEVTbhjDVh/JXxM+DrzLDrG1Eru+8z09
uvqPZ20t1Uxe4yuFWw1DNOD3mlSOagmx6kn8M9m2GrNvZ1LrBnKgA3ymMMnzCVbF41V5y70Vtxud
yaORL2CAziQEdhvNR/YnWpE5MS9T9q+3l95z1lB85YMuoGoU+bMfdkleNa4wenyuUYSqFzuszutd
UITuUEm7WaHyf423CsE0HF2qj6qqZ6p6JVntEB85iS9raHQ2ZMHrTs34QHbZhy7kMj4XuFw0VGXQ
vGhrAwtPFdFedDX3qGPzFF12WaUmjcrfddEnEMJVC74b6z61ZWEBgMJ+m9IwLFWtcyTu+1EsX+6m
fo9Ybqyxhrjme+SCECDQw1fbgNoDK6st1Thkqq2kV82bc5d6FRkuo2516c75q6h54ZuriB020NhP
khmbB0G7UcQhLNFlDek6XLEkoW6fBoWb4pcetUWMjhAppJtNgxYnfgfi3E8AXm1vRzffLcTY/M50
hmhdp/94xUaF732lzFDCniDuTqKJAWYBINjeYHj4kxWkPtcZXCXwhvpbt3b2octD6lYzJ72XSYYH
BKv3mLqAfJn6Ou6CZ1h0Lx0RXoNm6ykVIsZ3zvWCdfSCsYhRYTv1LybQ4Bv/bZPrDav0BGRo6jZ+
vCuYJwotw+hmibhoKNsNZZ/lk+/j5eEdvLER1rfZaCA0144zbt12DV7hDuEO9Hw/BsCaDfV3hbKW
wkA6xs+9EqhZkmBgirtYb7RSGRY6QFcxzvyBsZnhVADwdPUOx39kicyv9Nxc/suQQxrtdLlLyhrw
F4189uj3mFylrk7+kTiwfW1bSx19nQnXOnGU2T7xA0dL6y5IeXQZ/yx6SGLOomeur3xaJKheKhM9
dWCNsC+AX7ZQfNTrtDY61Z1663C+XNaGbSL7nb2hVfqLXHO2mwUTL3Aox7VGGb1YZs1OYBCOHJyB
zodIPAwpGVDVLTOxOXM54V6SSBaUsXLrZHbDz3FgatnnCtX574MSTcW+99Gm7B37vaue8xWSouGX
mX5HxnN2QcUvhi+ebIxUai8y5is6E3fGT+QF5a/i/4K0bJF7Ssax5UMPFRwio+hVBiWG0BpVOxDt
s+T/BNR3qvZSihLVLKP8xrobzCD9ZQKeevd+Y+yLEBb+4A7Ng55iChVZrzOTpz06L90aczB+j/oR
YMkg3gyHFgakOqgug6iEsvcTCGrvSCYZHwXK34+DKj7CvK3TEj56/q3nAgxwrUk53JWWWV3Bgd+Q
OcfPva43NI2I7oNytSd263wsYfbZE0L0AcHTaspLzG8vQq1ezmQ5jPdwmexD1nOoSXyCrz7+indm
gL9zW+exdFWm7FwI1IQ2AKtzMGp8UnXOInz8N7VLozlnzyvLafDtrAHdxXwXHA7lWEct7o9UWPHq
B/3WBCnCksEuWkaIvshu6mPrJdMX5ATIkliLLNab29BtwGPvyQPXeSKgRaBWhFQv4gQ+e5dLNct1
LAyXD/B9oEncVDSsQy6WL+zDT45+r3sepA6Y3WRnLWToksGkiGwNrTWVSo1NeyR5iZP1vYA4Hucz
BMjJHzPCTt1HprieT4YKxxqqy7VqEgKox5mtsFe47hSICvx+UGvkjdk6ehSO6K0/PPpZa/7DdWNw
VyXyVlemFZxigDvbas21GTlPjl0hklQfj65zYiPykKX7RcMGgKZ3vJDONdlH7PD5oxm+Tww1PO5/
WoD4v38QC14ubwi3WUKDewjatSsfY3h6CuWm6lbuEdBw+OUqRV06QJQmHqBLIUo1w3XC+N0eJ3+j
NaguqMfHrKrAv9F9vtQQ4xrWyQl19+gzIjNlx0diYdL/AYd6MO0OUVWlxL5aSjWnJGlgno7dviUA
Hx3+Ki8BAKjX5ZAZUiHsoG6bimvqpZf5kUaNxcVxriEpr0vCA4Bbja1PdO5pwzANRm5UIe46lqMw
QU8lWIHDTEkIbTlTNlyIxgoWeSedV0CJqG+b0VABS3ZLvFr4qP7bvKtKUawdXAdpPsWEpxJwaNsE
vBq+qQF3cbHSbmxmcjyLNq9lVgKKW10FIK4G6Qpa4Nrh3ujg5CfEfAQorsn3PS1Mpl6NBvddgKDn
jtDcTdy7cpH8bc6Z6xrlK64Y2+AIFheOBg/xC3ZMLyNHSxhQHmNj7lcPjpChSn3g6fOYQavSm4Cx
BCLUCwJ1f7kHhLgvTErQVr5lAUv3dBDrtw/4sjjqC/1pxTZ5GXBrO7fsq9NB4Iolt8+zHZ/XXob+
C8ZRV5lTgHqwIsBola26HogBKmwRAsdNWLQJMAU25Pi7otzE14vXPG7HByF3mo0pJchSGTJsxmmL
u/4ckRx1g4lIpojTrEtbBB8H96QZxDAGng9TjBF6fepd9TvErwMJ7cfc/Iv5jC3bDwKYpO3HKPwX
dyMOuy0BxZdKxpiuN0lgA8Tq80RSn/EtlEIF3M0tqiNEJUNL1PP7iSn2VWTKiN5QMMIXgK3+4rZH
FfwA0Di4qsKgq34qAb/kMnosgH8ocs0iaJm7iIGVUK86N9SSbtXDTkbBReBoLjET+1knnpipA786
EmkVEX/KflicZvbGERYO/7CswHBjg2K6qvfmytxNUTCWVWvQNYv7NERIqV6rJeS9QULplEW1reBw
zz0T9nmhXG+NDZTnACwsLI64eZvdrNwHof3pWNI49N0jmC+e2r/cjPnc3sIy5j68mpTLZk0aDNC7
6Fikptq84lm/roN+DaoQBub+AaF67UbrOhNXRmhMm1wyoBrKZ4cFFgWJ3ZfdAAtMFgyfsbN4zcv5
mJVrVt5ZdsDdBzWSpDe1f0rZkHfmP1dekzyzr5gTZSPOZzijToweMcz3sKoZxYC8e7RCwLFTapq5
nesEQaGFz5viZa7V2toj70aZ+9E4pbPpeaNGcsIXwSQGF+HqDf6om8rNNAQPWZ8qTSMx1Phnjwx4
Mkl6CI/7Ack4WYfFnducbHLiNU+v987S/C+3s+L8c472sJBAsXkuhoEecVodKpA2zTm+OX01xlCI
uW4CCUDGbF4sPKQaYekIu4OyFORviJzIy0itDum6SfemSbwOM4hkCU3dZjkgqDg5t6ZsxrWwHDNe
47GbhXPXppJUOsWDQgbrtUDLucW2O6YoCRYkqPVjQXTzez4ekHcmZ5Mpkt91LgGdSacqOUc5inFI
lqeOtzXE8B32qQzSkGEpGwnpvnDk+x4PSSMeOUW6TOjME05kFDOExCM2MVDhodvvn1GhZc3MrS+C
cUhsSB5WvSZfshJI8D6miL0GcV4Y+A4Ha9HlXBQORsxai5OTK5xpyf5W4GHzfBRqoD6pkttI4FzK
jVYmZbB2mMaPogtY4OM85F1ZVPllZGMbkGIMJZnwUYzdYRiptVNyOMYdqwPptAsZQuFecoBUNxvP
dmAysLh2Wngu9zbL0FoHc81Xd3hICJ3vj8s2JcZ39VpHPcaEzYxnZGe0dvpd1Taiij0Wspdd4B22
+3xZdeRAVjn0EM0jBbpQsSH8ScmcXwV9ohFiiIMoqw3jjL8lHUPywx+I7ZA8Nlhxh41eHWOyiC9r
gnsMPKoWH39xP1UHFGO0xZNMjJGFxPgns/cTeOz4qFMuc9T3E+ab8d79xWwh/7LXzhwnn8TQJP5r
5Z2ta5MKswyw1MTHSyq3168ovbZ50IRmgfD1DStEL19V0IzxFC/DlxTcz+muggly1uXXwvPzVgBZ
zJXcPzJZPG3lKz2jD25kM0MoksLzfnmtVXoonUoGKcrcyMmooIF9fDR56ZNGy2tNnARugBA/mcgn
95Ix6ZC/Kuo6of2qGg4VYkrs6LkWcLsBNKzRRZ+OoMxt/Yg7e/4gzVZYw9IPkhzIHAsOBqJttuIU
E6D+SYApKrYCYrps/J843I9E0USdosvgkLC3zu9JQnCnTuAwCg56MbOyQmoB7xhWWO1pJUVgnHvG
WztCrUg+fa9CoO2DLqi8R49UeOEF1vT5e45QmqF95alcCQv5qrdULptDEYRyOXuPAsX5psvWMrcA
wXFCSMb7p0PYnXawiRM27bekqDsNatky0mmB5TxcGq9qcCRYfxneeghkW0F9K9fYPQOzqgs8ZYSb
r3feBanqKBghcZbz645VK7DpQjP2tY6fLtUnaoqdgvf8cxe0DUmgovh5KJmFCbMAVd0gHmxezOsf
ql0YchnUFsTPBowZLbD98l0AxcIvbzUVwgtGNLHF7LZDu+lwR02rkm30hDJ06YkPtUQcnso5n0NH
hx78hNnul7XLDAFAir9GHxd7n3Bo8QkGScKikvKjzM6XngfhYCHdUkJcI704ku2FPbFP+oANe+A0
Yxj+sxPq/uxoU4kMJ40AOic5KpKINyimyya3L/G6M+sncXD5GeUBanLz6ZOYaldsBmjY51uUNOxt
kN6nQJb84cX1DkMRjX4itc8HH2qLTIVQjLIv6246S3vPT3S+7emvHpOeRfj9b2pPAGPsd2UkbPXG
V1pNXXEgo7w/TRLagzJ6UYyZx2vGNXygD/ppeCDK/gnBaEcZWwxxtQEEcSTolEu70pCumTGotmXg
fXAq/WvqfiEEcmIyzzwdYcJfvTI6DsNL4+5dPqXPxdpo9aKx1R9wonO+msEGSWZpJoyQ1Hk7peDE
aS/eb/jx++2bMna6u48QFVgOSCpqIH6QuhMUBWZiymWbBPQ4vGW6ucu5djdjya8K93Ujzzy5xsoL
/u5pMqmuCTtE+spuuWfGshEnG4Rg6CL22fgwm8HIRSSv34hf4+hSoxnupALgSInbUBkVZVBGpYhl
gUvm9a5RyqUi383i3yyTFr/nt8J20cEBzAZCSdwbd1ugxn3HtqpuDwCPB/MJG68MKkXTymBL2O9F
4EWUaErPswEGS87SMWrCYC/I2Xtm7+Xmu1vgr93tVXr+r6np0NUeo+ltVrsJBcKhTo6uHt5gTMzd
SASc9SxGhH8XMfoFZFl0nu8dHx5EpeFmv6ln0OgyVUU788PwXz4n27G2Yo8HguR0zY0z7Ec1h67l
aAKRwp1A2SNj2RC12GNpubEwX3dlrAv2IHVg49cX+m9PHFluV1ngeHSbxps1L942l9Y4C3/LkD7G
h3Wk1MKUuGKu94z9EZwChFSELV2KcivPq5kXx4e35dd8A884cfebwgTul71fMm1i398EkDqa93yw
XINkeIIp3CHNoVoHV19thGWQVBjQFaqjvphmR+3lHgsQiiOToMjzyTfTFAU89yO35Ba0sPqplxlo
wZ7JHZBxh6Kx2bTLA9rAUPWjKZlKF5zbQzX8Np2P41kzhmpt7ltl7nbkEE9YepGJCWUY4CaFMuGv
+y5ybV2BmvLz7ekLjWqVUfW2Dn4AkSU15HOhRzD6WX/AjHKT92I4dLWZJnWOPAQo0lHPL+rqku43
iho9Z3vi82j61maB4sDGQhsXzZzjMTglhB0gCGOoYWoFbo/Orf7DuNSS5wZ1z9YXqOcWdNlFEer3
4S9IiWUPNR4xOcXdnbcYCD7oJCJgTEqqc+Fxy4FkzUY06uxDB34SCeWdr85AzHTHg4y1KxRAiijF
ngj0ENMIIIWlH7BbxO0BbqhO7c1zqK8DhZ/SU4eLKzvQOP+iPMKoBt+EGYntnRtmV7tGTHTrrY1s
56LZROmkYqJSejAEfbVgWo1PeEpc37WgMt6M9tqxTgyDmcONKwkDjfKca3uBnYCEXmj+F1K1aHHs
owsNFI9hAxhYM6trPMz/mj/X0lje1WbtcxS8ii1WnCr4bMZNy1Z5gW970Eh4LxzgQpXrcnDLICvC
38uQmRPPHpQCnhMHfI2Q4IvkNbJpH9ZeJQIJqGsf7OeLPmyWgd74RZp6YJL7GT9Z21bWEfvmfp1f
W5RRM7jH07kf+88C8ir0MYPIfRScfgNFHMRlIk2XIH47UPKBPjLXRTGWVUq2UFAqj+pUgMe6VW/8
jpMY1HygwNVzTPnximogjWF5ltUeFw/7QQOZ3+jf3uq5q9KwoClOuXOStYQnQFNtj6vkZghSTXWv
DHc46qnTddHpMeo9er9MxjCVfK2xJ8oOzzksOX+K1g9Glh+bq6pvrnjiew9fW8Knk2lzseFqUnaF
6lvyIoMolW09hZqFIgigj/Jxtbi0yFpChHDkKsx7GkjsKoCPe5lPIWphZoNYb7M1Cc+zeFQHF0KX
i0DHTSfpVllnIgWG+KZ2E6b8Uz9VOtM0zUxDqx9IkqmNudgm+1ZVgL5YrvI8FasqlM4jjm+S1hZS
15ipzaeOanIZ6DE87vSkxatIT7FK1WgFhVxLnUzX7wSgtIRPffOqEg30/qHQx96N4Ig5V/J9+ItJ
rxIzYKgR6/K6nO2q0l/2/QVKlgnSd2Dc58PQN+zHjkuU5q9ynAHCQ5CbfHDL+lIP9NIaCNHoP0HH
RAJUbU8Uvv89p0gyXrEKo0kFraq2HhfFnb4172k97lnPsJct1cGNXxnb+VxCE2IYOOe11ocjXki1
H3BWe115thFolrp0CG/OqEaDs0O7NuRyF1NABwp11ZLZW4yxbRTwqjI7rgOwTtFWLCh3ec48KE87
RlvraLC9biL4y2h5NXj0iSt88/nGfPBrTvFcteHnGtZ+0rSwii+2+OfSaGt7DUkHcQoKyytazBVV
QOBERL1sK2mxEAbeLlgl9vy+dxpTB4mm88bCa4JOCcU8KUwaWeN1t/G+EeOyKXCRFOEpawdegkaH
GVB0wBeKY8JIxj77sVIirkBS4qZLIYiV8gnEzHNfTfcG2lcoZXqAVBe6qdKh8zVayUXk/HcLnV2T
+H52Fcv35d2emPdJbwO2hVMb8kn0XYKPiPX12utJ5OEZMIDOty0Rz52GWdAD+CgQmAYhH7/fL9G5
JsNec9q1UrOKp2F+AlPpJFkIcUL3RdbK/Bqap7+37suHYvmJVjoHoLTXb1TrsBWZMSbsh1jluNNW
+8ihv3m9adQ2xj2uJKlgTP00Z0SbHR8dW9476Gs+UWsF+7ICRRF3M07CZh1/G8gkRq2raj24jbPm
gmFBQ0LNlrjtNbQ93vzF0Xk8O0hbAUp8El3A/QAJ/fM0WuQduTXsjITORmBXGkL6epKTgo1UTXU2
XHBALa7+YNc9SNLDcH4tzCljPl5xjv6758uDzXpEhh4lVVciqiUB4FbS/RqpUWAEzZBfT+9v3hVt
lt79dxyXwe1NTVT/ZN8jriOcezqtIiktEk0xyhLemtK3XVK6UkMVH9jw0igncy3Rpi3N+Nhd/epp
1LNELSDnC052rcXvRkDKTDgUV1FNsV5U6mn2uBA7O+FE45JVDQxwRNXN9gjcqwQJnDgKsV+xcPZv
BNCQqQz1zmf3FA5eMv/XZv1gs24evHTHLliJNfO8lRTPfBhBadGmn4vrkugMbO9R7D+Mfp75OSPv
Hr3cET6kHgApCexvqUY9JJkvoJySRrVpsv31IE2NpuN8Ynz9FzNRQ/baIXbKRhkqMeNBm0PBRX7R
ldv8ce00U+p+g0ENDdTahxXQChVRZAM12/3RDzhTpCrwPYb5hzsaGvcOfNY1pySVdN0/PbGlnFqO
cSLQjZkmyM1/Pojw8y26b7Fw6xYhgRLlFhwarRktoD9tCKZ38EtpKM8Uz3ORqkSaZt1+9we1G+Ot
y0Rty54rvCKFkSdG76llQXq+tBUAbKOxd6XlHoWGNZZHnCJanOFZpRW15fvF7p5aK6X0HqtqLmbE
PTVDt4tDtARioYRjGhKPC/7KPoFeBoYikCGNDal7P37YgKFIkpI2NFuMRloghwCXS3A6oQPKXbL7
1l8pteG0dAU1N2W1XBbGjsoFLEjFxlEetp5pVgfTrk8rpIQvGhVmL/My68SzuiP7w8Kpp5AWqu1+
H53WSZUSWAOgCRKpBkr/RYwiqmbMcaHuTYqf1fetHOFsCYgZg6nALAj/pmwHkXtqvQvE4CTrOm1q
DdHeRm63cibSDeVEgwd/yixAsbgw79iN8DlNhvE6XZckbOkGxhOtUCl0he1/wL1aq9GENrtcKg83
ElV3HpFmcWNWEt5PP/mLOySKpc2BZblHRhcfKlPEg6pMTu+HsEBv4ZFbIIpuyYXBW5+70gOcnrJd
tXE1FuKGIuZtiwngCLx8cAB7dJ9PdxzqP4lvCwl1Omh7AoGP0f4E2KzBsMoQY5uyuhlehL3nFG2Z
ZqkbYxyTM8eG/RH+upSkSr1qycs+ByvxtMQ7Rk2Ltn5ypS6K8oG+3rOG6a809w3m2p29zxKOpyRt
FsnuTXJnAClLr3FpvmNdy2dRpC9FAJwzS4ThPCQonKVwBaKRV/3bpTXaHp7dJ0bBRscq8F9VSjda
870ve2doQjV77ELUeOtNnoQDSHLwHrAs/ER6nHirVfmtMeKqefgORbDF7/XFhktqCkcIeQSJXI6u
0HvuqomOJYSW7MUEPe85r1B3g8qENgGAD23MHbDS7jaf2PW86fQFx3OBI9vh8KNsW1TWhFmY3evk
H261QNVXLhoAhUNOrOKP4L7da2IQeruPsmoOD7aMN5Fu8AqHshcSOe4GoHhu7sNrNgILeLXpMvr5
9pA220whxbQcCr8kPpaClY+tF1BZtMr7OEDyXTN0DU7xI02KMkN7HTMVqfYRK6beU8Yd9C07RUaG
vkFW28cLeTGoKA/37QxFR6IRRE9lJwuQhz2RsNcVuNxmWZhV5KIiV9Sd3LFgZ6ak7ndYYFCqaMqk
mw5dlwKyhIf8tsMlqyU0iJbRHlzKsEXsW3nzQg3tb3XJy133mxSX02CiXhji93YjaBCT5X8cacrw
KY/rfK0IlAJiIajYGvP+pIYm4EEvDDs0ej4k1Qje8Jh3hAGDpx/xhTDtK4i675hRR0j8AMp4u8J5
u/XsxPIz7O3MYo66ASkfyoAqQX2ufM39UqDeukVn9KnCxTGdPvS3oVUsAqyImE1V55aUB7M+GZn8
LM2+6dWWjHfkCZpENWVBgq3vt5QVQGO3CimQ1R2arJ5lUcXTe8vj4tyrGMcQddecmAHGtjFTS66z
Jy80DqV27wRbUHVKqJv6nK4gdXcESVAXVOg4qqZzdW9ORw9PNzNQz77NlqZMv39Tm6iN50Sp5pox
54Z8Zk5gFOKkUSrEk26pGgNugbUnOeWXrHeIZ9ltv8ZvCfun/H9qyMHwyyx1AdvGRgK+XIppvpJU
f/DwJvYi2vuLwPW531Ph5/6uyyr5toubOJIUoccKf4F3CCCZaWg8Y4wPuGvRE6Gqgjaj6gjyTERr
HgR1Tt71b/2R/GHuJWSAeOiPzD2j8NZ2qwVdG5XTW8l3WGuC94/piUSyxdVwXNIMQF6kb/ngBJEy
L9+tyziwKm/o0gnFlnVxPteT/Tw9qJbDe6OVRicjs5gK1EGPAC+ESeazYtk8BDMQ1vYEzWhBrskv
TKpbSMUFsH/djOZI8mirHRNTt/IbNo57aFFWEHLeBwrtTJvrAXB3RFHDtbtEunylhQFU1pAxg5w/
66FhFEwVLCgzdHz7Gq4xP8HiuOpkFzwQwUQKqSPjKAGOqBTncvYsFlCAre4qywo/ontJsToVHk3d
RzYKLYo20uFDscboRtZyiDwgQTxZUw7gBL0FSBJug/VBUrIERfT9qZCQGjPVKlNxabISDfVM89Kd
JCGbPfPY81d/eQ97IVOHs1bAeBZw4Q7foXhGHZOlTUVvn6Bd1EWvHra37Q388pmBzqmfxRq96h9E
1Ry4WGMYR2WOc3+8ai1LaIXPsTxp9QdZ7kx8xmA8ItjapysaX5BtlyU5lwQ72PXk46fJOw9q15me
GDE2uIlidcStr4p0wtMJgP8pq8GIN+SHDiUwupR6Iq0fZnHSt120oaW2xIJn/CFBToogYT+Y2pA2
raRUs55mUVGqFok2CfE7huLPzC2WHfIBmrl3NU6IQ6MQwspMgwt1+k36HCPmro0lvkcOIBwcrSep
UO56g2KgPExlrhIVgUXDHTBdj0DH0WulvyPcTjzjkGz4wAmgXsBzrk5lpAGY57YReStaorlWxjcY
DelND+eIH47PW+gSg6haPOBiGpN7wmio/N85uUS7wMOFs1hifBLT5Q18x/X4wxtcQEV1ZMPa6Tb1
3MIv4uUG5e1nSUlq//zkEblJC50jyjskPdtOrALFqCeOYekbjEbhBOx6lZ2IRFW4MdQtOVr3NfSr
VWyS+qBqKRZ9+6KisdVuHpW+D5jY4Q6yrjq9Z8yIf37jBbKfCA+KhusI+wKnuS3z+tLkIX98QGgu
8+XXUXN+cj53DUAhgod4x2LgKxAWldZGFrFTmwGFNAvJ/ebr0AeIRhgHb11Yguo48YTUbL5W7WgF
2HdZhXkCFlQhj1CosyOOias8dOiNdPArg6jvj7f8Cetp9+y8Ue/fSitrj80gC9W+5uC0gzJa2X+x
O5Xp2EeVWAPta5o93crhcMskwFpq5U64LYT9+S4ku6a/dBFg468Qm9ULncNU2MD+cg+L+r3rCCJz
bEgTTZLeivPMngJP8Lodyn1GVAkZ+hfAhTUxz2dD3L62IpJNRxttZMXy3ycFcfHkt9++kRnd6D9s
1VfSUoVUeiYHLTtv3q6/ZWzgzsnOlVi4mxbFjhmxpabypCCGrmeh+mpk6eMjuxS+W5nofY18iPv5
9BOsCtUa8CZkaDycXcTfJa39iRvOD11/47OngicSFWbgrKZDGHEXfDqZSwpcwraStgSGMW2axot1
NkdQdemqI2YjruvTTLFqmMHVC5a7wZSLUsDhqcGkSEEfVu73Y8u8KrrInU6f/znVMRwIGz83Y2SA
DI9w0mub6K9sFDrNaeZXnaowCFbMyulv+CjaeahSyC2Q8iuWqRg6gjtJjUI2xRTs+qNI6nsoLopX
iNM4aPzFVkMPluvaULNtBvyJM7q0fS7SdxyOG+UYoEQYCSPOoyATJh31a18sgiuLsOkRij5hSn5g
aYRnXYh7vkl+M/Y36v3WVDwlRoGxCKKxQn5P8zPm/Nf15VX+ib9npzQDf33HS3ZQwDBTZyfnS3Ca
DansBqX7Gp/VrtnTqRA8OHCKqiFPgCWZLjks4RPMeUNkzCWw+tEe6nHTUfKigktTZfY55PCkE4js
1AkY2GlkNb5vv0dBPpAFd4AOi8HeI5Dn1tqJrWTL/zuS5kRkKpDrS2fSOUYz6iLR01Owz7fTQ6Zh
Og0BrLrEdLC+jMwdcWDJY9E4mo4OdVJJGHW0cVhoRSp9CDjBjjsKyt3zvxJ0uu6uBZDgTbLhSM4M
QOURX6T+4B9XvRjZ5fTWQC7GK+j+eKjvBp7/tApP7UPwZCBZakbzLS5KMsPRC1a1+SuhpgY2ryW0
KQbzi0ifVMCLQqcYytWl1sBFTgA1BPI9KfjcXlMOlh7riKwfo6zYw/Pv0ATiQ7xX9jAt43QV3qAU
HophyFH1jlHZp3urawVe2Rg6D6MRR3v7P3aC0ovG1BMVcy9DXxHnUfoLa5uVma4HHbl7XV2jFelR
6xqV22qgkpyO3EmeDMXDGKQWtg5e7eKXcW1aD4f86q3HGjNemMzQGgUiPcx9sftwVziXcjSUqIL0
hHe6DFfvIanBzLYuDSNo9XFPlyaZ0qSBm2dH51U4RAUZl8Otd044DkUn6xI52fGMWqEtgGR0aU7p
Hqpi/37IjQ0pfHkQ4xneKSoAV147hhXY/LBGt6oOMAvm0hqvvHh4zZ0OlylMIunZtGC519SbNfwX
/7vS7m22XAHA9nlJawmA6k9+hIlQ0KhZfSm2oub+7IBDbVA/TjDfzmt3MY6bTWzHWZgQ/1qpzVsJ
+XbGFSOG+BYA9nES4aIhCtfFBqhb3NpKJR9M+xSqvDX/mA0i/dRTtsJuCv6D2FYtP6mbBhI2tjiA
UEmIQn22tula5vyYrMJbZP3ke2PPLP/QPVZNnq+1wU7/nc+RR3Zzf6A5M5ejbDE6IUqUoR7IINSK
jVIh60hzlttexeh47L8+l1six0dmzjlqJ6fU9Vtsbq3/iM4Dte6VbdaNHUHIipHOtHyZP7C3P7rr
1cFvNbeeUhQgzsKeeJRISi1KC6U8LG2VQppklQ4H1I7Tbml5L3X3TJlLPZW4MTXw4D5H5N0+Nfww
v2RtVQxGMii8uTwkRf6B3L2YF8RLk6FUfzzhqkpBy0d5qh0STlt+HHZb9dygHWMW0M0anix3RsZY
bL19L0F9T6vN0tTAMBrRc65rkcx8AwbynBboB1mPtoNPNUyj+j9Z8JrxzOSep6az3Zq6jFC4UypR
JD8cbRRj9KtCvuwdi8RT+G826Eihdk/dNjfWsqXjfzgmZScIwJmTAwXOz0Ynw5RoMtm5VmApmc2F
rvgD7bW/LrniEBic6qmRSRPMUWTMe8gANcibrjj3omYRfjpla/0QSMDWb8/8XIZOpGFtcDdsSbmj
El/cezqgYHM2gzBCn29MkaCUx/JXjSgnf3C23/fTeB5VuhtgTsUAim4nQ8gwPD75nRbocLEgUsQ5
DWlPn9zUEWZmyAWe+ORe/VuS8xG8p37YiY7lEEc4G0TOV+qpUlEEXA0v8ocSP6jLQ9dIg788CW6l
ghm/zKGXBPFaxNdvYG7XHkcFv5XTI4jQU/A4hKePSsXkAxGgPqaMA7OKCoK+PlPqYCiZ5CRimb1t
V+Ouu726BJeYJAl5palsYq9Up9XXiFDjDtHToZsV7tuyWhkMhC6Tb+7PIFa0VP6phHorRTYQtuGf
KJZD44s/Py7RnQXyhb4cZU1oo7sIQFj5/w2YSAReNyXP+JHy80zpIiE0SnqAnaNd5LLn/xwcdG7E
8IVREb3F0rBb8JQCLfwbQJPYl6m1sOFCKrBkPgPlCLZMj+actdKczKc536F4bIxUW+LAsf4k3JWb
gUZEiE12ZOAeDQ9ferOoxNb6Ev90qHpdK/p9dIYZ4OXDK9lJOKko5ouKdJ+eN3QkGlAVuh4A/xMW
fG6+C0hcgd85O0WKMp5ePxLJCExXa9HQthJwjCrynQH2q/l2Nlt8xQuYEHZMtOHXK4q5cCPajWoy
y+tmD9xHCq1EKa16owTlGMYsknPwzRU3lR2ATDGiXaRjHFoo4V19TUk13jEeqics3KN42W2hidjI
GLZlqA4BmDEU+KP9amNxvAG69x1rtCSolYkMTDLCi7ga1b4PJKve1a5VrZQURQ5C2A6/USlbT8Du
h7SIUC8s84ZGaj3VdJ71SkiY0xhoh4PXT9or3KKMJCKjVoWTjEQ7s2xv6vo/MVw6qIk0tB11yiq9
HU6x9BvWOy9JcsDkqJqwnocdJsbHvoJ/pM+/RoPA3Yexfw/JV+Gr8olHQ8asosVwvkHuGwu8+vj0
GNfQienzpnYWclwjQMZ9xdIdwO+mqz0UW77fQjLhUGiI/m/aviVBZEvLLZQ1mOQ9KGlSxM78XlXC
k53ikaWCDWC3VfYVA8Jg6QfYwHV/M+Vg8X4OoWky/gUXac2kHRFlkS5NRbwaBVXHeNCJck5AnEtv
LjVa8HHLnkKzguWWLOYGuHUh+M13aUEi8pOK+tlI5UmQLHnaAr9jlDgO+vDoieuU2tGZpq0ThfTj
qtDx3mNEFJHhS9Ox/JlFpKLuwi/8ul6i9nzSvMvvod4UzcHTK+BPIlNga7Kn5nB3DFgyv1oL7oU0
JiPmV8VmehTjN7AFRWmlhA/dmOqJNj6MFt4t+Olbe+ZzcnUT/7K/V9N3F/YBJ85NnTU2oUAvkZVz
YGB8tQa2ZBe8CCoLm0l2BI3yDKiuoZRZy10ZXt+ov/qKEh6BJlOfgRrkHZl8uLQFPyTvFaEnR74P
vvLUGv2W22Gxe9VHhAyTcJtLCcRZiKioY04jx7LiHxz+3HaRrKck+/BLDkCEDBw+QLxntos33YD2
XqIWvWb9uuJLPzyEjkZ/is4QiGY8Y63ZO/1Ei0jjjuvHALmz0yLlHfInoKB5AGbt/7xR1Pcst5wQ
55iqyZ1K3lVDrz4COneOUSEHrfT7kQVW7QwA7rI5jY2l813gP+/yk8QaZBsuItLq7/bbq05oZiMo
/3O1zd0mDBSCC1lEZ1HBPRmV5C5dIZ1KUKijjn+xsWPLnR1LqPn9ZhRH15cBCrFkeFGGBnNmvKX1
vbI8ZcVQPWnxdMYBHcD99gu5QvT0rcG5kUB96ZkwmZ/RwxDY9ZQwdK29LyyFdCcUZSZ2q3Nwm9fY
vs53G13rN+AVpC+0PYKvooe6pXZIygb50aevN7K8MF6mjcyRyteNkQ6bMJM2W3dDV9G6E9d3wdTr
F6bKOxlMhgbvDStUTfz9McsAAFl3ZMGgYgIK+nBTVA1nxDstysA/B+GvcCykvt8KjvkmkQOp+Wfc
7GbpqkZGcQSPFpv2KEFCiFoIMFEpoNxaIV8h1PoLCTXwqaecmyZtOjNJAmPwOCM+44XlvGlhoYRn
tAdDhGlfOQOqWHvJTou3UsWX1hNhYsrW8XZTLYU3y2mTW3ZJR6p+909VGYE2kzxm+l/22bYvzq2N
a/Ejk0KnV/Cxk6/J/iNNDpP4RfUepOTeVJYOYiuxlewnwKudP3Kc1mI/rfBCqhxEUg8CujCXr0RN
fvKvecpinUaVsfH7cxd2Tr8DRXEkwyvf5vFxCSClcYoRhOsb7l7owAHv8UUS8HvH106GCkeEvF4H
rZQKFV154Wi/cUnsgt9gNFmhWxOURMlvIkTOFaBvpLEhmpWbd6hpKinfCT1dyhKcaBki6TvSZxYd
CdSwTc6UwoLQJ2IbAwEyIkiH+AJYajdu/y+0ymff8i2l3qelh+QLUioQAHOJQrICGAqqpLHmEwJY
iGNOxCWwz4dtUyBR7+LPI0A0x2JlA8rlds4gL6FGP8NXfjamMgHkqVcZboLegSChroW1yDTbuABw
sALBvtXue1cUJE9wa/ua0GjOo21OUqK/CDsCaliXodY/ZCcKqnTiuBYfJJDsg1ajVS1xEeubVaTP
WMSSgrVoB+oWp8tspQ8Jvw1mhTdmQpd3sr7YdQdrmeshlZabQ8gmLZDTmO/mj4EQsCffSmLC7Rfv
3Usfn/UH8Z6Zw1aaoQlYv4r3KMKMQDUPfJNLaRB5eJJMhzmwn/yQy15YN9p2BXXO6+tukOnrPKcd
6zmx5l43VXFZEbS1XUxXYFCjuvsMFJGfT+Ctte8N+aeESs0G3NEkYt73JYtazH3RUR9ko80RdBbo
bQbSH3EmJmSrDsu/dM63z9roMevgLTaga1gCNJFqQwkS3UO5u6AGCZ9VMcSsHcnXvsQDXw7ZwKKO
pywPKJk9jjx8NB6WNGabEY/ZkVW2LPJVRfrb6iu4ZFmkFNBLXaMSVEl1jWUm/8RJZl5Jlkbo/vPI
PA7NDrs2Jvd21DPpeHTtGTfytV6t5ZyiRWZXFLlESY7w6/M/RUYJCKVIU+iK5IEu8QODFzapZgKl
8pUhCzVbRN55meJO4JNpMFmQemTs7vIhbK2ohOqxF15udasHJPQzxtTh8Z9Cyg8g5X9NGeqr3BZM
+ZgwUdyGr1Mcg765Lo3Xt9LZ/OJE9iA8264uTrSsAEQZgR4pImZ9cpSNK8B1jXBmLaInW5OE6nLl
enE5bhJt2Fw67lamMmNbb5BBwgkiD6kvpHihYS4xXE4ArrPaJ4zO4V/vSKZkC1eqr63dBwnp1fXB
dqBKez5pLuEB1Ymv4ZWHV4FHtV7EubRqwnTa7eON+08kdBPFa0sswmqM39VkdupPGhCrebIbvmJ8
w/XhAFXHC4pOSz0fxki20nbgb2BllVscbNdyn4KoSw8AD+cm/VTWgpQNWxdEZg7ZGkDexjdkoHcO
bMCG6EAydcaRs1iH1nEUMiKlsY8bxbtdTUYoRwogsjIYOidjGWOSPQS5gGc22Lc51YPqtXhveFSW
d8C5n2Sck/tmlMFtWous0/dil0bgpGMDhDmI5qbGkpgwCbwzrXXxYk6TKH5zvS9LAjLbS/IV7RyJ
xgX8EYH9W111mj/xov8FSJtLNQ+KYa7MiE/mpDAp2ZHlQ+u0Ezny5JlLOSeaDrAEOsOUnSgmRryx
hcVBGpdYsG/UJHTbKeBUwCtGm+rK3l+CBsJfPcQo3uZULtrqQY04rf8PEnfDTIaYWZHyk3baSJOU
GyZuN2R+YSHmcpgSAu0oFjyv6aNX6Q5jV7z04kszoH+toaZoz8xYDuLaP9Lsz44xX3m6bV9IYkNK
cct5Bk1nP1N4j56e+jzhpqWqM+z5Go8C7GpHFzZgj1/RP/pjTUwITVjveBdfVGeSSh2U5239bTfP
VYA0zXGSOpiMH+N4PS4y7b0C5V9PLxbiQUxoomtOU7Tn3nbmvP/RXrnVWZUxoqnQ88q0XlkgVZ9n
97++5noomcBQncOyEFEJoxWKjGZoIWiAtsyGfBbwx5vkEZ7aolpwQLDjA7scVQVufI/3RFOGMNHp
P8FSZtWCx+zv3TAiCSwKGtvn8sPzIQqrBDjaAQ3/UjrzvG6AmoIMFNNxk6Z95GgGDc6REMrDUvwE
Z2F+qe0lJD1U3uxHrKbhquBVe8fqnzZxjyot95Dd/RARtwIltVkUYnxWegG+nw0CzmOiVQuX+xzn
/l622CT98Iu9PdTGioYcJ0kMukOuvLxCQWbdZ08Q9wCpNkKbnHz56Ajt6xAW3VfZgBa/7wXvERIw
tcufd8+ol1AAMxY+SoOXQArDzZ+YcRyoUZSL9o9jV0DYaun3VtTwZ4RSbg5EKUf++LM2u3MZZqAx
9+taIycLUxBi17k1Xg7QIbIXdWPdT1wcSl968XgIUQHJFX2KPB+27JiY0CH0d+HFgDFQ5X16EcAW
TChuYwFQAqtr5w5P1o4rX8kh/9bCynC9GpUyKXENdhFxY7rqFVhvhumj0xY9n3RO4sqN99pG01WL
qUGqAhIXMIznmM7kPvE3wVXvsgXVB38rnBV6y4Ze+Aome+3WVGbIKi/61Z8wOrzyWojw6qV7pe7b
mEBNLuHTDpq7mw+fe9xojjVvvSPNdlTnd5ota/cZA6qwKM/G10q95do5S4znMsjzJ3Gl9gJCMRbc
xuMOOKkR86E7e6+JiNrp6vJ5NtW04u5IQgxRZivsrnwIypmhagAbhZFwG6aMyJgcaFGwv9UdBJz+
MHEOPB5XnIV1MpRJK/hm/RrUAtByION8mqesO0jJpI0BahDPU/uoD+DuQLJnfDEN53ZgNcbKE3Eg
Rhy7JJKSq5evmR6clghjBOC2v3J5dlYZ6WYq/RKtTQ1fXmgv9uSgnVqDHyr3ED15POou7tcnq3MJ
OUJHID2q0YRWUUVhtdfL4/loNxC8PjAYUFj+PAxbhLsQyd5g6gD2w9+5PiYJt8YZxmACIuQFfR3K
9DO9oIY+ZjpC75D97r2sO68MWGHi0KfBK2pQyLcjZL4hn3EP9hPRnp3+NfrkAjC/YqRgb/XwQLF+
WQ06ai/lEkl+CwtPLgNBRYDhWIjFxtbFgjCnWaHHm0+/OM6I8yBG2+wvIFpBLARF/8bdhYVmRGhr
opJ46KhbvfjFOdKa5RPJ0936QTZ8f4s3LguJM4fJIe80inF2BxjDb3zaiNDpczxx3kCTWdZdlWQe
ZyKxwMKZtYPOKjQ1jViUOHJhL5tsyR6B0lZiBJQ66MTBBIE0uMOVCuFPlAdov3xS10oFQxlIapzw
esMjJDnYxtcYhhV1QaVuFAAQqkwNhkAslY4SaGsW2BR6wKTLvzH5SSM7n187EEUppeW7m7CnvkNM
Yqnc7Bal+PQxIq+0oq/Fu+5WVr8TE7nvKV/CxvWwNSQA7G0f4mTm/njAE/4OvKU/NVHT47fRcgal
+0XR0SauXkNL5uLuJo1vYlHYXLc9LxvMD2CN+QRgyz8teChBPOWVitXADWzN0xKyLQxtjUaxnkg0
FgIfbKROiSnylKptZNo6MBOdza805q7hTac69S/HsPaFslINMCDVDBn42lqwnallmHsl23F5NYXv
KtZmZ2nQLeoyls8PCB+Antmf0PC0fLbSK6i3292uyB4Ge63oABlpsjiH+aTYicKfCe/kH2G7R0UF
P3qBlg7ZIUgrOUQzQHIwK+uRip5bmR/wg56pb3jy9iYouXPFQwfGZfqIU2QiPC4sZeMA23cAgRg4
aNFsLEx/kwTduqpgsIprt7ANP7z2b9YsVv+mmkHM/7hIucB1lBtT9T7Hs8slpG/wpmoPfQgr3dNm
sPsm/dYPye/iJY+zMqKRPmwKX35eLBjVWe9ig9u0NVItu/4xbaIyaq1VUL44739OoVQbg354UKEx
9oLe6Oz0RmH/DP9yebWykx7k83YkIyLUUNnaoNkc2sc0KywC7kExEbho+Epon0LYgOL4FT4wPPdR
HSr1wo3xirpP555/+acQS7WhjYeEvmbqndv0HUamm4yRM3z0Bb/CdexNiTVJHMXp5RKS5hC1bnGy
5chTZYyaKx8v8dqnHUzXqrDKz082EV7AMrb4OPcF5KEEs1bo6d4GOxhHjiWtBw48stxmdfG7/aUS
yt53vM1trdRRYhMpqGxY+uHC9Mhy4ObxzxftzgYemk35tvcatIfqLWQ6kl/wU+iBVewtWGkjDLVH
QraUx7fR4hE8GcIljDiFCB9m68yeUzORUpzfzGuEsW1ZuQHRb7brweaOrKcfhZ/IL7n1ZXK+Dcp1
EJy5N1ZOBKeOFuvhmXIv2/rJtGHrWHMPCGPjdfywE/5oLffRh5gUaCrTirdU3CSzDHUUcJWf7v/Y
+b8ZpCM/lhQ4zjrwroPJ4XJ5+X4oInE3we9jmmme2oow0CpbGcA6vour2t/OCn9AmiXmc6rnVUZg
ONSM56KZt0dlVpBACdzLvcR/lt+L48CjPmBuDhuAqAM4c1j3lm0+WYttswupFIPGLVRrDA85ZKJP
C+wN47Rn+UALtLvf4xtqesCX6MnsbJcGRAlL19uXBJ4vb0OhIsvDMUKulaHuvXV2ahwte3MdY8TC
P3aGFCMjcg7QIjzEJDBKG5LDQLbtjb441D0Uptz3Q7wRQbbxd8TBsstY2Y0XaqWzO4p0zJFrXW9F
7aeBpuL9ZIn7rmYgkNKLTHRPuh8v/YBD3cgFRZmKdP85iyYwkwvA6x0ymfn0GR/6y/Bw52e6+4IH
RfSX7cQGL2GomwcSguVFHw+VROlWC5p/+aX1YGUJIxzUBKQbj7kQdw8RGpZ6PMwcdnLLznQgMoRE
qQ7grP99FslI9YgR2icJ0mikiGcofqICtry1mmlmSp6PB9W8keGNf0xhFnBxU0VVP7qW6MOhnR5E
Ae5WMN9ZTu5gqL1KMA9nvdFBonIX4tV39FVLyLoV6Ac/FrIb2WvzcuJCo0D/fPIOrEfVRZ7Y9WYZ
zWGOhQv8r60YDJNTkpSIX48DcOJcyEGEXLNOc+oVz2RPYHwIBN6jhtietbrAqBC2Q9TL6giSAbMf
1E42vCPT0hOIGId5iw08uXY+rDR5hO4Pe90Li9SiEm8DNcoDTMyEiQwLPi9WY6g/wA7mZ5tSjw2d
SVFc+RB8g4m5bRSnp9SPvq8Y7HR/bq+dzw8io5wNjEACT+rpX+E7uC1d04bSaVlR5YTHUasTOfCb
nRjgeSxqAh/66N2xmrYkdx/T8QNyaTzMK0Rm8rVBk/KfqmqgZ9Eu5RoRfOI3Ck0NDya9qR8/L9Je
muBf5FOc3+DS9SfkBBsAO7F8fuPTDivlYSL0Dixls5gMttYl4OB30cun9KxaNr9vjD98zsinwZCf
ItOrxzOWgNgGjwBzRPMwR4OXLngknsrqSqMPF+lPPuUI4lTYGx2XCogeGOaTWuNsutmbvg3YDocO
teGsHg8PzP5bQN0d+0J0qNpHGYei5KwdPyUtFc+pLyV44OC3wZTHvmKINKxRzgCTPy6g8LKDhI2p
ELcs4HE8EzW9KgaPO8ew/Myx3sp2vv5lH7nh7DNPeCIsKgM5cmTOVRKWaGh2+AKGwy35X5kDS8zX
UwQYICcG1Ab8gVOjGNNP6S5VEwn142l9zVOEuK/Aa3CBiUMDwPXMavWH8M+ldRZOyU4XFAlYKTeA
04yatAAHyrkRWFh8oyYk1SqSZFvjL7aRqitn6AgFi8gDjk6FPb6momaeUWyGoic0jdnK+5xZu5kP
H4Dk5ayBWoXRsJulZ4ijGa54std/wTFkNaW236ZfcaFiHh2aHuNIumyJ+YQumhUU9I/2tWfymVgi
DYOXGLa9/7cK0FwcA7YuyDQO/6fi9zBcJhqy+TPbNlJrFbSf8kiqCguD4pGo3oWb3C9kQkM5Tno0
itoqVVmW0uCrFuW25d7tKEb4zCjnI4jQskgkeOEXL1KlQPrmQUUOir/vlJUQCrI6mfSQCvaeaVGz
jdcogYqV0KLZfV8TygrqdRMWb7ZfUQ/fvCSEFJhRW5N5Ze3cndS3/bkw5BvbH76l1Kaa8PnYnV53
ARCOGpYC0NmMNqLTDYH66rWnslH7NCHBaXpIq7KrwiLwlepeEMgdBj1t6xC9EbKLwdz98VKWqorW
mUQd6vNDWNGcR4OpFVRyhutI7heVzM62zAg9Go3ysWsI/Lal4Z6UFzK5bcBLxQCLvAIKmiEqoUGc
Sq42Yq6GYQpDfbmBYHocEr9AiVG/WCecfbN8vEOlCOB2nvzSQi5ezmVXj/ifvYlZaGg0ATEOfZuz
EfghpFSAZw4EekGxbFA5c42r/+UayAnTEk8UVGxQoz2SbCXgk9OERnUbhnyt031YXKctJAY/czaF
j8rwdnbgrNCM60LZtdBhC3Mdoiojl08yvuu4jKGROdkIilCwEonS/g6HvFI9F5NevBECjp6XghnF
JN5F9+1AHVFY5wxW3xugML5edQwH/N6CX84yNOeTaolpDsN7Grd2Nxq3MKgy56rUYoRPrFA7PDD7
Te+Ey5JpRXDRYVn+C9TEEnv+UE0i/EuXtvtQbmFNptedC82akxD2oWkEV7JB+mj2foYXuQQ13He9
0G1r0OBdGJlwfaZqgtbzATyGiB5DJ9nkxZnD+KmhJdZve7eWsgBYFxwp7nAdiaq+oGnxByxgjTEl
CMi+wum12aA04W/xNyAc6rU5cyJqnOhBqnOkdDD0vsVpoKs3sdjx4SULmlX6xebNJTztAT7NgaFF
J71qj0oIZwGxoGhFsKWoGzuhm3oQ//RgAcdUAtMwYbuSvo/UFwKrC7Z7ZOFW9FZOvfMj+yCXtf46
OzRMbtOqbkcWWK/xz/PtoXW1PmgUBvmengWU9SlJN4xcTp4hFssNu1rlyO3MU1YSyfQOJk7ZKX8R
omOBWphTn8i5L0qDAs9OSEhm5dX2e92m3Z8leW+J6OAHUtzQ+pS9Hk/9UyxzKQUEq818lEPbrKib
f1BvwbY63uq3zrhuYXg7Hf4puB4bOGu+ckcgk/rSsCA+YKV7gG+j06CDWPwmbKhcGjdU7gQAOdVi
kC80C/HU0SBhc0p4fkMBsu1aHUXeUUEHm3ao5WqSEnTJLOu4//ESkHoDfP3gnYy9yklnM90anInX
+6jOMSAjsgugjVRjjgcaBGqjYutpMvuPjsuwsl1POiOKmJAAMTGHsyPatxKiFcjE6biY8hdFos1m
gMEr4QfhDFwfzBkRahdC2ydjt4MmMiw60CVU8QycSuVYc8yw1F5aQRNBQj4lpg2pPMlRKCk/mu9Z
oX31wcml8PMSk2YB7Pi5p6lLA2Le6G8QhKj/H285j33n4sL26UTDPjWqsXBTZlT2eFcNsLkQTI4V
OXXEg9NluyzFnKxgTZxB28B6zOuPDzmDL93NyPW+xLNybfJ0NxMZ7355p5jxDoBnlBWtxe83aiCs
p7ZI/rcSO0rfpfiBZvup1rfYu9okwOqIQ01+E/Lh3+B7TlJmi0GtlJSrIC7oTIv8tFUDD4jL1ErI
qRD2eM+6n8VwVBYz7ZH2sOke/xsOkjmmNIaq8omU9AUF483NIX17mtaH7BMYwHSeWr6HGwiNwiSb
cFVnLB6vYf+nRWmjDN+kcVHQ7LTyi2tnGgIn4XG55snfeV8Y3yi5Eu5FqM/6dcA8gjzW/yA+9/wO
QHKq1Ahn3AssbGUNscFn+Dx54211afpCAxtERK1o52eQwUSYIvXlNlVaxM7i1kEz5byIYj7jjeas
DiLl9DC4+Cz9XczffPpQIOZ1VSgOgWMC3fATAD+0ht615gcpFDw++RqDpZ2aCMIyOcpcgw8+CZ64
7bcNdBBjL0+BztfNRYeppq/+MUfZToid4KBzyXXHxcb8t6/dj6MaFCnjAipuGvsJYJckKtQC11qp
lv5NVeRT7cqpkxfOLjn67dDN5ebiaOOyjAgR/9MocT+GEkt76hUZ8BRUQT0id8T5pvnUo9w9OeTW
DUVnrL2bCto9kF51d8JpRG/DpNw4UCS1qEGlIutPCSGqn5GdjvYHqNUlaptOjNErWWcrfudVOy8a
plmGIwsEEBXoRN2EecBQheP4EH5gv5c5img+WNnRKBMyNn/QeYDM0wMaVMnlrDtMYZADktkqLnza
4EQmtAI/AA/ygVI6yEL3WBvyCww2Bn19+Vm2+vSeXOKdyhKZRlTI8m5JrfuBjLcnYzJrNdLQ2d1n
jgC86Twu7FFOXLnZbuMV1s3YEw9tv4i4hNNX2bwYxHcFcZyFzx53ArWTOE5q0+Eie4xUeHDXaO+6
ml7+1JryW1zhaiY9RDsl1rjTvjuUs/WVHFY5TYtZKWHkSb/afvjCyjW6yhqZFAsu1/pUN7dCFoKp
X03wlw0CKQKd4BiBcTfgnBPmRTSl/ahx92c70LYUvAQ78BbzKdGIXV0ybElEQv6TgLsul/XWUpwC
nBUS+mH9uK8D4qWLHUm6XDlzSH4MIl6D845vB56Qh1wvY4OfCQH3upR8CptV87glCDbhKiYn8vB7
fO7m8cb4XZ5mCyXq+tri83sbfzWjNSBQKw143q/jt5qcsqIcNOmOoCzPHQeabgkG9yujIMWLUW9G
r+ud2fnfR44n18Sbp16ur/RBA+uxhDgvWIovdgNQ0pwcFbCnbTURy8ItjGTMNpsAe7HZ/24aZNCt
GnixffznjdPoBrLLXf0EdTEmBzGgB/SGWm38WKdP6eX4ph7dfgqoqI++Q9v6tLscWZB/nwhBbDtu
oDAUDoSAw4s/aqpH6nPpuiEtl7pubvOof4NnhJLla2233WMyvmiCXD5prAaeSMKRItDmKBet2uI4
LTOJ2mEL+OGGYmHmrAKbNSQfv3xBAIaOL6IxITX9p5vB3tcqkICGYYS0DXtOrEq28vT8Lv51ySbU
BAicJxmrVqRPvCtAcEhulcy+f1NHyUWdkRTSWv5Po3CJJ26Qlu+W/vQNJnh9BOW84rivtkKhyTPx
5ueiZjpnFS64kxZZ3AkQIsBHZlsCfuh5n3gmJ0AMm0DydM/NimyeI7zXJ7pXx3kDSaIJlhR3fdkS
E2gmU7iyK+un55XgM3auPP45bvhYwv9Wvae9s46fFnlcesCEIlwVDkPRtJJPzEfbM5VT2pZp8JtY
VkxPgUf2UjRVKeU/zDM10JHFjA13EXhQUUiA7ZqOKw5gYuGiegvM8//kCw+WlH4qPN2+q8ESSxpk
q04djI+ZlWzzZR9uT6flwPT7+bMMgMMNw44Jp9k9gq8RCzpKP2lXWycuTvibOI9Qq3lIKNo9zdBX
mu+lRqBcxsy5J3JxwWIL593NJ9lldwx6ZYh3v478T3zsdTK8GT3YyOInBHfOCvuKOaRxJxTBukSd
FUT89LT8kLN15UxH93qMLz41Or2MRaX05ZUrnygxK5oGTSn0hdTiDdCk0nFWN8Pomo9qg7UJvzWs
+WvCj/DXn9EDuJxqNVWcMGZ0PuiIGdIEgh4PRre85u++D9nGtJab1fFkDHpmUU4P2xaApoKe7daH
5hF579gQaBmMP54pnvNwsi+mbBRqv8N7RAToGYGLxb5O/y72ga5cGSNDFUU7Ks2Qlxv7Soz8vYX0
z/h2YL+DVTLqOPUG2OAN1uQheQOEfj3noLBXBi8LBjZYHBYdpcTYtEnUhg0TpNYHXhI91UAQLlNH
1hyF4mnMge3hyf73HH2j/Gax5dE6xFXcwidhmQgrg40qtmFxbIpEWAm9XatIYVMGF25EkZJqGwGu
El9d/ZlsN7A/QBKh4+MJjqmD1zkFv+L5XFreXccJ9khhUa4D07Zi51Kn9pJ0Yhwx0S2CjmOAaMQW
QfzaxDy4eKv/RTkeEquOOEYtrAY6/q95bYav/Rf2OrwLPQhiBi+ATkxxy1QCZSugKudrL5CPCH/6
OSasEBA3sZ4qgpbLg40zE+A7oP4OKPCwNnSVYn+oFknMYBYEM8XlFU1k8jNa4PUX2nGJRANXkLOg
96fjjUGCLs2alkgdxLwWPi7tX9WAmmwJXEHp4HTOq4mkQsrudn4KbuJBQ3t6wMHiF2LGm3cyI7eg
0mSq2EX0vxVGgospVSzNamd7a7l9/yAmLdOcyq5As2XI05As5mUD7X4/XTsS+ThDONQLMJrV3Hp5
EIVihr/tyVul3liXUg81/DCQ+Bokfq4tbR8DKfLHuWb1rffbMTE3QFkykN69IlNaw1kPQ/sIqKxH
0QEXM0eg7O7H5Nag7lvYr8/HxVrNp4HIF1W42dTVXE9WPabH+FB6Zpqw1Lo/FYyFqzFf4ubTpVrk
7Jw1Haz/arHz55HyOH3TnomLLMWMU0RTHwYcCxjHkutIVJfYeGkI3IS7OSWJmzIgcX+vHhPlPEtb
mdOBWd/mykM2JyMyrBdpj4zBmAZNINhD0lfJQccgGFWH3BGd39Lrue++ZeC6RNW5Wc8q8tRrzBJ2
Ew4abCCqbbLbaj1ViNtiylvv7QoBEL0U8gCZK1q9N5RJpk0JnwLJ2HrLukfp70iP4Td2/n8Y40WM
40uRgDGftkq4Prm0/Ryo8OguWyuy7EKVBsKZMv4wNY+wwQekEj9U0Z+qZX0Qa9wYg6MVf7uCvL63
/xL7fUuH1sGBNYf0rhQXXo/JUOu5JSgrB7BLn2dHRoD5EHX9fjWKrJb7LSj55vkCmw1kNpRR8W+z
Aa1jj+l+kyAysxO1ctD/5Y/2F1R7YziKU0jDWMyuOfDjJ0Hj54NH7wJYjKAL1HkB7OTfDbr3MtJ/
Kaz9pdgyJWTD+d7aVCRtunudyjTiMnoNKGR8G4f4TcFh3PrbxSLsmY6dQDX7RcsK4nadkx5XssRc
TK1IknGyrxaJ8Q7YSxTR7RSYPZGujdT1D8C0ujFfIucbFij/reMhf0zQPcWDnuIkhVFdPrwTenRt
p4NMD6nytWq+btJ9mrxSeDtIJkdETy1qgsy1+K7+SGz5kWbuNVODwdO+VMYF8RH0t3Pe+M0Vym1N
u1dZhcXuwCCcO9DaG7zW4a/04uX+aQPT9G1V42fme9xaJWKgaVCwEJz9f76GoYdYf7csW0HktkkW
8kbA8i+GLc3FIBHxTQb2a5xdcCvgzZrYr8DWFCjXiVwOdCANjMTOCwqbf8yOl1vsBZMf1F4dmpsR
SgNNBpI6a4WdfSNQvF3k/+lOU33nx8b/Xv8lCUYPL08zDRuMkn81vTDqcpHowZmllg7Eb7WJM7LO
apYmWjxYsSsXxlIEyczo09pwwjXNuV+4tG+OGoaoUV767yQNi1Hi2qEO0A5UksR2vbJvZqGxizU6
5dKtK5sJbH/CfbrKQ4UAIvH6+yEnKlKNhdbtd5EdRvTN+9I83xvB1V37nAZNYV3OnzY57NipXX17
hpEjyQBScLiqDEpnco2H41CT15u4Jqv2VwGaqEMsR42O9+Kb7wluC/I+EO0dgdwma99U61nOH9cI
NP7nvM0oiSAtXEgQzcb/WCwG0Hd/I54vNgsA7dZjRPA+95OXJ1snfal1rE+IgcK5LdKAI7RFXM3f
4nQO43/Xgfy1N78EmMPUfeaNuejlQ4tV0s6UTAOWa9tALbL8vNGQoxQcZpHPUeZyntkuwE+9HSsq
iiWj1HrOZerfuc8z2PncQYPxYINXY5PYxcclRiuZ9lzGJtAcrWiXWVfPJlrwDjrzvCXqQvbcD6f4
RODKZHvtf9SqrgxWQrdCm3bcjw9xhY5gboGYhFY53RdF782bTJ6Hu//F4aFipUj98ltDlgWdhwdc
F2RGsXKC2rSusDT1tJdztaF/cPx73pO2Sk2KRyznFts5ShZUNmuHMRGg60qbnu34V+Yke2NRtAWl
yApcvVHuuVu78550x/DFPM8Y0k7P3wPzSmHT4sT0oEZQWQkTLBGJjsDNTfT1HAeJKINXfUS8aexy
nwkQJ4lJ83A2oASVzyPbXRH40Twvs42VeBjO49jOVCEJui1jiOjY8VJmSfRKU1i3RfBN6s7a8+gd
pIdX/h2k4C1Bx4phNNivF1VasP2NjDb1bl39RzUZSvuFMgQtK8N16FU54lJnK98pkbpq6NPHgcJG
MhY+xi7DChtFoSn/KaWppbiYbKpwwK0RtxCr84xj1J/mNR5926EKL9Rr4RBE5JOVFW9rgTAV2eJC
mgqwTE+SLwtDNtDoIaPuvg46HmVemTk5s2F4WMcJewf7HPltRv4KPfQSMrgZXrI6sOlfoKuZ+HFN
FrDx434nk0NTdX59KJM9BN0WVuJKFESIWGnNmRL44ArKe4zF3tp8kM/gLPvP7KSI5HyvPNOiHSC0
4LyjdkqbDEUfPCAOgT8Jlj11KAGoKF/v3igIsvGDIHsPzoDdLxtlylTjAhzQbsFQ5wNq3nTDwzon
dJ7uVEFlycBdtMwkJJTYu3+3tCv7tLN6CgicYdtNlxfyW9XJTNiPpvnXUh8f3olnEicYxa9KrRCc
8r+FwstWfI91X3yDOt8+be+sBLX3WNMdI2UFe46BJ4j52rDoEmgKtE/ZjxFcEjRZzpAzk3/4sJpg
mVxoX+E35mdgeXrZTgTNJe7a0E2/gw77+cGgf8qRxfFn+OqIOvpQ5lsHWU/DImQZ/iLN+nk7H1YB
saKeSpjrhbKx1yRuLluMNCYslvsmhyt/CFft14DcfK6NbKNP6KMhKTW1BiFXsZMgIvrS6hTIb/hl
IgxsPyCKlfOt8UTAGeLd7eh48G4QFzZ3RjXrT8NmLF0SALSl2sMAzXDlBY92f+9YaIqO3HInDaKe
54WXuCMnBYkb3C5zKZ2E48k5p7MDhwvxG/jyw6V6DHO5Ao/gjqRbnKmvB7OuWzAJLYKDFuC6HuWK
O/OoAV9su/SGkYRj2Zoy5Hwzsvtluy3xEOYENzpF2jEJ9aBdJEUDwjHS4UJmtviGvAza4uNyWpA5
mlvrTgMrxfb71uxQcxYLZnKXUKoS+MKkfnNbBpZ4jFkAVJDsycN1QspdVhekJaIk2fqDtnvS+Qph
Bhh7b87V6HS8A+ZrkotfVwJudq3fkZ1EJvveK+oTcSvgwkhxH77gmrnFUiPrEsZGj5wGp9WWdMyb
2eHRujICw/RkHkA6BoT0XRwWeBIT1CzpgKDGZVWoOSogMIY1m8xjzzNemE0qy2jH8t5e102DOpsZ
fliibEL7/RqfOO1wwQFfjpCHLt/im0S8DTGE+Pfk5T0aK86xy0jCqmW2BgQHYyIXIrHUW2w0ac7y
L7bKgYvH/jwAMr2kUNxmSPIG8SSWQq1IOOuwK/hRHxifOvUtZoM5AZ/XsHuZEDd5KBdTOg6GpxBU
g40YlZxRpvxvj8w2UzCE95v4in3zyJdZJYSFO0+lqgplnAGzbFYRxDeFdsVBwdcfS6q8dWnsfSRq
tf1nueoh0s84/4JmmIw6+CE5mFwcdPpTKLxD0KHDnsQ4C/tuZqy4URIvelWugPMHZigREXLAuNTj
Zq0pRxb2mEDBYklwISgZcFcLsb3bK75zoAETKEssP1GHW2DobFJueA4/uVVjSMCUgJkaN6TTgCGq
n7nR+qwDZzjai2ESRyQ+vD7P6+vIPTPYVXASwv3vwG329oTHOIJ6r5hj7LAKy7rmMshhdXBBHZ24
a1sX6TBbuCyKJApn7MEP97h5A7PzuCm8+Y9fwRU0HSi52zZIQYSlXuPbJExSnecxBnLL5J7vGlqT
O8eWXXwuduBwm4DWcBnvD4rX2b2w4fVqwy7CghpieZu9l21uYdEncJJnh1eozjRrUNmvWPxp3WuN
ziXeFpi6IwmX/98keoQnrhQIX2UoLsqhdbBuyntw/mTSIHNBAnTjb9CVG60JCDY0/H7NZJ39gSan
APwrLoYVmbnTMIhjwUPkKoAMw3GFvTeTwpFsBMz0LsSkqM7a93aG4doJ9dCroRrx+7Kn1Zqu8BN0
sXKq9eBDkV2N2n1SBxSSiZvErluxTDj6g3rS3xo8RaQ5Gmj73Ypdyhvwo/b3uDOhcdOchz4KwKBg
EzfwvJnMISD0mezQFmkcePN83vuSfnzGzIuB23fMKv99XN54YHrbEG+3e1F5q3wWAGsMohLTwDfU
zBLbPAUiWb7Awcid1B0XA5ICfbMhGAjXukaqK2Jr7NDHe0IW0JiihlArZ5oSUyDKze39gjmkwLSl
fs8puJez5tcmuAD7YhYnFTXt/IPHPDQK83aW6amQxPetLsnixRl/5ojuc9sRxCLXFqxVDBAznTZX
A4V8ZcRX3hNObGNDtrIVdpEKAETYyDmOXLQTFsqr4gb8OI2/WDQNNqrnukKCqEhKS9kSJe4H9T8s
vHLqZKhVK78qUGZOCnG8rCZm7GbLtsFhNB/fzPzK/EJzNyn8L1wDuFjw46sxd2U8mTTcpo0ejOwZ
mu04wZosmdP71yll5kUpWfWG7uczV1651e8lExyZlqiz4RGeYNO2GaCqpAhvG8Tsnjxxu/MWqpa4
gjkHSKl8rTa/rMiGMKvnls7K/6PyrOfa3Q7iRVNHe++KmrnxISIUfJkc2pzwFUFyYsGTgTFfot9E
ofaW/W6jaefrRp5MGrAZggqKhT4Uy7yXriz3a3Meu+q7GXUTv/cq5Pi45Jrytaxc0KYGAGgfNhTt
E0H7qO0SNLzOYJlKCugbLO2VkX/QG8/iumOG5SxziISvvTQpSe2etpxmYw8TpVuAOkQWcqJwORtC
ovnvcPNolIJDC6p+bxau/hKXawanPYq+U3i8wbYhfCSgP+eHvt6gpY3JRn0aHuD4lFbq8R//+/TN
lX9an0o/wrl2Y/MclhAryO+vjJecnE8EE1VrWMYmPpv3/wjjKizLjN+evTf/e5CXQDm8jPtHSE3Y
qeA4FVYCGb6OJEYzvHSzb45iMM8/TrMQlklm23oIF0Dc+2sQYa9m8XrqMzOIOogDn6gGTHdndX6h
gsrduahSQW9JdWa1eZNLXR6B96kcY1a0v6GBD/suv400eK3FwUYuXS+xEobsVP9mbRbISqE0Xmhf
voU/nKR+RFe1+++x5bWuzo/EnRBPnwcYzU2l0vqPc7h7Lt7PT5qu+lhAa+yi+6Y6qHxQGVcZ4gBZ
J6/AYlFwm2tdxPloOI+SSoYvzUo6Yu/6VXtBw7JuPOGOUOX/Ng8WBCzRznjxFHAydvwV0eNK6axk
gPF55nqi7OVgdDMLRzaP7w6PwVmQlhAnHQn6lF/8AeTX04/AWuaDTirmlIBJxgexSySiqmCKdvq7
zJP5TYXsrGSnC4sMV292prd1RM+D9r+nGoZRk6ortFWCnSDnodBpfgQ8MZ87rpgd8u0kwSOj9VId
OMMzvhN8HRpcgakWLNoo/n5ud5hJ018DGQd4ROwRxwg7cBcpnCEKWMo3prAaMBML3axYvmFXVd9D
yUE4pKLmBhv4EtiQ8cBTgdAsjOOZs8jr8P9co4j+/2F/5znU+l/W/+hI2/929PSSOcYitdT7vCqI
4DTY/1hT/T3LYuHuQI4ngjKMoLRhHS7JuFUC90P0Qv00bj9bTj5mGlK5oRKqXbfJswAV3NXcO8lg
mEdMTT3RChfQbPu7aBsKxcOswzHJu4pf/BiDanK46gj8W3zJWebMGNVWVkDCEi4vXhlzB7ZDYR7s
TmDY30z8J5TFzYBRgfEIDKg1Rk/fMX/SJ4xQXapNGb775DOxJJC9p0xOwk5FhlXZHVQuP4+ijd0J
saGmc9Qrrm1GCckqSiVdSMQyNwcFedgDBPaSMJDlXQH7/5WFVyZ8ylzMX6zEzzEnetM3kDyd1V4E
HGtzilJzbZi6J9q3QsyPZ5/AeQFRycJyah+TsN8bvSjYdOaYBX3z5XCUKfzH6TaxiZpuNRWKfhqt
LJx2Wja81wKcM8qrMFLacpmuMIXtSFF7ifqoGlaBVt8Vn5nOKWbb5IqicIHgOFxr/esGwsR6mYwS
5SBmDHEG9vbopz6DwNJjP7scHesxmByXvMslMPO+WIHLmZmfiTJRAoB42I5fTNpfDVRJjXDkkFX1
Bp5ySE1pYLRNAOUnTiNlPXt7/N3596ejDreJK46Pywb0MYTCb0/iQroT4nDvkE+vanF4XS1DKYun
OJSQ9dzE4Q9mOj7j4Kh1pxFM9JYvOkTPnhl1aBMaScmigUDopK8CfLUdtuKeZuDoOL5YU/0aA84L
GWzAV1NUhtEG7/aIDiyL8uqvc151Zrz1xpZpNzB2k1ErgFdMMcvNxqPZou6y/MIh9mVxAZRzWpGf
BAh6dsgmJoIGsOkH/YFdE1OgrAENXcrezoM+JBMNLHhIYwmbwIoXN4BjsBg9+g6ZPcOXnaQ94JDZ
P1CBAj/OEfCurinO2koRwX6En2lERjtpOiMrYXlE1fQyAKYp5ckkVWKJjhl8vgJHIBRpGsuzk5du
DGb3R0SNWWQElGcUbxrMi6xiVqzZAmpclvNHRnRDy5U9+FGHCgwJA6dkiOZyBN1D/+9MeQuI8zYE
+xtGeUOoqnTKGL2NGWtRcBLNOAr8EyBWTi1rV7QzSDhUNQr16fPuE3zh+doprw/Sa9XtgVEKNeyn
l0SuA0KNm4NO+xXNfP9zs49FOU2hXG+FRDspSCx7mR8/gwY5s28PHf2uzqVC7unbNEtyqrKziSON
e/qXiADEywbI7/2puwyJvEVyOYtjysSaCDtxNoEie0yGRmV5BFllaeGedNawTMazG3kLrWrVKfI9
cdKExLoIxICBgc7RgZ68EiAdMlHOgqb/uco95VRAegg/svYgDWZOmR3mQE1H+keG9QrKr2XjRs4n
4Ut8cG7r32IDR2HVeZWXC4vfwZIpJQdw6mZ2UuRsNvvK6WYvyrli3em9rmsgMO2cH7hwcZkk1tPp
jUDGTuXMlVZXXdKia4Mf64LrHeCFgaRqwBIK8UE/ECWFDQ1u3FCPfY6Mr6r9TJUqIyz2pHiIvGo5
Uea4y83Vz/IX+1dyIB/YcQo5wSI4Su+BTO8P3gFdDdPGvym3WKUI7sbGGzSNb82TVcHmZ32qrHhy
RHjRpUBXdH7OyO80X3Svga54Cs1pOAjObdcyTxdm7v86M6WdpHLOet7Wb+DjTL+t+05AqiDvHWwG
tWfusA7dPQjYoiZVmmvOEDkgOG+xJDHpBdaB4vCiAazKv/58PW0qhdoxOJJZBjhiko2ay12fWnGb
guJzeIa4FFK8mFvg3BU4tHcMZeXEMbHqSWt1FA53UketpKo7FI+ZqUtR0vV6Q72p5v/BL9PbektN
SLSpqZrn9JLAH+oWtvvrnS+7Zsx7EBpTKdscwc4otjj3wGcMAYRt39DnYUwi1PKOCm5g/QceOGvB
U5yKLFE1YyT+juzEfzfGeQ8wGn1ZanYGv+vIaRyCTNLwqpN+f9iLPN3ANw/FTX15OyaS8onfQqWE
ixcMq1XaXbF6BOFGOTSFGmxkHVLbTPzZGKMh2Gk9e0E1MM6UlRXaCohLCes0au0+8wD+jJU29gC+
FY1EjgxhfshUGqnVhIdO75NoAT07XXVkQXYfsVE4feybqV3L3lshvKsQ79jM7J1q9Gow4C4mJTzg
/4lH+pdCzTYeilHBQ0LtwI87vLRF+aOebftEytgprTQxk3rKV1JFrOYeluZ+38QeoHaPuszOpvcy
DC94cgEwJx669BTQssJWPrKrF5kTVrPVkML8Xh4znfylHoFs4sYynpXoo69AviVnc7hEGpbMOUVR
dsGSt+RDTMrRijUkGSe9PlGy9m8gUSsQgA3rEu5jJTMGskWey+77hcM+yuP5dogcgpgi3MCHdoBw
4J0/B03wGCdEFS/cOQ4C7edhXLyLEf0LrgxZJmkB1fhwZ3nk7+RtFW8m8R4QfJAJV98Q2fVM/4xB
BHlVFXxlXopiVj6nE2FpOyPy+zoJ6Vogazv0xt2+Zep5+i1d9Bqu4KAKdfdutgYfHSzGqc+smGQR
NNBphxsy7V61IJNbq5yq8i1EFujdRhTRjosjkAEaGQtnLi4XpAsohnkipOsWy9y7rWeA47xGhjCk
Ue6sjPUwKnpfA5R4ZACNVjZxsPz6MD8PAcQ52gclJbHX/GbjcKb4U/JUqI4ymEEgXbdb+u0WuOze
M1Q2xW6NYTxJ39KAjWYd+ZRBTWL46Qr33HHQxh2CfR07yWy07e3olo6wAWtsxm+KpnmxDpt20ONy
QzSh9DEWNLi8IYGIwi19zy1KHQde/ZKLHuRQDQh3GPHs5fY8jwYpoStd2HMhy+Vh+5t2Un0NasQ1
LgcXAnKQ3zgbFYHQZjh6uZBIGVkSEkUrFPvk3GXCigS33aN4E5Njgw68cL6Qh+RHUEBy1jF3pZdQ
7CgByPtmzed7nVILYXThqhGNzQ4d5LyidCC9m2rg14Aw0juTj7rVOjENRYBVd0UaHbeY1rQsRhvS
sey3+yMEuHStqps7FxvDwVWnBkYhS/fIRZeus/hz+CFjC5Dt7ti3msAHYsikNNIIOAE4i/+aohpc
HQLgOwmE77X7QzC64v+JTzuP2mya7L9EhOP0KU6eBa/4a05te/UKhXSZULXbC30u/Jdmv9WzIVbm
pbCBSwL64QFF4KYzBRBtooD7gEyi3KbtKKVbM/62y3SAck5YuZnLyZJJaQLcsgMUeCR5w/xJJOLv
nSN3IMkw9vWB/Ngwu0TBKf9GQ5ut4NJpYoYfe6ehTTqGZyK1rOgP98JNItPDJ0LSJkX19yRbG82j
bAtDYyL71h59XaEy0i2j302Qx/PWVN1yhpa6XjwxKPS3I6hmK8q2t8OJTo0xLChuATiwt9pOMF4w
nbiSItRispeoAiS5tGPK9l945DBI+21eGHOXjkwiHzcWtFVu34p4xuJxArTQ4XPg4s8wIEv3CHAY
rar/pqmm/KMlME1Hncg7wnckZGagNnfdjpC2r70GIaBWxElV606BwM0CslVrBc7JQfgsQup01l37
5V7Z+YCLiQ2RHRnMpe6PqjQatw1zG1RKZkHdTdf2OGXs1aKAr5cUdnyUd1bwCyilJyKZf1wsLgRM
UDOJzmH4rPV0rjZYCd3S6TVVXR/4kOOEAolN42VxpkvygYOVz2QwkyG1Pj03tuf3K+YxnGKxzNab
qGnJuUmBbLGNOWl++EUg8vqsA3mMs5dS2NS2S0dBLduWes9abX9xmIW2MBr6+g3FzyGcnWNn5Sbb
rdSBGp8MjzDVuE3mgTq2RzThqdVeqlDp7SGYQ1DDNDdKL+/XhmbaPNnrs3VidSjfrueO0CsZfhtv
R+UPegnoNnc6NjjC0MF7W5G6CvoRZSaxC3NJsaNqpF9nA26InJd98tpf2NmiG7MbE5+yK8QCrdyk
ZvYUpvpSLcxzvU9yEDunFkR90tK7NecV0KQxNGole8XjT7fdmMJy4aG+MQqm++KUPTAqci/btzTp
ezIHD+oDtdjmaAQllvZ9UY1FTT+N3mX8jLG5DF8Lf1Dfi750DVLVAtkeV/wpE8ENTgbxbduYrQd5
1er7wuoa+4D+FhYVt1xQSYLpmDLLawGCtr0Prerzx0hBEbh7FDK7LfXwNgNK/SQfLHojK9QgMTsH
btm35VnzoYp+q7fVLoYhB/4uUT+e5GqSouIDhcEpHoAs7/gHee0paGI2C/5rVphe5HzMzr5YS9iS
XXhkUJCSpPhJDw7p6EYtfUFY7LV/seG/Yi+5jirHNC93yyUqTP+LeHIpvyQCFzuJNYbotXP5vr92
iqHauGeeB8DWaZbTUuIQy/hJT0HAH+azPDLaPVDWYDPk1yYgKuFNjj9gdHlIqsJve9Aao2VonqYQ
qXYcBCQlipvzMoa2GylM4t4MtOYto/rjgfApTCRD4xBH4TjErEzRQL39b01G/umOVCg7UwFoeirO
Kvbdu/OJk7gaU4QRVdXOmO/hNMGXq+2aNjV+vMrqobJTzD3C96RdA7xYWsoLZm6KsZGYjxGXRitN
bR+D2GsnIfygplHiK3Bm9nqxqS0AHigsq5nuu4GDYkNXwQaRNGr2OnjttAk34eSXilmpO0ZW5lca
ege99hgOhKmTMLbxy8utRYxym5tZgfFpVI6yKsVKURgTMM4LSWvSTVhWQtJz81uenfm8x3LQLnEL
pEdVziOhgv0csPHgxQFG1cTAc3q8DtMwQSD6OJ1lAQSpnuSPdUzednrLuugd5bqUkvNGW5TNzaQe
c8wzddCdT3uY1oYbp4PednuSOkrmdmcxnmAKi1VixOzFYc3whmYgkAmCIZGRpqQLkycvhcPZXLcZ
/BTJ3rEQsWZNIVtupEcaTtY9rk8rR9iJp0nEteUIayqcS/7l2tWiEG8JhrO03s1bbwHsAnaoJmKE
7/qB+0UQhi0fmCj375YW2zy2hGXmXhZwNeMXI9nnoeYApjXERhV5q4bVaKKlckfgqIB7jkl8Piqo
hXhVfsROzP4rlsSkp92afZRmJTuVF9mHY4C9Cm3BOTV9aZR/s+W5rjm2ms7jFmBGO65/ckBQt25Y
W1/xigooEOY7ZBmh0+8lROkc1n69DbX3YTa9d7SPP1Zoa7Hgvaf1KSCyNG8rvStumLfJj1YpeX60
IH7QkVCOgWs2J1BLKzGTJEeaTNPoM2r/GmFx6QQTw+8i6f2txRSeg/QnUjdnsjf9ivnRb0Fqy4xi
0ABH48SkNobi5EeaBzcFMlVJnYTF3GEImrOCya2XscP4tpdoX4OE9UkQVlCMU1W6PGxtlQEL71sq
gt3ueRKJUqNSlTy6RJOpD/d+siD9rosVY1za7hO1BWNbs7wUilEDWZsqud6rdR1H0gqPJ+cOXtoh
23y8LiU0oDMfHzgrNmvbZC0aV3DcvXYgZAlAKlJO3Jrd3w5IngPqcHXxVTLFjvacJBQBpQ34WBIk
LyxmtZlaOuLGkjJN+CrMqErca/EW6W9uUpZz31x7bc9pw3U4BdC2TXVbYhDB/IzUpX4y03xSyHfB
4TGaMIKxX7bbDdizTJcyHhtX3j9dAlal6C7a5qzSDKV3bS9znxl6Gv81pUDyWRlcUPOE/9MgCBfu
RGH+HPV8GgsBJn0gVCH+hQfK27ptMtpZ64IqhKvzw6/cW4rVcawP+pIKHoxYUbShCnivi4AsqiOn
I64z+CpS/u+NqToVKHUtIejkvqrE9P6JnlL67K3tB+6+iO3VfM/F5p3CeTEgp/1/3l+FmMv2WvjW
utyTxnJA5VNYgxKdgKPNBylQKrFjnrTSgV025F6WDV2Bi38lKVaFWI8PX2uPkW3/sH//3EDlwvSd
PsK6xl+AvRDYqB/FU+59BK3Er3Cro/Fe0jdbHxNc0kk4AwWy/DflVMXHLB2VLw2il+DoIWhYob9l
H5RrUsGPNQaBsK8oKj5CEDe/CPP2DZiauam94L2p3rqIn6j7NXgX/M8wOdO7NQ4dzlGuL+2telZg
0u/CQfDY8UR+AeuSES8y5h7K4bYegST3J1vTxFbC5+GlwTnxQR9B3mbKdS/FShlWJFGSgQo1PNgF
hYvY/p5/hJgxfFQchHXmCsiJBfmKQwucl8+O2t2Fog/uzpAsi51wODFlRLYztL9q2/foRt+W2O86
NDQp3x79VyhXWZECf7HXRv88J9Qqc6408yeYxvkLJSlP8Vmf1Qh0K0hkZXgO2A75YVZAA638kMs9
oMfby7/iV9VaAtbbJLbAxe1w//EyAZGj8c3bxQCWvRFhgNqlHoF32WNxr7aqn0xLNUWQUMAUmd6t
06Bky96V3QMot1FqDxx+fCJzTxrvZUqzApFanZZSleKC5E24st5AW2yPDAYU9ZuMSuea8hH0d5GF
WLlMcy8kJhWkd64j6ThSMuYpqclKKCREcff4hGBzXsLvvjb6gmfUFafVxBxHvlx+GikCqUYpwSlj
oH9r+20AA1JrYTktXVxQ3QL/Q/VA+HrEF72+GsU7hQi4AZo+lAB0yb4T+3z7zZNkqe4j17iR/vOL
oJ8k+H3gRrBZcSw5Gt8k+oKzboXn+TxypmBjmUd4pne4N/Ln5wX3WQbuCMZti1mN0haXwPoRYpSD
SSoBMegWXgK/bq8K47nIx4g1UZozRozT2i85C7Zt35pq151Wav+pr1yc4qMLA9zXOfH+vpUoTToV
o1gXqxUn4qv7k1e+EQ3Er+AVzz+0cHui0Ew8jrEzkPInZi8gdNX46/gkRHZA5mjwMnygaEuUNXIX
9O3EngH1iWhxo0jeUfnk2q320mr89q86KvCMq58/8bV0u0oqI/ZwxVWjlsn7oDWdXX20/VWHm3Cw
eh9veIGHmPOea84RCP9m/Eb7RrXq7zbnkM9b91OxsitWXNqYn6LzaIKdh+o48dMVvPeO8sBYhbEJ
kRytE7lrXpahxKO9fhmpAd7lyBCdyv/WxHiaM+KJrsV3+RJxogft2w/4htsN90WWtJHyXFFiPagq
SR58Q+mwAIR9yIIFv4gTvf69mIqyXGjmcoj/il93iCNbPsvgeCzNVHH5cFPUp39uxZS5CP0VPpT+
pqlFDHaCDMSoEHITg/WjS28vWo9jmJCcG/Eno1RnoRbScYBnKA5sJDUFv2op3p6Syw6HxZY3tyDe
Doi3d8CLYuRcQ8kn7tGoqzUHgV2ss840nvlSqH/RrieAbWihNgPH4Np53CBxFAST1uEYpmIMFTF1
OJJz5lqlRRhqymqXBqoGtK/rOF39apsRNBjbMqfR1OKPAYvKWfsHaHtMQmt8kkzxsQDSJ8X1ekCv
CNrjLqn2RCgsmybuw5H2Ae1j8/APlASQaFt8WGIatzjvm/1vljMwrfS9+BPhEbbP6/YCnDKDo3UG
Tucr84AqWljPFouEgd3QrHTkw6vrYQehuIP1Ms9cxFHgO9SUpcl/hMiDAxlC3PENhRws/kakzMd/
Om11/s+WQ5J2V16MmdeGkO5eeQPRZ4U4Lroufgfx7mPTztVgeN9B88+YVk2YkCWLRk3EyEnCKzZr
lX463kERV+lNNfZf9Mm5V5VMENmVDvLZzj4KD6pMkynKeQmq8F4PW+Lp0pPARl7qo79mwaZU9Qlm
iaNUrrNSNsl7u9TpPXAO/0fDz9So43GeLIVcJP4yZbXDj66Fij5cLEcjpeS2bUAD5tHLEBZcNSFM
qB9hp3rhaV/rsXRz4iHYMDNoi6GUAzv3IJOY5sZKkQKtNepfglyu9YKDbeRgi3tV5L+HbngFVWs7
KJ3Ol+x8d9C1df5xXM70VTN64NbovfLCA0Au9sinKKTtfqOmwuRU2vspuNDT23CLd1ywVr1TXBdz
llmVjaFsoRBSBNGaqrNuvd8+aD8usTOLm4PHB6Yi6QDHzoNx0CO5nkrku4JcJ9edTcP+r8RKnDjQ
b30caL/LTOfkG5LoQ3oAlQl/h0oo7W6F6eXa6toj1wcX3f1dM+bq7QcOnJJdBfW69ItI+oqCowL7
vu0JKmrAyQvez68fRxcIyTr/JJBYUnGu1gm6q1Z8P2N5+zl/aN3YyoWqyY9DztwFZygQf1cVofaO
xTbGQLXsULj2x7kr16hla/UDVVK23j60Jmvl+WKj9zQS3knuNaEQG470y/7B+K90HbNRb0Me2Bsj
tiBMa9VWke+qP49IDjLQNjSDGKy+clk83x3iMy6JieMm5JaSunJk/KTvjgQqCTinAphcxV1O9j1o
tWPjLXBWKy8UT5Gqst24an+GMwwOzRONYhD+/8HZ5LDMcXAwGUgRjk+SP6DwBgs9ZUt+K4KUYEoD
t+qgrCKjtX7D2M5bRHHRd1zuj9fIlhp8ir554GCVL7rN9ewW+TXK42mw3z38ItI4Ph5Glp1rqptW
1KGoqNbifoSMuWHrYoxV1MVesXiyIBTCi2cYprbJGggfSMkqIRmQhey80NtwmJtNIKEArV4DcyMt
PN0AD9/oJCQyGzaP4urNf0aBm2fld0GI323oh+I4lZLJzCPaEMirJhpQ+DauBcOjBmBUbCk44vys
3vfTjhS8pzNjgTLg0oE3ojnLXqYjDnkKXpJAeB0iwIsNEPjg36YjrFptUKG5AtxM5wsjzT9+vnm8
qTP/Nlr9tjrDQajsSiDi6QNY1ui0sFE3g3cj3lA27eAgedftgukgXi0gKUh4MbPkSo7AD6ALxEuk
4WmFxb1k35ZYViKvwM9oxlz4QVorn0ncMaBvzdBP3jb+pBwg44J2p55QrwdPbsdooS18G4P0ogTi
ZeFVyVEFCImxi9SIfjX3lN/KNPnbyOR3tq9LDId7Ep0MiYNnQa1uDsSfJBRRuUvpThU0SQei7+31
O3lbb6Dka7eiDcc+4QAKUhLyiEvmDKBJc5NWa3l7zJIyDFQPaYV6BJR4slTomhc14GKEjkO+cw5I
WNXQSDrqoKT4csuxlvEODW1Jw1CXVNqncwxZgPAfpGjD63+tcdKLfl8BmFs+g8xNURL/8d15wmAK
h+AL3ClTTVyJbHwDzSAnR6CBHtrT78a1CnHq63FhbRTt6cm/Pmr2X1Zqr0JPLDGWDusyJTdU0SlB
W6SARjPPhI6OW2pWigxgFRZikFeFPedyoKIYXjsUtGNhriL9LcwkiNqJVYI1spMBH9OB/f+iDope
d0qfd90YffE56kuKsbIqXTkffH4xu2XiiKvSoZnbPyryy7okjT/fYmEOfgPGMTfSiHvYYNm2FBch
eOZBVyOZ+e6orRl7Kz0zwVyL3GJznWnjNJPZpOGnsuc/cmlBfjbChe6qFoxvblBU+W0FGqSlay6R
5gyvQr/G/FFEGo4O+dPUeHoqHEbPalr1pfrYkVA7IDyFbVvl5RvN0M99uX0Hta/R91ZaVEgyI2mS
clbpxCW0phRvlEIBC5vZKFODNVezbAPUVFMflC0YWAsUCAwYa+do+No9/4ctVh3+k7YYGjRc8Iki
eFGtcZ8B+BAGe5aNRBeere2n9bK6USWiMaWcSuLMHpns6MIsyjjmGfTqDyTKcup+B8KmZ0X3UmJx
ug2Mh++TXQUhqSMtgk3JYdHC2sq3nkq4ETpyCcazcYf/Mq/tznzgyhOSUDaQmAVyr056WfUaw+SQ
us16BQVN4l1rD5M6xf6SpumTZqkhg3EMTtcBb5SdNu1EuJynt1PJ6OyzDAQCdOpKRLHhOyhDn+kO
ZH6thsQRnaF0c2xRgEATaKOBzbH3Mxqs3NtpaJu+grjaF2UeT0QOuc7vtL8QAguq2Um2lomiE5vN
e3sSrO7QKGY6+GaXyy06P/9k4us+Piba5BCWhJvREjcG4g1HVqb7FFDoZo5Dpa34rEnuUEFgfUe+
0yqqZ0lC13vQkCANEl5HyEq1aDVLmIrqOB9R00DkbC8BfMgBkTHgl/Qare3grLAqDjdG9x5aINzU
s4DjplHFQd2NPiwovrZUTJVqIDWeQQwEaBR4uEdRNPEcYQXZLPUcq5NlCloq1IxF9GAd+y/YvX87
nKUSrhgSqS/lcXykx2TQ6jeIjj4mj9DQka06dY5ZRubktHvHx5S7SgLhsVX3XsKxoS9sLjPYs+U1
QoSZWbprA4ZN2JJe16IuL5FWfwyVguRP2vq6vVoLcmuTCQLktgZbZ5VXbsmH3i/6tWw1Xhm9C2TG
poMSftuDCHtn6DmjsQ+MNaSeXcQt7iaEO7Pd8LxbNHyVHvD6yPfLyEXQj0yREyN6GycBvGSBbzS1
GSZAr1uG1erxRfxzElFH+5ou3bYxntcXbW9h++sTlnGrFvNFagJADgnk9YnH8qYlsKKDIhqY8+S8
pck/oqYT1uCrkPwoCJNUsepDQfKunUHb+ifyYfiNWfQdh80MwP6P+ImLKHfWbtJ4RlvFymESfI5b
q6HGGnNiBxmdRbKWyps9qLkPhRRdYxE1kJ2cYMaA8vucYvAVWBonZ6nAsW5mx46XULFja8sr2htL
znUpb4RMnznED2X0szNOt8BZH6mD6hSkZ6wnfhx1rDYAAilDf8mrl4NFpQ6Ce7PZ7AEol6uLWghv
jHZhE/ZmbjPcYVeEAp+RU0vblAiDxD67gqCnsb9gBmkMhuzh7zaSyJU+weB0qVp8OKf5hPD5KUOt
v9f4yYWge3vU/2zCrkx51hNTSm1cFSMxgVB09m1P+lRUQiO3Z4zvg9S+tjvVQzFShCpacKBwkCJF
ACSWrIqK3NNORydZjvrVji3YAw2/PAY1D66qmFQcJytWRIKJV9KOrkznrLXAP/XKNcU/Q7ruCl6r
Ye6bqGla8l4lQLiKxg7k5LzQgBEvuj8lJgu78OGt3Hrq7rRURe6nsaGi63qkJ/tIth2Nx8+JS3XV
c4xRMAhMhyv9H6hfdcqBlBWg+Qc5APr3NYwzk08Be9LL1tYZQo4bh0xrm9nq8/iEUs0RCCOHNiOB
8mpXBKmoaIuzJ/c5q47TtTu/lISturOBYie+00MUeTPn87ts3AYLSGJ9MJyjurJ/YPnYL8zV3i/Q
pW2IB0MdMQIVNs9sA74uXErU1TY54U4Uy+Nu+n9RYrVoxNhWFBKP3cC6rwmQkffY2NZMH0S7MlZy
bwA/5qWahishAg8E+Hq8qRvoLKPRYsb+vv+mEy/ytXyCoSVZctohOyQGmucmMfQacagyED+ICRwH
V84i52aFmTSB9xV3CcMkEE3EJrqQhBwDzc3p7Lf9LUf4o8ScqSydXS8ruuzec1aMH3E9ScnVyBVa
jDSP7HvXAUJ4uIBfXBJbiAZSK/j4/+Wyc5TSyee9C1cj51tbqBC/8EbFZNLr7AvjN6LyI23BSoUq
HZyq0GOT3lz6OL0g2QiKvmv3BbOzGceB3CKfoTyw4+SLcq0dlztFG1WEVTiAzBGDakBQVuRYOJ2x
sJ2v99CVuYqmrrEOjoHwR/IYywaLA23cqsy/m9crEiRLG/HrQ2f41jbDniNiUfrAyyZ6mCPoOubW
uOoSw5/HRzv/xi5VY7EGUEgzQjDrz+wv3YS9XKq0+tx9phNsecs8/fiwExoIxjewRC1CAeo6ZiX+
yVqLsDzY3mqfacowBIlLslfzhi+bI5u00B76VH0EbML+CYpWPIgMBABpbGUqxJrpE1RToYuI494/
3IaycRlkXCp/8npLCYVnC25xvrMtWc6SgcBNuHFYYCuJ6Js20Afx1WcTDu/4+ZtR5q5mbfX4jmnJ
v9zeWAEKc/S9OvRg2rUSv64Ref3Q7r4qnr08eIvCm+J1cc0FYEnnDownDC+S+yFe8xUgvMdnxJ4A
pCRtrxJNNvAHSmIqiBVT4TfdiwTJVrEb1XvdqteW/3rGBDiWXS3ZG0u1xVmHcRTsrymtrqP1U7DL
iGvJ7lJgpmXDgrUMsC8l7P72gGQe/PvpGgWxtQqJljAwHkRKrtosY7ymtNozeIA+khDVvh14L1oA
8dvsJ7qbF7vKMr3hE6U7x5rsGF9mMKkWqb68gXxmDejwZ+8BmhU1reWFa9efWjCUG0+r6eCtttJZ
7pglQOORsujqHWhbO+MV5ozU7+6GL/76iviopQbLz1tAdEURqYmtTKWZntBkmrXSK24hEO14/8KP
E+OVmzv4MlNFWzM3sln+0QMPFKtJzpK7QJHSY+TNh5U9J64GBMCDFOKlzizhfWOLXsk0Hzl0G34r
6fM9Sr3NlxC/QUt7FjEDjRg+1v5OoAatv0xWqza8/iq18xquTDCFeEAqy/IakxeA+9FYSikm50IY
e0X2DTO+9rf+rkdWhN08x4M0Owf+4iSrFuNb1vO6VYcw222M6o8qRP+DPQr1t8842N1zU7oEC+oa
nbNinLKj5Q6glSyUa5mmPBZAEQg5m4PPioemb0RriNKYnkSfceX21y5dnr9MWna9lzp96GTatsJI
+hROiniO/SvmevBC4xd7FjM9bRSCd6SviXlalP1w6vUYj8Kpg4bhSk171AKzWMPwZr97u57xynsN
gemSK2lMVc9krQvwUaEr4cOo3F7FXQ2nXhxdyYRKQUrv+/MWy278hDTInkZYhZy3U7xLNc6eZXAw
dIDOGrjSRARYYjttYSzYu3L3kqPqJxxZamLJbj6an2gUhh0i5XUH1qgl1Lh1wUSjJorMqkTaC/C5
8UYd7GGMF2rD8dUsWI7Kef16IoMmbdnFl4qUEnogbQZE54WzIi7L1RhJjC0GDH/gZ7DIQTBpM/QW
lRrWz6XgdqgSPHCJVtHMsOhgZLZtcwD16eYcHyPjuZmgqXFrN7SDayrkoJN8xNg2TT5Gw1oav+wV
5alyJAtEooIk167M2ZUUILoAusnxqkZhCmXvZAMzkQ31sJLpTgOHVKTvm12cliP+LmPW1MM9rt7v
zxaWD6w0rCC7aFgL9nI42YtUilH4kNM/Yh+sQZJfgAAufdnquVMeWvKgWbbiY7OajeNap9MIbASB
COCTjA9fFGZmdnixx3warAnhmwheCRpTWWjZW4swn0QxWQMNiOxsAyUP6RFRnunpaWpd51WYkZTQ
O1XTjtkf1YyyrEVYqSVuNaOy4biXCsRAXkOrWkKNYMZnAl16EjMGMDuHMrwoSQKaaOofUt/y9j7J
D8PtjvbPgpvaMN5ACvJmzYiMDzV8BGdDhxeGRsMU7Ztkj5Z9UUpFp5jK/sGVbpkTF+HwcHjLDxHd
lGH2rI/Naj/PgTB/cLbBtKvDOR1Y4BOMDVal+jMVl/GfbnjCAJjEtZkoYDf8fqQpMAvRnQo3q5KK
9LMCZhs2quT1oo9ZqNsLCO9GN77cg61VNY0XOjHYtVIz8i+Okf9yLF59JMxhsNe4fa6y4QMRYkuk
VBlw88mrOyx6xaL9G+QW5ugfdURLjndC02MxZEehGfW058C6qlhwZzBqisib0fBU5iiiEVkvVkUi
zH6+8hQggtYHLRN2Nyvpk8/cIXUMW0khhZ621uYrK244PF0b1ul8cwdLQ2v6srmhc4J7au91Nhlc
Fezugs+5moQyXkO34u4vf1g4650ZDSj0PSadQHf0tglJZYl+B1ZvaTvx48zkPmwN7e/StQGO+31a
55C3PWbIMs23ybmDDBu2Vz3uHUQRxLHV8EzQvr12ZINlNtdIK+y0rOXICKA0NNF/7l/RMJyikv9x
Vhr3qd7QM3mUlr3Gt51jdi8HV7RmLXzaudbsu9QrFrB6NUuZ1iwOo35xStrorOcYfw3BI6rFieag
lsRNDPmSysVIV3WjrYxAKWASDqNS/Kj64p3qHf3H5B5vAgmokVXwcda0OP8/Dnla0G9U9Azsl6hV
d5GNwOzwG9vjW8BwvKndEk/SoQkZWCUO02aGK+PNT4OhD9PXmtGRgXVsJmHN1XR74yoiCIj8pG4m
G4A6BTQCPywMszPEIw0EvYcHmKLJFoGyErydvvTL5qGHt0AzFjXsIQz1qHhWbRP5dRc3IGew/eSn
e/wILXNQzBEyDit8ilSEczUSH31ULgNgeF5cjYPY0lZ371X3JQb9e/eSPtxD1pN1P6U2BrMeQmIL
WD8zHqljhBIgPZmP0d2HD3Het7QsoyopC9mR7SmX+JMmNVOnCY5qiDF15elgp9eqIoq8rMqMhP8y
wBcqlnSESznnKtEjOAsn2qn2rn6UN9Jms5dNU8hNudwi3ZnoOW8+4Xio+4x96Un29ebTsAtEiO9C
OmoGEDddOdAA4c9/UY2Xj4AkWpKMIfKuAvwxfqP/6qEF08Nt+aoLaWUlWGPmODvUFNLTLXxuYMBS
SAZuM+l5R43gmXfoZ/J5OizwPaV0BpQk1AaI1SnCCApscHXmxvITL87Wd8DsfKyOINK5KK9H+xmG
HiHaVsTGVWPCqTCOS3+MCzM4/QyBOhh8IsfTDCqDSyXNSN1/bsivh+HeTFvLurpXZNWSxN88dEFM
5y0kI0E3P8iYNQBV7AaOCzAW1Vu4e4pmeaxWAFKDGzb1EmyXKkYmPfJcT+DLOPhzixsdc1P/xiKt
X35LzBdU3eJ3raIPXv/ypk/A66CM9k8yPxugcq4OPWS3wJftaP3mFzeo/V5GrlgbbyuWaD8Eap2E
d/xPktxgnWKx+52I/FMY47Hi80sWT8uLEfctoc/1237O0Mp3buuccSIh/oFcxw/wWxb25Z0PG2dP
DST4i61mAh4S4hBVI+fhRov76AkcaHsljA+avvn+Vb+f92eyySiIGBVhCVgSgimCudAvi6KautE6
x5JpPix7X2GJI3XGcEqW/zB0b14GjWR6zbEGECPzp7rSAxE/JYxS5mgGepIsJ8i1rWja2jgslUZ7
oWfchH9Psdz1lXvkDeUwiFOwqxWTiFgzD+2H6sUS5nEfvknxdOfCzftsa+7+lZChgWdwk5dPKU9g
tpBC1VrTnlWzMwD4JhGvmPX5pgb6KfS4WJpSMDkO8CTP2KTVSAUMdod0WpJYeQUcjjPxwztlhiUi
8ewxOPdsh5tmnsVwO2vbpnYwIL7M4ukYnJffrsHpcxbFZq2l6OzFwtnq0Ph+5/6FA/2vm2oIcQbh
exfWqX4kpas4i2YiGsAQP/iCCAQHtORGnrjUYGIz7KOCgfN5Z2N4wVdKTFujcua5lcwJtCR9JL9d
RcBlJ9oY1L6EfuAVAtIcK2pFarG+CwwVuwT0pCAB1acLkeJG+1s3/lTLC0LmRW1tEZ6LDI7pQvuJ
vGsL0zO6ojg2XOZiCvdZmC8ffPQpRRPlpauKO1wHlCclpThYxqkmBaDTHuyixx67eri/SLvKZZ6Z
fGAz5w8ll29jAJ6Zydk4RrtjV9YlwnKjrOGZqebl7LC925CYu1lP4I0Aidr6IRpcLdDdLsE3EaER
lFCHspHuxLY++mCcNQ5gDe//Lxy0CMEkAOdtngB8Ifr0gflR8ibPnK0FHRYJAT5PAUwODg3A1N9q
y70RkMx8HLK9fdrD5qLvNNqBdvdIVyvoPOXxnbBRXl3CMcZ/VwtyEZRjxxuzgY1v5nh/Ud8MDqV8
A9dOdoNsu8l4E3Ul4GYBwuudj8PVAdJoyOk2U9t3bpUuHhQp+sbF6qS/gPPU7RA6YgRW/1d7sgXg
l8vhg17nse92H9kS8D0ZpPZrrBZR7D1u+ZmbL+eAjcahtUXEMD/WGjG/HHeTbR2GC9TAd5RONuD+
bTjUVNpCxOJMXtveyZ5YNal5FxDn6zyvLzXr51v3cQ34DW8ZWWqxyMl9Lpf8F5ZjVCX8a0YCNWCu
16pYgOUcRF0EZ+QX4djD/ZDsky8rpPzg5vbrl8p2tovKvr6p2Ug/bgHUbC5EWtA4HVnT5aHo5D4P
1/GDouRBRzQdEkbMBNxFZnaInNMZgapIja2wkCLcI5nxvK+VYyXdtuU9opryQbfGcM+mHrz7lPJ2
ZXQOBfJ3N2HZBkjCTFZOuDpcWrsWA9F7jWMUEXO6O+W03/XjEdueqR9RwYX3YEmbxu1KA3ABsQDi
O4TshbqgM/JNh5fHM9VrAuKOd1f+0PBIICHIeYSX7snGl9KSWA+1q5bnpxc0u1SLhiBLZCKtXRVO
sf4ZQctezklUPqP0LJOCyp07D0DMB6PvDACxj6pZNwpwnCgi/6mjt2MvOLAitA9pzPKrSunfSDKP
fvq4vhKVWfzBIxi4CStkPQJELtMpzqBMeA4E9kLdkylDOpEWYh6QL+ODlIazOJyZjZ/75P1/8nDa
55T3sxVExvX0nW4W+8GApSRdlOw18kCnm0M6aNspbICMkqLPM09jRJhxnQQBMAp4VKKCA+T9R++Q
tItdYQW8xc9NOVzX8A9eIcWe87bxUyS1W30b/K2zso1WmoEHpefHUuaIw/Kx1/+oLcE+dv+aNYlt
JXE0Q/aQWjDasiPcQupSloZsrbjrYW4kx7+xCWFmvB+k2B7cEkuZlJCPfVAhTxXuKflk4NEx2dUH
YB+aI9ncaehEWe+ZIi1hUYRCh/QeOaMLjgbuVxNBBN4I7ME8NJ6wO67qjhgMAWk1cB00V7dVgL5A
CzYGqlhTlL53XLMcrJHmfEYsGRc7oEmLWfEIDNjU5uE7BD9rcgUTVUfi/CQ8pAhEVpK45/c9RBDM
k8qj00vsao4rexQJy0NV8K66xOhGlUjOjDtVnAAtaFKpB3BlY4y1bzaQjhihDz2oGIdmAM45pk20
kwJ8vhDXv5+MozYeOlnSgLb5kgyM0qA7uIIFXxv79EnxTMFnhQU7iAwH9d4Xk+MbZw6loUTpgkuW
S7ITY6Whq5d2p8TTMdufdTKusbzlmnzd8L+aT7k5BH43jVtYdsyCi8XE+58nDY5rP7rn5Vtx9/V/
fxYci8mTcGu+1a0n3FHCvTa3iMel5Dx2LljkQBPTIrqLWOrUyWuJqOZyUprSyvGRnrJiVyfD6Tun
VeKUTq3aYl7qid4vARA7z8GoaRpgKIN4Mdxil6TmgyvYo4W1F8neEwgxtLwjopuZOHTvQi/nbbQ5
HutrT6cn9wOqyqulLPQLaA2XdQxcetS2o/u8dnXIjxw9l1oL7o/xM3qnE2Yuy0MR2sCMH08KkkuZ
KjQmEpLvurFoCGgiDOCB0xkRprXIq+deKfPPye2NRKbhSCmMTXbO7uuFSTYzhaNYb1VaRyEdiMsY
Kggw15G1F/6G6ECjjrvi0rG1wiUXlgQcWBDLgtV9zyVmmuerX9cdFP4xwhofX8IA21Xk95eyjEzn
+TW1TaroLLcb5o+4GVoSCgVTMaqKsXgUvIJLC6KeCmiqwx/AUg5eAhXy1JMpApx2mJbFwVKely9H
yUbBfOK7LuVzwlhChaXeUY4nBeKS7kVa1cSutgtS/N3ium7IXPiivEEIdXF44DFn8LiDw+N7kWAr
XnBzBgKWtWoW9CWyXC1kBohvldElx2b2pp4SFzRs3pzgA2+QVnHspoMzb9IVQo9CyZn4iNwCpCv1
V9FMwYynXTOzcex1Fz+QaUsgG5AJ28Jp6+6ezzvnxELO7YyiHtYn+TcfEQPGC7S9Ck2PIty7/0d/
633y6rLC9+YLJjD3H83NkwxtuC/LEFREoWaGdU62Z99bd6KCu+icwo1SvA2Usli5yFQC2Mvds5mQ
bmlRfK+PGTwDauZZl15NgskzaHW2DZ8UkX+wObVFa9nHU178AB5FSQRjQ1I9LLkFYzAxw4I3rL/2
4GDadC9kg3Um88O4B1A06HcCcGn0ST2w/8u2QnOEA8rnUHF0OLmoxDeVzK+ROt0pU8dBPJlQ9byk
cOqMUlt8S3jfQjiaQycq5NxpjP7Q/lI7yciUVVFrXgPinEeS3BzAd64ib8xGVOXxfJG46kaVbFL7
oU0wNY+hrlTTmnZkdmggna6xrGzBW+xOxjpuKLr2QbGuUYNwv5eRBq2DZ377Nd3hKoKt/Fsoeg3v
AgHsd3TX2dHb1QQNyqC7YyasmkLKeo0VCgw2eGvsr5MmQGSNYoInvLYNqaLi9uoVvEXWJCcYvvbg
pIKISWPhIUO29/Z2X5inYTx3ErqpYrj6U+t5JAd7OKXgbMjQcBsIME+pvlCl24LXgjtx93K0QsYT
4dIZeIuq99lxKbuXEi6XfyKaG2GvWJDjsltD2ZADZNxRHgqT1pBLq+6jDfhh+tm43Y/wK6SvwU+h
eH65U12bFWgpmtom72SLQkJkmIdgG5itVnTrPFWK/cjiYXyT8NXQ0yFR57WLhK+O06Fzpa/UI/CP
3FvGz68QcYDiRDWUh8LgzoyERnyVnqCdLAG/FHc1za3lKr7ddsWb/bRDpk+MqxpLXWjKsy9b0SZo
4H2oRL5RsCywAnwfimRXTqKxg7Q2CofFyt84aMDKXxY6TClAhR54wgxszpd6/C+LlbblXuYI3EtC
cGkfjHhUoE8sG0LbiW+1rzZu55vFvtyMAGEMKldb+KoagWuf6EDMW9JHpvQwucgAGhLKmwWYnpwO
7tQ/aQ6fM8wvdVZ7Z2JU+KE5C8AdhXh6q+seSPnKMI/fdbzKKhfcSZCN1RspYNsyU+2IwY4GoBGz
htdhZ5uJ6HjrBFIlxcJl3fky8BYn3o4HAw0khVt3qcTjGJQU0z4jZqVBVWeiSVHThwMbHHI+dUSI
u/vNzm04Lq0MJka5cf+R6TA+nQu0cw4g7vusSFETPFRWEoaqbX6/n60TIA3fAJh0ZP4JWbezeZPW
JMvEMLdy73xN88n5zKR7OEfpauJ4r9KdpgTFFiELQNw45zKQQRl2dAos3KLtCCIjrcBGcgKxuZYV
0EjGfHi0B4tiaxx64e/EYv+gCBoRWscIfve96/qJKrd8oE7Z6MoOo71/0otfcf/SA8/ig+4pTC2q
CPJFuT4lNCdS8imEZc1XTqKL3/AUXIT/2/zMTNIcx7JYP2KHbzNvsO6wNp5hGUtZ4ExxuQe1UypI
PZqe7WWCd9iHUIcMFY65k+Gf/kIme7CXlpIWlfkwgaWezFtZBCO3r8WL1JSmWjBfpvTl2Jsukmf5
RkwCcnaSWWEsxbMi3iKTSOIRlhqxUBQFqUnmv0rI/U67CkR9yhoyUJrRwVwKiKlvm9cwB03TO64Z
RrSNpiUwPVnSlXv5c0sTZXOSljCK89FsNeeFBD9gfxQeJ++3BsYyCta3yCiYAevwD4jiieEPXMcR
Tfui+lHXd9P4gMVubLoPdO0NojKyKoUyE7YnL9IEvf+l9h8p2OXHp96QTY0KhSmdPSsY0tJu22Xf
zk4XzjNZWUeNZhaDZEO8pHj8JbYNO507iCoRNeTCsz3yJ5IaTiPwaUrqXRYAgvl2w8VJyfRQl3f9
JsGc8Kzne+i8/gNFJ79a6J+2Cf7JluRMFCtfXJxb6erdWBD+QboPOT1yewXR0EJUbiKAaDAhHNAK
oZQwFwQ9Is66AtRv0BkO48/zjOD2wQrsaTCRkqAiHXZGtTMZ0tfB2QSvYLpKmVYpGGvIL1ijxdvP
Bpzmh2rt3KjwyuQliCC6kOACKUu9dP0ezpMdZ8VIRagtw3dhRlqnvgxW/7hbtoZgWQxHpVdzilfJ
8mopP1KmDxTCDM1hD8wEvqDRJqUFJmLnaPR67qLo8V+SwypzeCRQU3a72ID2cKrCg6AVh3SZ+ft3
8wCS+iUHUfE4aQknF5m69VoOskbOiZGaP+lfbY9RxioiWHmBIGq/EmCRv5nrlt76m6Q6HUhPxkAD
clHGHexZmhasphbEuJmKaHY23imDz98JtbdkLbxhkdgMwGuakCN40SgpVohv0teSJ1mPVAhf2W4A
I7k3XBDuQsPq7IkP/kvdBTbmkDXNcFwqN7WXq2G05WWeimhPC9+hVx83UkE4MlyjeaxXY0/yv+81
/FLL+Po+CQDLMQqP+OU3GqVy7KJCbj/p2JynQ32S88Pzr2sqPPH0z+TLf5sLpKWE05/dAmEXPXRL
7hIHbQSaasv7QmIoJedoI1l7a/IEAEL3e7jc6r0rI5iWzArHtMtu4U/OVBlxRh6AYL6FLk0qJ7tj
i9cwbGVh1RQetTsTkxmQIYDlyL3y1N3oBZmhkncsHoaJWLKPTahM3IfqHnkAkmO5U5Qs8Fc2Kqd8
fU97qaoyV8VZ2jXGFRRW716v5PzVBhGXgDqrnWjE5ZDO5Rv2mtzLcrJa9ol2JakXjaV3y5wjqZQH
zIqPfjmfT/iD+x3C7VrR6uA6Q7ydhiL0YmDKaggCKZ/rm6A61KRs2BqWrKf8XuCr9wDpqOXQ99hi
xIKda8g9FYSMu3N5b/FBOKC1qchT1Uwub5Ezs4dzrkZyks3nBFQ2bruQiKB78AouIaC8ZHPCTau4
aDccCMUL9xK3U16uqLk7ENYH4tBYCcEZV2512vFUExWTOSEZGQfsyKFWq1Frgyw6MmI6nxjmtScF
Zgeg0aMjFoMDCbYx/A3zcFs1TWqTvI/wKC6DzThoRFdQm1gjq8TTc1cJPPq5wZQu1uFo0y6/518z
3clfrQ4bbZQY43RjUNznEIFWznhWTGyNWxuWVkWCNmEM7r2K52k7xYTbQWdE3Npr2ia5f6FaS6Uc
57mbR1Nwu4rJjNYeKixXr6h+gt7/IPwl6WZJIrTlUVXa823Xq0Hz3qkT9r8JjlG00S3L+p88QNQl
4tCPB6D8PwBqjryk1ZwNniLJN0rhrj6GIAc6yaWiYDkJSyhbC1kT36U+FpH5Rkyb7LY9V1/fOjNh
ksKPVfXrjVe1nnWGY4Tl0479EEEBylynegOc1208c/iqxxrehPJyvhs09K4l4BjAm18RcKsFXpaW
6IBPS7fxjrd16fXRNi6ha5ECgllYFfDeVFGP9BD74DNX1AUPtAzfRp0U5df45eBfr2p32OyepUIS
clqzUDxHj/CXnpMO57HcrYZMr2xiNy1cyEI5XtPz9LhAvN48wKzM2sMBP/evL2EE8FFVbUiB++fL
HASyzgofI/PssfaaBkxL24hRUhbBJLcwsRfHQnp/pSvacda5Ef+zhbiaU0+0Ggy31Q1P6gQglMVZ
5UtrXia/NSP6chccJsPk7VsT6C1n1tsopOwkwh3xbN6CvhzfBtP5FqgXNn66TDQJWDs3hx+yWgSj
ctGvsM/TLQ1PN9Z9ZB2jCLi0SCTw1ZQyFUtLpDSkjoUa4ZoDK7DBgtU9951ygf1LWaO3ffbV2XRs
nACeZYHubhdceciwcnUfeJuuhc9tmbDTqEgA0pWN4h8ObCdrIjF7nrjacSwCogLAY3LJO+WRUrC1
rpt7JP/eo9Zl2M6C4+zVDnhakz2kQZsCAy+h7Cl3AmMfevuHVRmuoaztdbZb0eMfS7YYv3hjuRB5
OvLHlNxvEE48IEqXLVaEDno4NO2ZChAVLY0uNvfWYvRlIIlnWAEHUv+2ue1Iz17Ui/Qtc8LFy1bV
EXfDfnFGwKecomA4EE83YYEggjY97s29rBjeB4l0dvrZS3Z/g5nGiU9mPvI7LI4zJEpQEwhNpOTa
T35V43U/y39Q5qdUAy3GrOl1JjPiFNvKdpZrY6BfLUlQJUvf4M4H7B7SVNpkQ6HolwfGJojE+aKK
G6N+Wrws5c4OlWN5SDY1v8NzF4ivBwzhN8vKI7mIocEdbkPa1EpbWwoImNzUrOsvUNOYEEdh4PBN
4+2cvNOhZ32b6WHZKX4lrAGoHrrrnmX00871Uvo7jt0nc2Ag1LxDhXVnys+aJP2FPcGaHxKOSaw3
4PeAjAHR0qYCs0ElovPpz+CrdsikRW20rghCXN4XdVORcG38GNueJxcb2sLdHWrFcE+JYZldSzL1
iBV6iNhLRh1/2LNHE9ejaSZzn3PveFEIvhiTpDw+n/kwVGKMxePrdLRrB0KkqA1fkFvRFaWychwC
0Kts/4zOxuDjlZhAf/Q8MJ1+6ECLZjxHRAG3EwvsxXYXs+o33s8ZK42KnsL2OsJDvpnvXjfDX/Aa
1ULjhmLObtX/qBcmGG4nvtghfGCivgGbLHPz+UI3vzNyl2PmQHyuGKjBkhQsLUIY7ESoHoiFKdBj
GSz/Pdz8nDzW6Ve+MRmMma5ATY4gUDiICM6lYgUvR2FjUuKy9XNmOKhcoSgEJ6A3bOA15zfui/X8
v1yBox7k8WrHV6V6QJBf73a9ZCswgLS148x7ZLLyHSzeoSQc/lMbsrLGIeP2hqkml1RXoKrpiNu5
LnkqixidMMum8/ngJsdyqhyOSeZw1P6+QPOnNPcfJRhwanf7dVPKLK5m0ZlmCOhVCk+5QIUy/1y6
CZ/yn3OtH7MMoWN9nrj9Uzl3ux5VKe2c2Ey+uU+BERDJ04nUVvuZpTHDrcNSm+7Ng8WSIOegd/a3
lSq8SLIa+q1p3yS+k+DKwTPHV3i8PtFyLrkAl74pXmOHSgZVQcHN8GKjJdAneIb4KzFmxwz6nKEe
W4yHQutrFZE7aBSuCy7ENHlPS+VcO2h1ORs5pHrRaKg6ool/fOa/DlXWug166IOLP45f0b5jVndw
QsyqyX4uVFUX3is8XTztKPppj9QMFCJqx/XBWSmY2My3t2Guy7GYFxUCOXwqQBvNxoAlhXCHK8t6
wCJzcnJePb2pTVIGnxy0d9xgrfFDvu4Znk7Q5WD5rHJuNbIT04LEs0CXC3N9fyHXz2qtVbUaoCDK
hu7rDY70dfdYJUGtdFdAHSs6/2rbzMPYDyyUb+snHvjzInrSaGCffHnyNjZnMU8W8UmcQQBIRLCP
cRYOawnOtoDyaMY59wtXsm5JrlEMXQritaUY7FnRncaBYSehLi66g6KwPA4QS8ytWmchQwVE9IZY
URa0GEC/2/MU7QVOQNf2RjypHkjnqhlGMiwQ26tRTcGq7X0t5JLG3ERGkfhhdaUASo5KsFqbhra1
M+86rKRGOFt7XnbV0T9Qg6XypHHCd8QBvuq4xoImfTx3CqdHiDfuLptnruLlrhm/lp0+yWe2LJca
B1KI14F4b9sxO+iZPiRLYUgzOfLsopbTnac4t+yxvKVOLVVnMBCu1kgQ14Ta9QO9TmntvYv/Jwy1
/COU6n91HiwnxzLDkqOU9BwX88T5o/bOWE5QUn0ZNYqUST5YLOjsFYF+d9a4geaSj1ycjtK2C5Zc
IOHMNvnThfHkG28L2QC6fV6j8C982CYsOWHrRIHrTBuCGNMixNgGCe+Vr/k12+aT0QgSaZoyEXeM
/CGbMucQc5zag79I9LNzzrw+SXjhdEcq9sNi5Vxj08CkqwTRxffE0KzE5IRXXGE9SlGr2lcRjLWH
mwvLZJ6HF5zUOzJPEamL/Qfmkerh4Zh3McdLugOHwD+QhBzdJJsemSAMc8UtzfaXhpqo5RF/TZgc
faHR43lpnUKXv2sEQRpSmMUO6uUOqsOqDYFu1B24FEhTEV+amKauE3id9AZXs1YZYNUdQFw98SbM
LzaA63rwk+RudARkMuMVs4ErggBW6Bus2jEV8SzYeiLM1Y64BVPvJGDOmBfJhWvtkbzjkxPgQRrg
a6nFZFmBaC+rDCe/w3KLqPQ4ccuXJKg3YSfRmLuwugQH4GABXLC9Iu59D4BDmmOZ8jKbe7U9+4nq
0mBEYszR0IRrHPhPMCNtFULu3bh8k24WWwLtje13fL7eDPZc6IV75lpWEUNn2TgL2lip/nJeoWLy
KkxNQG1mH2U4RfJJKMvEHUnx2SoHCJBSgPZUD5bM0QAu9pkAOF0ZqQQVac9Y4ky7vHjkINwVsyNF
paT6WF3teadaoYnPYxX4kg6lnrKhQBMdmZnJJxYs/Th4eEXRx4Ic1szxlufP0nGzvhIgRYKQIcAD
Dp3fRNGWtxryVcJtYm92uQsNX8bbCS9n+9ZCVeefCvRRyPW5GGtEbvrpDER2lfqYVBbJVEFoM/5H
JqNE8sqw6zGXccXj2LJIYN3ZKSczw2kd9bjUYgpoUobeddQh70TOA086MTwNMMLMm1+gR1beFIk9
T1aZ7/SR+iXkpNMjsAKLfvU/28NUPPjg3kgWRTp9OgUx69AJ8d0ql4Sve3y8xiUlwha4jWaL1CCL
MAgrjj8E+Y88tI69nJAVA8HVb/LUIPZ9wAFkS5RHtCWdLVFJXLbD8CREzL8qmPueKW5hERrzTZUJ
eeMQ7NnrbWZtpU1CaKpE0wka7/exzja/SjfbyboNRfql/SbbTtqbaM1LLv5/o2gq5qftpQCMTSEN
sJOE2MJXDDE5pOVdUJMPyCaB7iFFrGWBSl7GBs2UgHOlZYKBSVYCCPkj8qNfiddbwZI8pi96VaeN
T0fkoJUUh4v5F4+3ALLoKSwoBhHoq41Z+SV2uKZB/XQXA4MxLNxn+jvEKkz2OCVVYQDcsSpp/bya
aDb3wh7Ogo3nbFijVXZcYPZJPAiSFgiuuBQ+POHUtQBRXfBFK3iS53lXfnv8BHKBTCVRkY8FOCIW
10diCR3kiH5+dAEng6UaEZHkBdjCyaGFTDqvvOVBmcQLoIY1dND1rI3yggS6u7ROjRQ2EU5mxXpD
bQStfXB5sv9KeWeZU6TySCnzdV5fAVfdIzcY3C5CP/DyaJ1fcgbdW7eF9hVUV8ggtGcSHC/A52E/
EzehKHas0w49zyaw/Q9yWbdwGljXrAG6E+9wXUZKp7QxkDbRwsUDx/oNp1JLU+qK6qiq6uIBHYxD
9F1hb88PUj251ggxJ/NnQZ+4VD+nU2KHw9n8fsp7w8eOTkFkt/50aW+dLcMlV8gMgFi/oghceDdV
Efrz/aEj1hZzsMk/2ctngD3iTCvIsTczhROVJm7aKCp3alA5AZJDb5cwepft6Lv389CyihvoYvYB
fuUhJt2iiAIkWQ7TceF7yQqF83l8Yoc9Z3wIzk6KF9pURyBTq2/+v5r60C+HYHa55dVGvLWI5kUx
C9+P/qQmaiunSZYFx/QPhF8fd/S/dOdLmLZdQ7FaAuREEGvdVyVIYyaq9cZqbKJ9piffFyhaUMGv
F+o/E8X9eUtATiMQSrdneAKXsJ64Ri+hYgU2Ep6j41rUNqxsPjwnan42H2hcVxZeq03wDoifQxkb
427lkJwq0YXRNwgpnPAVNZrSTFfJlUeJMjLEM6jEbebH4Wrswyb4X25F84cW1mLVS3OQd+IEXskp
dNvf6RG4zTEs/s1J8dKYtwXA+WN4jTn1rAw0HhPBD/nE+bhOhRdnJ1QnQX7n15Y0cUh2slXoMclh
cQN8bHM40XawDAhIr36m5MYXQE0mc5UPUa6so8C5l1EvNmDrI7adFig+HbN+YhGPTmmpknKMtcmv
BICqCd4ScUfd5ITVhcxD0dL5LIUe/CtDEsdDntBMo+DsVjHVLpRONqChDVeMH3uTmYrj+oZ8s3Sm
78Id6xAlwFoqidpBY3qXqEMWo6uy2k7gAJ0ecu2uIENy86xXzIqA9SOgabMcJnePpdTgiu0Irfm9
X41/XNmHJLsDWx/eZWk+kQlr1M7vaeNfeCPO6qXGxbvp610mrtFBqbJ/EWIDBRwGmipe5+8choBM
wwx1gNiTVt8NtQmhTFQHIufwL10KvFdkHTp6q+7b20lMaUVQyNoQUFFBytqjXbE05ICaqkkuez6b
X4arIhu9iQGu/rU/9N9D1r+HumuYbdTWPQNVJIJjecNq3nY4uYa7vDAbdBWDnbSlr79H89XBkLV7
gWupHhfIhCBTbuHMw428ZxpXEffPxmzvWxYpWYL/r4Qp5RTSFq9RJ8qEE3aBlYKvhio8HMhQzjzH
W2HZ/VP+O25GQI2VuHqxHWabaGDs3om8KBAOuj9fLZ29wBzKpaMvbiPuxD1Z0qfyL4DGs2tX85sa
N5mJL0bhwFZhHklR8G41VS4Pr8qK03DwsNENm/jua4nGj4ufbE7i6zm1Va0DKXoQ7SmhJyk88dkb
EFCStrhCEw3BE2DmhMbCCzmOb/d+cfy5pi5XDpDv3lVrs2lXwXkCp+QANte3DDzidHuRmxVs9mxf
ky14hj+8naS6jlOIG/hMgADaZ1T+bPNwc8++5Gm4ah8Yjo/9rFNqh1JsnND38MqiHLQ48FNuWm3o
5Tu8GpeemruRX4mKOI1btJD1fmeAp6wy1o1WM3gIULWdcTaQwgtLzQdMe9QnoDkUJDUMjC5FrXx/
Zt4gih0AykafAG+Gjn0bRJTTuqbZ9G66ZQE2EOFGyVirJ8LLwMfUK7CWmdUoviUMJT0zH686LNkj
2WHVcHudIDDxaobxufNgdymLo/XWHa5BHxbiK2uecqhQNneJOC8bhyM52/00aobayiyzJgKB3o+I
Ud+gqPAaXimW1Q9Q6Ubj4fT/OSZKxWW5ZpXfoXgbypld/d5JabafTjmryHxEFgFNjc51D3CFVcpd
2tHFbQYZu3QFbNca54H84A0oBtv1vrs3sRI2cwARunMA2QphaW/jnmYmDThEHTXn351MuW8wNs1r
B3HiXXIqEnNrwXOiSgFW1luGYz6cXvgsCCDDpeyYpe7aDoQQVgwDcMpWuKqJHCpUFKDAcDS4iOA3
V25/WXqs7cOJVKUeE905/1OJ9uc8AZsQFeQKNsPLGV9QF6DBZUz0YsGw6mdju555I4zmBwdObEKn
DcBIZ2GR118PNP1gVampTDewX3/Yf5Fn8UIzzz9e7PQSWR3/wnS7+d1Tina0pTfeR7FhoufV0K/Q
fp3hMO8XoTsWk+tr90vZxtLkF9aaNiYFZbZETHi3hE70EWbCxMQ+Xh6/eKb8DCc4w7liZYXY5lQl
ahhRossNIhT4Lrh07uJAG/yAQ59jJMCg+8KO+VYWwBjDv2KWraLHu3qGfPTncLIm263FMpNQjB/q
bnyugX9YjnslK3qaDGROnc4qn8PNGdEDYnEHPvR4SbdjcFKB+PMmbq7cYfN7dpMeVytqc7EhT0Hr
T1PddcPHCX3wx95UEtWmFKLfbzhSIDI+7rFk8Raw3jdF/wvgQx9IoRYPsPCR6EkYqhIO5wZDHfuq
3EX4wRdAfLNzN4L0Bu8v/jIjackVVjho8+qF2+mOkj5B2pmRrIWHpTYyY87fa/z7WNyda2msHB2F
5wtHP4ChpNzQhsilR7EGeTgOo+SMKFyb22yF6JR0zKsvZvUudZr/jhkcJE0ei4PE7LnhPrkjAPsU
j3d82vEA42eHdVvsLmAlAbsoRBTAvu1kKT5fwYbdT5HvB5Yf3bz+QQtsVbd50CtwCCoC4GByKg6p
OvB5VUCrpysJiE3taommXORNXKt3dpYeA+N/KxLKlUcIbjJDjjZkaw2ri6KM4hAX/4twyF+BoCwz
ntvtBEwWwpml8QL7+NKh/an5ioe+dBs7wGyktbGFYr41JvbRFnLpyUfjC1UX0OKZMZntYDd8CFeu
DPozoGxY2M+1KTyGVJaARow6JoBY/q0ADitRTMHoTOmh2fBRw15fPti/oHli8vsplk+lHw3ZBa28
b29E8oMNKAkDODB2vHIlIMAkRFB68kjxv2cmyBIfzsfWWzmgjG+2Hh5FgHtNkpRdCljnQKn8ahTa
thcZk1LwQJVEUrTJUpHSjXT3bLo0f7gPDeYDmq8LAv35R3qlcvLEMoXSYUrsGxAgYqzwlb+5LTD6
ey/ttqeBX+AZGzueQbUaJ5ZvjZZAaCaTh17m4CfJPfM/Y43ySYhVVFTZcmNEQ2pB3e3+TTXUrJ8r
gLc/cD4kYDb66acdq9tp4tm21IZk5+DlQf1Rvd+RlcxbXXjNkRsGm10t+ckNz49Cevi5sGfQnfPG
v1Bga3nzF5FihdNwdglnNOq4ZK6FkhlCXGBr+uLaTdsfRR/ZUgAFajjvtnY7wQafJVWxBwPr10O2
De4so6pb7FDaDx/my3KuNjeRLXxRJbNQVcjffayeRdoY9N7r2fdIHuSLi2EfTJAgoupZxnQjUymw
2hjSl+wJ+FyGiVJAIGtG19uM0R1csTwyvJV3KQwm8wQlTOSNwGNBb8tletonG+IFaplddrUprjcr
MVny8bz2GeTGc2OulN4dEr2jWMY+VC5JYOAMiI/wnmrYfFKlTp/h8tlxn4InALpE+FvGUIucQlSq
jcHLLd4fxUPyKm6yVE5SZIEBcFKDHSmAvbQcpzYY5zDsXCU1f1KwwhbxGkz0pSFduPVmJ+WqqL1m
4LAXnuyiHXI/4nr65FItJfQvYW+JMIWZWoRb4eXox+5YrPFDlSevw1hJmgf4Ff1eumBMkcLD8dny
Rmm1yIa0QzIEL0rfs1UvURzU9+ialws8+PiedXQjhkuZIQIZAwt3a+3CN9w/wMCQ8TyB2QwtOHNN
A0JCkiAq6cd6Mv1VpnUOgj+ws5R9ckeiMjP8jvwLJTclsFKWpMvQNV7ztwnRMSAStA4pSlNtG0/S
LuoOUJlBlF/dv68g0Hk9xSAN5XUmcxhvzNmJkXlVKB7SFZGHAPadq3fL5fyRuqLMaVvuAoE8Oirv
HBJaW2svSfYUveo7uMJtsdXcreS8OddGqJ4h7/sH7ersIDhB9fDczQsJ1pGyjNJFUgrNk93f1cs9
XA89m96r4pMH8JXaBQECw2QBWt+GjTud7ps2B0hPK+5IwJPbbw2KozDO6EcfsOI82kaCRxImXtOd
GLSP0oFklmSJCVMuF9N6zuFL+nINLMwsAmEsG0Ht7ziBGo/iH6kaTKebJJmfXb+siIw4qE+665Y+
W/mJB9dAmMHnf6vR4KTf/lrkPAeo6ViuRAbYudaxY0l1+TB4nVZHXTB2PDAAmxE97AJLwjErD1ZI
p6irK98CxQiHS+4rUfQ5f9FrGUnCbeP3VBcIjGAVS6iUiT0blXzD+v36/jaZ8+S65FX1TK/N3BCa
6+wewSuSPf/8GMdK5ue2QVGfFDktdughIbXujqpt9aZJv+fIMHIaV6tGKFB0z6oYHsKpml9mD48m
QVB9WYEtB6uHHwDWDniqdcQpfZ+XqCMdYU9vQKmEj+EbPA+gBN3sVNOYAwc3f8etVtGbHRQxWAlG
aTD7vOvF11qgRRWHP1gX7Irq+DzaLod+apVo1IvCMw8aj3pmXHgINVF3FlAgoHlFk6arsC9Az2fX
4dJ2rnAP1n846E16ygMDgmvbU6FYRtry8P0/2nyB4u/gDOP0i6nuPolupm6KUGyX8049UhEbm5LT
PUyaeSjChVOvcOxNcwoWu52wDTD/FRZ0/lVauE4tZUvq8LcGde9D7a7vtqx6RNIG78WdiqzQTEP5
dtxVnHH6thr2Ox9NwZsObouhaTuvwSG6QxQo0WD1Da8zwLuII0tpP0Yu4x/bHIm2ikeTLyXEP4l0
BftwrSyXrWMQlmWOe1oIA3iKZTCpkb/53Vu6+bMzQiWoxfseauBQQCQ0UpNiHKWNCsK2W79S7V69
2gwtWHitI//eMAK6vpON0KD/8AQkWZ9+4c60CzcsoUL0GnQXtIB8o0Szdtx5LxxFTDQ7KDaFCo3t
bV2p1j5Ls9xIhZVzGkysYcLThV6hOnRjQDY/oidl+rcLecZ/opJIZF8xmggdF45fT6/e25xP16lo
p13YuoKyZt44qL492pENnMywJ+pWPeexeSAbi9CN1QVxLxtQ7kHlf01T3dmNP8ozbHwpjCPvz4Nr
qVpY3o1v9fkpeCqBQ2aPv78gza+1KH0pcCn2CTHLf0t1IGcN6/IJyUMGzYgcbFF47BvbzX+lD6Bu
Ta9sswm+8HuX8FX2b+iK91/8N3XQdMcuDqvm+G1nUb+DWMFvy09zBzaohYWM9t93hBXbYJMVs2Wi
SODHHAw1YnavHXEbvIQE42PB2Mk7tCoavmtnhuIoGiUlx9TJ0a4Q6pqYSno1dC60skwuSsM2Vh46
sCXMhHo0V2ht3Q0TYEeZVA17xg6e6QNf7XQFSRb8KpI91QsYdd5phR+wbUYyKCVoh6q4DwxUgMZO
ayJdhQzPSjyLpvL3pIqtz/cp28PJ1xmp+hiSjr1wJTSeDAo5La0WapwN5WtNqgn8mXW4RuWHtQ8r
duQMhwQq/dquY58m0VISG3zEw/MFM4U/TrGK6pX1X6vjGXFJEPXOM0YoUQUKHzTzzYLV8W/y0wWC
j93tF7neC8phlm+11N48KWSaTB1KM2IGmWJ5r5MED1WQfaw4ucNd9Z/U8xtQcW9gIGr3JGtWUuKx
942YijG6AeeyIea09+talwzuMSekHoFuua6PL4ziDSz2uSs3MjgRqnUeBFjuxNeJbYnPamN/H3XZ
HzOPZfwQQFcbF18f/F0l477UCwIZG4CfFGe/HgZBDC+a7yzuFN1dFZrptudvlcXptJxVDod6YpEL
czfZ42Aqppp7hO6YUg2JcEU5O82GlFZ6gkdS7Y+Asef2MiLsK9hIZo4E9O9T4TsQ649wwKef7W0q
cKqgIq72bFae7Zql+FQpRZ1f6g768g0yPTDqJjeeb3gids3SitoAEoZIv6Pf/1C5ImBTskALenvs
O/EcXhrpcOapce1LZIlA4PXzm4MuhfLBYsoQ903Qu90AiiskEv3JWy4cWxBr/0jDK3jxwmOgZ9Jq
uzH8MZgDYykrZANDL9Dp7IgtJFE4D1HmuiEdtCly4MlPzKJ6HxtyZRNdKHi357u3kNczDVlDExZk
sc5dSqpjkhY4hoS0HsglJnn1Z0HuWL8GFOVYgOlioDCCQr63vYouDeMd4d6MCvtR6xxJuDzsy4vC
5YljUH4X1TAxbRwdkySUbtTs7gSEaXvq/V01Vnpq8BvN7NUcC80wx9I7+wqpSk9/FSzu8Wjw89y2
C+CXIynPWkzsmTmpFkwvsNyX8VJQIkJJsefyZOkZkO/KNbT5pqyxlbO/hSt/xkADdJHej5Gn7EYh
LfPET1Vt779i+f6jXN5Z3ZED17gOU8reMV7lLauiaGIlwPsOw2TNoPLzC08HDjbO3G/I7Exhc26A
Xl7SV138KGz+9pCmSr4vU+cz9YLm+E4TrBqYEBTBfLSsPxBCNT0PVIMFwwnnaVW4udROKuu5mfPx
LJCKDW13C5rOqFY8TjwAWEA/TCfM85nqdtASb32f3U0fbEAVgwBVklZQor9lGJe9AWFf0GBU69Rd
A50G+A1tDoDLfvQV2EiNW+8mx73wlVPDnY3C4oj6Fp4wsWBrvDlANDQeg469KOjcHH53El+1IYNQ
POJngxNZHaTzDAMwEaBSAYwtcGt/r1g/fvcQxIp2f/3FX8z0FyY5kXg/JuoC44nHT4/mS7hn7T2q
ewUc0L2F82JKRCTP/BUGqafecPl2DBcDXms7qdprcRHWI7mjQMJrMZXkrKxxIO7XYVeuipv9/NN7
KWoke9lCs7xbNYZ4jCPR4NSzWXzodc2wZH4FgDoitKg1jNsPmaEPLUFkp86isgJApu1IUGD3LPqI
LX5+7c8UtN87gcQ8jAEiNUyK8AnWy00TS2o8deLCUG0fyYDJJfmmCOyLCkT76XSKeOT3XpZToizG
h/dQQENVBS2n2D+t/h34ZEXislTz5MoVVKXUbwx0qtsvZzp/bKrKFzmYziw0TDzZf6MMVewwM2Bd
czdiEtg+YH4M5Q3rcMrKpzygC0ch9xhWDO9MMVPwGV74RhdqZKcOPBNwo2IdxcfQFiWIVSYh7k+3
vZmxPqgm9+PB3CAugcZdVKgpwp1utimPfEMtmyi647pyShzkorl0BEq+bewBbfbpV58NKqbCM7KU
Ja6a1pLkGiVeMUKQWYLGFUeVzxWfwezqJXz5/0GdrFrLxgyAdZICcP0C/EfFajURtNncvUtiMame
6H9aKcS3Udw4d1cMTsjK/O6r1CpB0LRx56hm/67PVWrx+eYULdMFSvbQ001ZNLcfzCb74sjw2rQZ
up7AFAA3k7s9UBfYRmcUuXIDBP+owDgcBvBPfVyPOzvtlUyTOZ6B2nTF30JO5acsoub3TZwVgz7U
NBBFingM4lPBRsIjR8dQG20hY+/M1BZk2nlS8CyFVnId4L3KdAkpKvMSMdfBpqJvJ2T5WKP/AdN1
31eTvmd7zs5bk9U6HCUGQc1Qth55D44KJJVhX4qGQGcWe62nGdQ5GjblbV7IDJPdLjqxbtX0459Q
a3qH8Xa6KP3e1PZv6s3kx6hp6xj9E0EVAeoGQAUb9voCbyqzGAZNmH9romvOZkNQAdmNTrSBb5Mj
+UegBmhAtE/r0WkcQDYP2SqMp6VFX6/jxyMegWFA8MSy3GMR+9VszuZSZ+JSWcA8r7gTbNicTT1t
vIiL/L8X4yENXVTtBqND/iPVI+9/AmZHTWlw20hcT2YDDxYmV84qVcvJqN1us1Hth+HtOtDwErm3
P2ZhUNADcU9U9UswNpVkCnED7GVHeZUxshcgBWQT3iM6wQY78aV2swi5zyKCU9L/aSlEgWKLS/pW
f5yGHKCqKZ0z3FCIJlun5v3oeDQ5jQoSneMIRd6hMZfKZqiKX6/8J3asx0Ut34bWlSD5P2VjQIru
wgElRFnr/rYiBSPV4Vfsfkji2CWzY5J5P3jPNq57Iz47hoA9qTxnfBeGRVjVrYWtl7jwAMgNQdrP
JRUGXZwDxqRPFbfW/1KXcm2CricHt8XOnk1jWdamiw938oTeTOJLcgjKPZlZWaTlI7cQ+79Rvpjm
HAAKooeM4IWT4Np9GknbqbNHKRgf8EwY6nuLBd26vK6wFYucNazqb324XLHDmUt+KXMPoET3RzGr
1sFxK5D8SlWHpqJ+1R4559TyLlZb2QmkTHmDDsJ21DXVof3FiLtlvtjCSzM/SeQ4GbXDU3HJdwPr
d6/m8AtqXQsuaK9pHGSOajlq9lYgiMypqPtPkvIyNxjiOda6IpK3a0lC5nnxOXxI3+zG5MGDVFUv
+wl47MBdX3k/O3+dBAiiSHNx8/o1QYJmtd3O32gY9c0/GoSCzFHzW4YMQBKm8+XLMBSvc6bASeyV
qJWl98w05zpO2UNMMqg76+pZ8YCQC6N2+h4kLeMkwHF9wFHKLr0PaxSn9z+/UM2P4U3dM7NwUSi5
iwhvjsjJoXtK4ezwSeACXQTx/0NiMyVH7xr74ZdBR5MvTrelgJnQ4g1XgGMk22E8LAXQaPPpioA0
fbFYbOPDluzhNvjMOv5wfqnWZ/JSgCawAXLMFWSxWTKNi7G8dWMW6FQoLvrscfJvb/vZ1mYP94v9
Aq7rJjUqpHYFGDm/ptY+WYj55e506T1eEKfkRWOwHpGUtIFnhX8hoIDH/fZfcHIYsCLs6CegnxU7
ZfvoFYrMAi05/Cy5X1jQ9B/+SHxbrpWkb/E5KpnGWuQw0ncuL4m2x93eNrkfTUjZVjnt+8L2WyDQ
QlFXtRda/cka3ehmWZwzkVN53qlrSwgfu0oqnQ4JAAmCFk8q/UInzt3f9MbsFZeccsYScIFB5Rm/
dlwXk4IkyEnZSZRdhJjRmNlS0WmcT4STU4AjsoI5H9Ka6vX7Jh1+/Ch2ypxkndXWN2Es72SEaeiG
7WVVVDzr0Fwo9v/aXi+KkQ7iOLD2/rvQewrVGlT6VlW2FYrzcUrLXEPw732hYcSsXtRnh383s0tY
H8glZjk1XkZxI9j6qIVeqbO9sdZE2dGFLd8EdXDigPiYvbh/fTT6qiXnoiu53VgRwfUrnVEO/PjQ
lAi64Sl2/kF9e/EwTQDywJgpz2TbDrXLXynCScUMu6Pv8ifzii3IAxcNoMrHvh/jGDXfs7A5Nsp5
LFm2NnCP2tlJP1v2k7tZtt6U9VWWUg75ybOOzlPeCNt0QKd668pJiFDepgJ/ged2ziBaTZhk5LU4
88j/9yGr0UYPo6SGuifVO6FikizlvTNAzwURoOzxxK4g/tw+yKZLd233NwhsmTjRiMmjCT2CoiO0
36YuHy4ovwM1MkFt3YP/HNY5CW9/vpFH+YOk+Q7agVetHl537K7e32R1oy7JoNhwHBy4rGUUSav7
WUu2pdXOPURw7t0b3yI5s3Ng+t0pQnzzEYIefvAzEKUxw1AAWrh/PLQopJ/2nTvcHbW94vZqXDf8
freHnbsvVLjcDU9p/5CHI0e7ab/q70MP6lt7aaFHtqvRSBKgKMXvy1JLxl7XRbE1kDWgVOBC9zEw
8We6MXrjQMP/sUAMJ8Whf97KG5f1+2a2rzuPrXw6DykhaJuFYS2R38sttAPovNteGavWP6gGh+Io
rKcuNEo+LKXmKNv9+Dq9cLEjYYK3R1elwTR3FGa6jYta1o96tEWFHdjW2ubcYswD5zQnWM5ktlHd
rIywKlo99RDOto2TyKLErf3G4TATJ4Ye8bY4BCmhcSu3L7l/NhyVm3fOsqcfKT46jW2/4mWHF2n5
vn44cfxIgvRae5O4owm+diPaBxU51xMQ1BOaQyebAmmy0hd/JqtUc+3O3Cc5QQLk7NNbVXjoth1v
WXQrl+qN+LVAJba5DEXV9Xa58b0ZYltqxz7wXaEEGGBQYNsG28F3mMcA6wqgqh9Qd40/q/EkujMb
thGHpZ2Gvp/vSVoLlU7gD8URaTV5UKTq7OP/I+uhSSebflvrbRGqNArUXHl4QfTz7LfdydJx8sI9
l2suFA6SN1v3FCrIXwqek1pXHTCXQnNJboYCWax5GHSeN89Ue7ef2Ywy/RP1T8OHA10o/DaPUl+K
hPrxlcARBSZem8YPaUEbcK0oDY6vC9F6z8Ec+FihDlv1hVQkBfS2h3gL1TtX0PypCCS9zr2x1hpq
7ijMEFUIKtokVmPD51QYdwetGnBRZV6xNahlrBC28CL6ft1azI0zH2rg5p8gU1mEs7WIMhrozYJB
A5YutjkSDJLBSWJWfOgqRgkLgTy6E9QAnt/bLW2CgzQQP22XK5UcqC3U0L9DWWUngVuQVLyh5OkA
zrhoZx6itmBJz33vJrFhoVCMkpc6xnwJFtUS4+NZlsaPO/nKTW36ufWC2BUSIHkOFuVlB7mz37r4
5sJk8Xd7LYcOTiT0EW8PQIQczObegih0fGNS48QMt83XGfb/DwXnB2driseenz92cBtY623qw4bp
Bh2sIZxK+SgB3V54j9K9dvCG+PFz93Eby49f0Uc4nlSxRj/odP+8LwqymhvpYxAPl5G4MxqO1ho0
o1Bpp9pGbbK/bVHu1PXzeZpEy6dxBz8ftnseNMnDpl/kocKr5NmyxTQyWR+cKrFugEJgs0CJNQ4m
E0relHnb8Inyc6M/c4oPeVS9p1S8wOAySyMEkjTMfSTaK0hZ+tKXU2fWJz5FmLwFbQGTmVnnquaH
E9SVkBnrRoAbD/dOabylKy2Ary2Ezge4MEy1lxRIIe9obAJ8Bev64Ad9aONPQ6GqTPKzaPiwt8SX
Bto4yP1TxB1hoLExaeU5Zj2OhubKAtnzUJ2dq7PF/PSpHkOzYzbGozhYlhs/8+rYep2WGrepzTZf
rpu5xQh8c+CAJZ/5Ih4HQjdfIpBykTp7YT+rlrVmKauFEFIXrDZwwjDFXtYOuv7IFH4UI63NKGPc
98uRhBUi5jFBYBPJs8IJyCgZBSOvCgyGlczRPIK8PZiQwWc6+Wk4mmdbUeK1+ouXSDTPS+imHgDS
3ivRgo15kOKygBivLOqvVHTi3bNMLzn5HojHs/1WETaX92ZxXm4SUQOcfmYjwoD0GjX0ziJA6U6G
r88OhJy/Wgm/JSY5EHRu3fSyrFqvOPh6CILgwuHhSknWA77GtgYA4G24X5N1pQx2+QOIBbj0iIe0
Av9iKi0gkyBgjj2M58DgCHeN0eP9qGGOSpbbKvGmb9Qk2FHmcZoMOj3gUX2yujUBFoUt2q6/GTDP
VRksFMmdmvefRwIoqngxg+PlbUj8Fu8YrqG/efDAlKwK7oX6C0an9JHLKhNYywe71UT4F0UmG7LE
c5S7EYH8HpVA31plqwRu6G2tWJWXq5wBiI0da+uiqVlHUlfemm1jvOu0aDPjpCFkPd6hhCJP4anz
mOT3B6HRnAb7C59DU4kalHoM+RNQIOYG0Ya4lheaCgqOqavK+no7J5TjgVMZ3mhNs/daXgJgTf0T
hqmvNWbEyCJc4muIdfUsQOdfOT6ZpZi+DTQJk7wXo9icjaqfKuknAof7bBkQt8Y+S7I2rHLxI6eb
egC19hQIc7hRucEUGbQI/pBAYT2z89SYGn6xSeCRx28pCodRtsTx6LtpInDda//Ef+95qoiQBFh/
PNSPni+jCF0MU0MH1XFJ/gD79tX0Br+fALXotCqih201qKQBKDr2MdvHtwKB6Y/2IJHL85eSjqPj
WqyrEalk+aBrfhz4eXXnppUT90UvBsJy23QHuFrrQsz9pgvrr7KmN3unr4u9UYiwcXqEei0Guf9+
ux8x4SP4w/t8ZfYWsNftS5mvYJFW+xK0WgsFPzrvA8cyKOT7xdRQ7w5HGq8AnL2idVHQMTOUOziF
aoF1dXGouNR7Y3yN6tyPQDfCe86wROuQU6u0M14ppGRxS8KqjhGnJ35J+xAMdJUlrWlb9AYOHO0B
kgV4AGW7gsK+6bYQR9tf7tEzofngRJ2iyV9xLiwbzUgwzGXfZezbfQiR81hyc4GqmA2wTsQJSLyA
4KpfeMQWFQzBWXTr4RlDr8GbMx7JDCMVAULQEgdGfNkCzfcglokxewRDbwPMOC6juIND4fTIsfLq
NeYSy/qdFdH3uhWrnYSAz4XHxZHwBfNTwLRzM/jLXu0CQ/XVQc7rsPNW3Rn9nvThF+3ESULd5hNm
cFH9rYwCrkmEZYdppC/AmGVTbEguZtKK80UqbLOaL9QH/H42h5BaaFNiimGLUTnUxTDTFRXOku0E
tsvAJQk+FKYyLe2WMsSWNKt2i/lTDIO6ZlYoRVilWpiZwLm5bOEzTaI2TSgPuDftERKejIwBh5+g
T9jIuV1KfvierGErTzUIMo7aa7VHd7awBLL384yKZ/4bDIhOcjvmK4MHRQpn+K+S4atNPkaKkEpF
+bV50UKmv9QFf2fry0P6k5qVUZ7jK4sNlmBupqfNNDkUb+mUBIMLfSlQpqhDBfJRuoMTqDz6TcgN
WylnRz/EOOxBholg+f1yYqtD1GyBoqpY3r6bz9NxHg00M9BrXHI8hUp4/aR9JJuLd7Ol5lR4KyaD
Ya60QZGA9TTl/MZJRFdy900OLo9bhD0jZdg+6m8bix3fj8V6VxRoFXEp2mzviu7ukZjCaoyvpAaH
63xFFOORY2+VDLX9HC6EXBxGOHNkQF/ZUZ4ASrIUaYfZCMOGnsrd5RY4c6163fxQ0xnDNZGqFidt
SabSl63+XMBvT6jZBTZTZhaLtPwl9iPc2VdNNNDyJx6BLtTOFCObmdL9IJABF06AtQWxEns8f890
OIxEab70MGRmn5XuXUrMzhNDWRfGkJRZJOLzl380x0vrnRaDqsL0TFOtQ94U6n3dlA3pBK84kbfo
zZFp8tMjldMp4inkSuDFIvopHpHmrG3Ds9prkrgoXqvKA6nqZUTbHiV636eyy5dzOUXTdumOkZMW
UhOzu1GLLUcvWyYjX1h+1RcAF33XmqlcPyZsx1aj3kS7OYiPNtY7v+U90NwQEjLWvL+wb+OxpCF0
wi7coEH303xpG3srARGh+NSHfVY+Uyz7JB/iGaVB1yh52MFzk/rtaKDkgjk2sineOltIkNfqCQT0
p0sjLVDyuFxPRxe+CXcfhnE1Lpi8iClzyKjhNFOq/vEMV7jWTlyRWt/Fnzd/LSARdjSfME/0Q6dy
v7T6MJUJL4FoHkqdtbIJKweUPInmxrIICC/Rq2umbgRtOqFvQEq4anfy0cA/PbwqaHIHxlsaZWYJ
uAdy+/BlKsAChruTmTpbOTS6WMECtPdIt2/wTjJiOyEf/aropHT0uT6cdCX4hhCJamwJClFmmGgs
bfia+FLEBHyJXy/szr1/WAqw9RJ8qK2tZvw63Z+vK5VbDt1Uh5izzsblz88J71ytD1ZNMTS1JENs
gC6G2lHlM8JH9VdXNrTrfguozJgvcoDxYkQ0HEz7jo5pY4yz3EjPXtlJU5seChnTw3SlLTTPKq8A
8iMcT9gOg2vpBynCM1BTRl+pDX5lsqs848MeGRg1mBH7Mjp7oHKa9Jv9aqlCwcd7gorIGcp+jA2w
Ip8KA9OS92yYXU3pF2u9yImG/r5Kkntxc1q7ZTfQRBciAaMYbEXZzufUS4MOSf5HGzz6SzVgFwy9
lnH2lPAjqhXpOgvRYZdQV9/W/Qai2CO8FBQnkdF7MIkef3tq+vLfNM95Uw96z1kXPbuzY1r12qDY
1HRhZSeNpdlKlfdlql70HhnLHzIdAX33gwk43tHJU0nfVR7MQ2uNU5+cWMBX/coorVTSoX3CT9SV
7dJWsY+wGF815RGMNMlPTrV14iGlGL7niECLfmdNaq/JBtikv6EcMMEhf1x+S0Zx+XaN/2yzKEFY
OfiXRha3+IxKW5ug7waUYOTZK+3Rut+KBouiOPQOFqu6JYrZWpMW9ZS2NlOgl3OQmocgoTalmGc6
psh6agbl7zy5ZO5SGt0AlJ6Nm0Coq6fISeSlBLo5Cp0CbvIJLZtd2JGLXCMlBbyOM3rEJpEAvyDI
UhrnX0jpya0UfG43er0IN1HYTuCP7f4yTRCw8fK5j+6WejG4TxZAhHFlPBdYHRi55KvoLi3Nh4N0
zswW2VOshtXiZkEEIpb1qyu5UA9Lx0mk6lon3PeAnfpAjgxr+3hjbfDjwll2+P3zju0VS5D5f3ZS
+NzNPfRcX4DAU3ZIscTQsRBINxojj7R0TlXh5i5PXBGOrRX3ueUTWqoGhIqDFLBXgQELbrURyKJk
DIP3+M1mLm8sCLcwzZ6APvFF5CrhuelXbYfVE7wyJ8HFmn5VftYbtcFXwzUYnNePoc+dNzfum54B
7eWtUvl2ZH2oEtXAOYjJyR36pCczEUJCzBtpzFddsEE7LBc8s1GR4wlBEPhRJkuhU+DS52YvHIK1
vyc2+IsR98K6Ti726aYkQxfxVLKtAg9IFpVgkWpBKq0LBKI4Qrs+mCb2nCqTXNgDvQd1pY6soXhV
JHo+IbwCWlr2PG7mUU8uwdSdFtrY6v0wC2zK1u5SM38FTRLFXH998kAJmGbb5tGRQvsgHJaXncza
SD7I5b2BHj/rXoxB37dtdW72hWw3Z4/aPPlcwTfvVCt8JLjbX6UVFCfqw+co2mjAxVRO0e8ZVVVS
k5zwPYSvn1mLLBsqeTvOa9mMzQ9O8UP5HlZpo28a9/MnTt2TDajc0Wr+0r2LMg2ivmBc46rsLK7E
Xr9eCGyHk1TEIRDr0YitkSf6DuCzE6TOY8B5C0t+l18q48BdagrCOqHj3+d0sal+ydYlvPnpU5dW
QZkMNIofGZ3Bh91+ZiSrpGYWpFpGFCe64UzPPI/DdydL+bdd5dLbLZyker8gJk8rsj0f2fqGN+5S
F39h+LRqo4DbYNN64PQQOvKO9kdY7Z4nRLdN6QlzQAAJNUJYjhudl9jAHXdgLRWcB0/ie+kq6al1
5y73pKXM6rFPXezwzI119rHM0TtvizZhGABffLf/m9uL5Vr2/SXhilH6APXFddqmvLC0TchknzKz
r7kZmyey9ps2eFfJ3PnZaUjmAZJGxqyZvXaXbmsrLcTd6krfyjVknhA7A5lzbfqAUXbrTQJdC2qu
n0wwmeZvOxX4773AP8AcvhZfbhtD8i+UIi+Z4FRAgz+D+wRN44aYP4850Zsi0ylrWc8T0z4VSEA7
eLpzlLXtZDXa2N9n8mI5TbHnkXy5+kFsBSNOFNp8JvFf6cd2OyZCt+xF3fKIAVj0l9nknenD+acd
1udU/bNUg81wmpvnKfuAZH8bVO4zfzdU4FGACCFqGRJK+cVN31bobNpxoJa+HN0lcAvkcosK8AtM
jYubLYfOuwOK4F+CzDLtCG2+P91mi+zZ5hgaZK35QTkeCC/eqjVmx0viOMXEV1bfjWWrdJVk/0R1
e2noJd8Wnla5mimiiEfovqKuNknsbAtCn6zuSlzL46RwHnnP3uXRUJntA9FKr96xlNMhNrv6GxFN
UOFuP8jptR5bhQSWLF3BwvjscO48alhXatfAhNHgg13LtCtYM8qsVCJwRrvZjqBxKFIqUaj6kdfT
EaAsZn4FdRs16ab1rjd/9Cda1ZtvqVEUE3R5gVrcfLPobbe1sXFLjWFH/2OTgzVVSUMOzhp4X51i
ACrI1EKY9B/Fr08rOBiP9d9DbivrP/kD/y5H4f0wAML4clZqKoKBZ5vtFnQUg1H43eDmTJ3V8bdn
x9I3mE/46f8C0o7/XJ/qRiARC3UYnXsETxVjd1WHEyMAPnf8UZtb6ERjLnI2MQXf7WjjTN9pgz40
Ns6ZeL7sOn1mp35rnIBGRN4ZLPhzLhdZdLSSNBEV5qh5Mv4Aths9Ooo5XTp4wxA7du19ZQkO//rt
A2NiHaHwBTAGCmJEhvAjM+4WDyAPz1wjgqcc2Y8x4b1w7/VLXAZls7sNN2sfPRCrDY1fborSkY28
IwAWoJ6KzvuRYAOBfOuBd28RWhpnqezYXOHHuS6Idmj9hEYASBvrVuY9wdJfZGqIR4l+tQB5mCX5
zRR0pvmat4fQsTuZoniBxuY4Sg7VJpLNBquXw/jsRhT7XGlPkSZKBB6A+AxNG1/KA8VJDfm9pWf6
C//2x/ZDA0qqnk0ejoKJT05uDMWCutmGZKTRX0IBzyJfv6TnbMoPcZQ1DQLClVamk+JMr+ui9dCK
ZsuRVWqUgx2jzHn+tPhq0vAYR9WLsgAN3wGesvgzpCJWQdincFvYXSZ1j8YeDKALkAkASJ956xjj
EnNIRO0UlhlytAdV4QvI93kVl9q8hlS9nGwC+JsboRExUX8OOtWMW2pqh0O1SXwsO7vewKOp05+t
0kI17ZLAobeQi8XOt7CrwrrtFdiP4pOXDESc8lNNcuD33CMK35S4OisYTQ2MMIIeHGzIXzXsk5eL
mlzGc4KqWRLLy0Fi7qj4TJrDkjMp7dGL2kmn0EjnvXEWM98sRhSi9lZif9jYEOSQJtDrOQKiO/zj
8JCTzsV3yrfWlXGBhDekobdKxu8mlg7SxnQ1IRruH86btEpWyOTbjoqs7bi5hCrc3UdtcxGheGX/
tJbIiMhLVW8KzU696X3bDTn2wQ4blbYrG0XoQU+YeywGf1pSnBbksmlsT0hB99rtxSWeEn2i7Osw
S5w5e9nRpZciUCc3EjjZssjta+u1o+UKRFDAibLqCoY2aIuG1NzZncI/oQllBGerPkihGnvy6APC
8No+EkCoXeNiwOKJkMZvuQPqS17dZZLyS5oAPYdpXP/oeJYBQv4OjF6/EBz8vCqQaHwZKtO7X1SZ
OwQf76YQx4wpQa03lTIXSs7Ru8iKHctHJcRipfz5TXQaL7cxmB9hbLrYsbvgPKyYUTdM08qT3Owf
SItBMQWQHEja9w6NsXTGVGaPQ75fM9gF3FLZyiRpRdwp3rn3dWAuMa0ZHB7vKJFnMMJLITJJL84c
G+nzx8zpCXKxijYS5/UnKx2Kov/1/j1VhGk2Rjuc8n+M5QE2OqDuyVuqMQ9tcDGulOx/153cThdO
hCpkQA4BrCjJuWYtEn5YSb1LRxm1wNxBWcaUEWwCl3evhNcDPioOpbiVV1ac/GGuB2f6llv7lNon
1ZWWG9fH0h1EXk0StpLolIuW3rJZrYV7F5QHq4nLN5wtFgOAd3Gokhq5p/gLbwhb+0EDMgHshfBm
OPODjdlvkMEo+2wVQKVnEN/x218IDbEi4MoKiO0dzBnwAMVrTl3zgtr+KRNt2dYq+5AVv936S1qQ
GrwSVLfr3FZEiY0svNG3XY1n6nDbNNmwDAAlKjL8QF1atX0dQfojlwG6iB2XjudaySwAwN5tkxVa
Yg78dgwP70mRDJ7bzhgpImUOEQFhQRFGC3ZAX02w4v55WAFiknheLP5r7/KwASdJqiyVVEqvXVAF
B2oK6LXyY65EfDFoQUuUkNo1q6gHhH3DPPKHEDrxkY6D6VkTmyIryDi6WI5c/C5OgSP6YYOzL29a
VXpbUu4BA6PV7azVic07WXqvzo4HZt68zoLiYzcvxo47v5rlAActw24/zDF/q6jQUREQbC7Mpvg7
3xD92RQDzwcn2RQbPj/YVEtPWE/lRZxwl7kNTxYldzRM+HP7gn6m9Una0/dh6bj43R8ghQJW9aWY
3PeTuA3+YQtNWp2iFr/Dsj7uYX4RD0aGamwgQP7TtbgAi1HUElz3lmFxmnTuvtF/CukRx/ZoMXol
rB/ufS7s8bWeFT9ZBbzUoimfxAoYC5/OHC1ui3bfyVk55FR8fJKhVZxkHtdcgivI5HOkbDbV907t
fgHWtuL0X5LW33r8X2JLlyNP1VylRYX/AiUbxP2RKc7lqwqO38i0+A7hpfsdO46Os4+V7y1mXK7I
pMKllF0Q3qAkLNdg/A3cNaNezuDDFVTGTb7I6+8D7m1RpScZL846A/BVdoCPV+HyToG+Xz83cuKb
ncxugATAOu5v8DcpLGBD0lF8PcR6JrlhfTsEB8v3lSTbJiXfqGw2Xc4vmMEPE+GWKQzQFnDk1eTj
XzpATfpfvIFrAFu/nyv5iF125fkLdkZbtPbjq+G4xkZ6wq3pjBn3UinPUOr2FJm1Og61b+Jry6u6
P7rC3Vl1cfrxTVRyvFdOoNVGtvejIV/BVb/v5TwxAmV2ccEEYlo4jkfo4yj7bsVkeq8XKlX8KM48
7H9paQ2A34r9jmglNnxmerpGJ7fidnxkuEMukrpDCFyeHFUYP8Ft7V0d3vNKD4ZDsOxKigfV6FS2
Nr3OlQKIbE9jkNQ3ptJfhxuMT7a5q+Xwjt+EKyRfVLd3jE/TuRSErRu0LcX7Gj4Jpode2WTaAc3u
wLOmfBi8A/2H4hDn8Pn4Z0HD7LnAYq3/qlvjM9Ie5Cflanz55TwES8JD7XLuoB7B4BO6Z78bB+qQ
tqgfrJDeODfZsW4tXeZwRh8fTs2ewdFpwIuPIGQ1xyIqhXVXdpELh2khDavP16Gd4wtAYb0u4N0D
OLaD/qIR76T3y3qG9MV15GZz7muAYw9oxJJTN8uk2X7cMNlJHE4gkbbsgZ+6hc0t9RD0qO+0mR0K
easylFPJbofy3+KzqquwwLSg/8Lv5/Zs9fKwNVV3SaGocCcci5WFOv/gb7xwRwLbjDPey7v7bPw1
tDROTwQjKLjohmjvCUANSzOEtVPvd6U87XwK7JObpuRngRdLe6zQTfEvaVFjvob32l3NRvQ3MIX1
FiIMLimetQrwA7NsI8+qJ5MGuMLbHw9fAtQ7lojgJkkEq2S9fNcdYmAXBqxzS7DBdDZ1K7TtqcEh
UqRE5kzaY7rPUPm/yQLSuusMU8CB5TzxFhTIfl1rj/T+mRoqCJRgbUIwM2MEksXBn/kSR5n2Ci+2
EwvhBuppsnxYnLrl8KdLkU+x69hy+46PNX/W1zFaKPE/z7GnSPg0dzCfF2i6TZbk7ULjIE+zFfmC
UgYzryDfKhfsWVyWZpTxT1ltHG3KGCUZL1yWem6P/zZV8bxnECct6lKoTwbt/oFmGFCrVOWtGl8J
cIKwRr7q9/O/Xgyh4z3WCYziBaBMaXKrqI6fVpBYp3I4s60uE9w/fFux8A5qo3F5gN+9OLqMLpk0
54bobGtvDWTndzD24Ssi44c9/GDguVZMkoakib0SIFHADqrgdEiDt21ADw1+IIfCmyFooOrlIU1n
MV9ym5iEGjEa+DeeJ0ce6Lb3/wyS1iyxvmpKCUlcQD2xJzNC4IC+zMp18Xbs0seV4/Y/58hpOnPQ
vibdkJWgIbSdXfv6YFLllUQlqOzFjKkCxeGFe7k5QH55rFfW2A+mJbTWGclLv5UGqykMxYkJHeRz
9q2fz2ymrDJRmZnHfC5lMZx2WRL5MMbjEdPGSJmMu0llPw58Uemcsb9Azhi4L5AiCVghoe0tqB+C
iCD4Gzy+lR8bgG4bdt0o7TfGS+PVgkf6WFFo+osKjcw7CnpSLWAg14PTYpOdoKrNH+zdoJ3k481J
n+c46uc6ZOMkW2WZkVybCNQFS6E94SNlMx5DfuhBF/af4TAB1zcW47153LOCEu04JGX+wpXcWWJb
ctn6IMq9ONTPMGykbKcBuft0KoZcCoDufhJGqencyzfC9UPRYWE7Vm6YBJEsD5/Xdyx1INHQBZm2
mPQo1Ug/3XN8GyUxl1bFuqJTB5AAYK4sd5JCyoyoAvhpNfNktMzDylr+c35kvxlCDUA9D4m5cmwc
91TFHG5x7kM6342Nzn0w2PQ31Phx7/1+XpboeQGiH+5g4aNAKPC+IMAnl4916IP6UJNYcQj2sC1X
GCSXJvc2dTaoBXSYwRRDLKMckW3AIul9Fp2uRRsMCg0Q1raCakHRHWOS/WL3fUWO+wl38iJnCV18
7npMf5PLpw4karCVx46BZvAJrMKPbbsQFQOkfqut5cy1Xo8Z6c9Yoy7FobDB/d62K5r7lGG3L1ta
0PpUOdlBR4F9Lt0ODyzsUp9+uITZYyQJhSP5cTu4wWUA9ebn1yM2u1/o7Ls29rsILs8GiLWfbNOH
SsX1kWQ5tiK2nLzPYywOrey44l9omjqVKoRwKI+xpjceH0YRKCpJqNBONiIEKbKRsko4qYE72Z3j
Q0MpkbQ8XwE7fjFz65UnWSZbjarKN38XdxYCDucEbsd3vW34NJtAlKtun84lE3++paHIpf52a4X9
mOVHebP5Y627dcyKk9krnTfFdljS+zxiGFkxIRnKbPjR2pJDe+HnI9KOdpoOOguJqsHGAcMX8duZ
ahZt1fJVw9SE/gx0bXpWA+THLYAm2TBD7lLaPQoRPtPWbnp2BQ+xUk199Q/u8YAFCHNNw7CM/JVS
AhMWGnml1IIxaB+Qq65w7tVeNs/kblCCTpj73BobuSa/MJAJj+ALXsqmrtC5I+gIi1r8V3DYqzQu
IJNXh+jXkf/npqu8YD/LSqZO+Fi+8tyHBzsu9ziTxXC/LjH66u64M2VCSFIdMBU1qp55P+9oyqn4
VC7xn/sb6d0NbsEep55+8E0S+r8rGXOjOLphvWT0p+cBuA4ZFZr4YxCp/CLcBLfuJ0KmXH0uVML0
Fm/Q0qQJHo2TExYeBvd8neA5Uuek2LtGbwN1uzf/ESevjv9N7lFN6XxpG0F3FyqNTnlxXLjqGVgn
7tdyHxHkX4K9ybLnpbf1kdHWkEzMvo2+BeP05jI/oksjotQTYDkXAqN3uyOX6efXcsopphq0FWUC
ENiaJBV6pNlMgYwiTTZdE1QA9pfUcbA6ecwtcfEH3KWkyJoR56NwfXeqRY0NcHtPgdDbcnIr/ZkC
PzmHeoPPZiGMtzcdVoYBX9KQVz2A3NaMhta8SZWYGq9yPzOuHNNB099bUYsXKRXPt/fbB7Z3CZTT
1t962rJ/4Y8ZUHrfmQHzeuL48++KOsNzm6iRSmLOSEyt9/3uydCFgCJnANFjd9T3HnMPiOIgKgW1
fzysKx8H+w8miiVhM2+s2C8Lk5ELNV+SBfmR1cdD5oyMmVLNdsf+15HZEY5rRzhjmr1T5h/Jbbzc
iMRncYHQA7923nkAYFjvn0YenM7RDZ0Qx2NJtyVh0qiKoJxPcSAHaWeehlCS/b5l310h4LH9rDCl
UmG4LGVUio4qB4YP+5OZuizoTuUiFy5PtYQLnlFy53051c8BgIRdFhmbZli2snBm3maLnQwUtjW1
goXg+GCs31JuAQbB6v4DpidTARrPDozpSvYUaprewN+lQeWX2yxk/Fb1OcoVNKMcizl2W8pTPB7K
aZiAWLQv6QHSlimuMG6D0kcpaHHeAxWxtA0fGgpBJk70N78ZzkVGDxowBs+Bk4TB5/187fu88d3h
b2oU9Z6A5QhW8Xsh6TmXS96epIFLuR4xdyUkLlT6w/ZlphGy0tRMCmLMNehG6lxJ0uJxDmXFz+Jj
OTYg/FzKwu8e01MAqmCPSQkt9yyzfXIPUg4wWr8JmOHOCz2aOwB5yb8Em4yA/yVBDdb4qp2iZBiT
S5c1nhNCzTDzwCvRqr3D1JSWUaVs7/DYIFYKgW4HX4kS8dKtqmh0Th1MZH5Edb4b//zWPzGjhTje
A+KmtV6Zci6rtOfd1oKdyc3DHVIVoKZwA/h3H4PuKYQMZ0+OWBe5cLi799dNItol6FmOpG8SAem6
uFOAJ4Ckt/SqZ8kuvai47j6oq4+LQ98/4pAw23P6OO42ln9ZqVnjW4+/vrGSdnCJ0PLukanBSivf
7ZwckunUaEXToDoTApCOYEelU9D3DZEYvGcP7UYBIbuc5TwFB2cOG4b5kryj/czhMFBjc+N/8UH0
se7MQ3hRCqeiPZT+WDi/vrHSdbkFVwflHzqTSmi8vzDDesc5bI5TPKDfzdtb/VSq/gzjNDjk1MsP
4kdz1f7rq/wDguzk3WjwbJdrM4caKVmnjDf4tCAxJa4SLw1sk6ZiwR8dVs6FT4tW279mcS69psgg
z6ReMEHXLehcQp8AoZ091UwU2aaR9rTNDbSXqgnWp4tGBL3R6ZYvEO1xxK0Ot1UIERXZkpij+j4g
WyyHcqYNLM/x/zz2tbmzA43FlBODwDnhBeHSdljdCA91B+0K/EI6qC85ggmOqVjHnbmYTzSLqwiw
syfandG/y++lMgC6qVM1uei6Ne/loRpxsh6SEWQsM+SKevTZD3jKgEWwpjzNJ1yHCGuPE8heTfw9
O84pZj1wDZ/X7KO3a3p1QVl/6jKc0lHVM2gqoCeDAvdHpwPF0Chm76deIEMjiGyG6Nvd92x6U6J/
NqvlTvUxQ/wlVuBwVMc4YOZxlttiTnc5vxZp6whhMW5uEAkDH06HtaPaTgwcGyS3pTyQ8l7JggFs
U25vi5ONHyxXNWEFVD1NS+kKY3l/3CCv2N1+gM6nSzjZXqc07WSJcpmA36YaaFM0g4UhJkB+jBge
GBIL3xvr4LDxCodqPpiaVjYND0rh49tZeDUb2pkotvm74860e6W6TG/E4aVipw6iX4MnMxPQeGzk
+UOsKIIVzrlJhvm+490MEalbQ1OV/DMQWQpMLnuqTj2unvbXKNiUY5pUAWEph6ha0MVttG0XBdWa
Bk2f0AQ/tmjYJOD7JFdjGTF0takOR/j6ZoPKOpGvsrJvi75v02FtoJmhf7PvdXr/RDCeIPPhnaEA
X/tFtf8Nj2cc2qzfkmP5v4POHVWI2GT1SAhegBq5g9dPQQOY0mnZRs7/WnMhbP38cVbyxcyc9mAw
mQU2qObCHlrZxFZkjMzrLUTc9CIBbD1hnwCLjVO8mI8kx7Ek+QIKZewx40KN+L19Jd9UzY7OYMKl
OuI4SP6Jz7gbl9/OSI34vl+q5Mp7LjUdXoOd4NhXUhGJDvEmv2s2JsSeVA59TStNDOCsRgLTkrHi
n3KBHKcDXmdYy92vFIZwiT7oOm6ZzAT3zw41degj+Ontg7CF/Cjko6n/LKyCdJsMRQQzGiUj+dGd
RbjA6XLJuCOvGlTwFf8JItu03uxDnSpXdn2OH4GdjPQC5PpCGybcXImEdNLKePLFH08N6Psjcsrm
2d+TzTDMphqUx3L1j2Yy6ga/3ZLIqaV/rtsMpcv6rZQn38MuRH+NKbftQOmb0bVgY5ED0iN0Z6GX
lr2A1bPk+z1LK/CrS+k5AM9AgKUmizE/A703oiQcJjvbMEXLLXhZhkFnvAN+0M+cLoZrbvxvZ7Zu
oFf1C1OonKEFRf/GjdTO9oNCF+pUAlKXNfwL/syLp3dT8vfZHXOxkjiRyzuTbXuANiVxo8CbL9Uj
JNaTPwxOLp/5C7npqcj8A1j9cY8eFb7kjvF0sxsnftDm0CxpykVMF3Z+tF/VSwh3yf2TLc3XB/LL
T+o4HYj+1pJWs1ebT3jILmyULukgXTlF4PP9dRFg7vMlDe2ml7TokY9weOEzffm/z+vy03i5I5JV
lXXItC5eHIxPN1X129mbeOgGRH5/80v40KflAh5mTzhRLbo4HOkJFB6fAne7/WSxCQBFA5LF5aRK
WgI+3YgKPj4rDXnbZ7HKAEuQB+bHCUL2rcxtvFR7m50W97HP+9Bvi2bashc1FR7jdaDRv1S5Shqa
6kwz6vq50kCkZI3fiQnqXN1BQrZMCX9LbcTkEe6GsskT8yJafbHTvwga/jU8jvdt8ydzjRKHjWDf
xiUgWi5qvBhc6GYClWVQI5Yh26jNb3GK0+n8CBcuspfR/WxLzCYKggJJN1VmbhXcKfmktmEQl5CI
81pWQG/p3CFDKV9SGU+aYZeMau0AZ9a0CDYdowLKWg2kOl4MIGhIMRI97LhyUw+QtwOXieggiobA
L5NVhxGHPR0tVg8QyA7j9FYBnrGHcVA/WpfTlT57rmSs+KL3km9LYjs6VPT7+aDItK6jj76sVMvQ
ELJxrjUfdVL7WQTZgmMjWgkvlgkGyDEKPKOrpVNZUyIWh9I4PsYmufdIaM3q3RzIO80oks2vQp2a
K6liJpUbB7kTMGxuQjkxxhkBSNbKW5zha43QIBDgVaNxbpPMNdRQ3BRUMNwIm/6IrKROE+7UoUtg
xGKYJm/i8zEnN6XWHriJUZ50RlMPYQptykyB+Zjad4R4IBhAdQnyWBkEvk82+mP1wIC/8bV3tnqS
+EwWqfGSL2VvUu8ToQA/TuJNe0ExXbGm/Tn1vo3KPKDm4gGlISJ9YmW+XDOFiJ7eGAqAcU0Q1rU5
PQQ3uEM/6taR16PMippb4YC1HPepLLmG43VkPlaxsOP0hZ8JFf3r3Ndawo7HxDQNzZ3NlEfo9W65
gW8c/sHzms2rDdWtQxIGTrcP5EByKi/iGfxII9SYON2PSZQN+z/YMl4iLyuWOXzhINUiGStiMdu+
xbeO4L+3xP9tDhUK7S6Wg77K5Qzfj2ekDQFuVnuF5ouWjmfqDdEHZg5x+wHGfr4hcGq8xWpbi+C3
wJErsKTadyg9ErAirXAoShVFh8PAYcGJHbKVty045CpUxA9mHc5IAOVU6JuxLCRgXTU6aylMXhbH
6sDJJqNNhoaB/Q+pMjvsH4q46sP1X5qeUvP1VqUCCLCTY87THc4eQlqzsdTDXjNVEmPSX2mBiQNn
8EE5ZNKGgxExAAjPhOYBogEkPEEhvfN0ebSyZFi6odEuFlnx08xXGHQ9M8UAdvkuMjNYuw5woxoy
9cDABtr+a8ZRck0EaPU9ZGUKlprk1hsbJJPEyFf77nuPc3H1wPB6rzWrF/AlXp6QFDPmHC/J5JqT
Nvy6AcujP0xod9/QZPH0/8BW2w9xVHdm84XhHPU4wCylPXaKTrYzj+wfMEWwhDDTsbJ0LCwEyQ2P
ZqSlkIxy/5P/e+HjFakrurR5+UAIgqRzeFGCVv0YYrHUCg41Wi7ceYleE8CcNfjlOFK4v4sIB+lH
4U3VEcyDXzPWpQ36gdAV3yRS14T5ne8Yom/Ne1Li3zbPDjidkZ/VWBpWJ7BcdHG7ZJy0szYbdPp/
JCP6mR5lcJ32yuqErI+V10Rd/8Ig9s5vm2Nr3ZuM4E6vQIR0l639nhnHXat70OZmLkdRALVYsT2y
Dz9NBOQ+L7P8FEkT0+vWprkDregGGn+edrch0wudjWa96pkvbU+99DyYqSM5K85ixm+pTBnDHddU
o53pFgWg0fnBdqx3G/GzTcsjwt9FxHW0VJnU3Tbq93ccsOH+bdyfaysNsNgplMQg/F5GdBonkykq
C72Ss8xMk2GA2lMPtcYPTv20qqyIJvZZw/RZbyZ5K3qXYCwoFu5YBNCdtGnkqdRrh8RKbWbNMiwk
KQ976ifw13kFFHnGQ0VJ5wM7EVrjJGO0qI2oJLwBog1YV0ZFVwVRKsugkOKnNISd1JpXZPkzJv/U
69m0Kk5LcC7GQCmkKSRbeWrX9IxIbdCI0wqvEDIBc3jYV38dIhNu/AwmNVLFQqwfmGH93pgwOkW+
w0nUV8Te8vfjvqicdwKg+uvoIgLZvkEnJW243pgQxj8I643Mv4+Mb9ZjuMk8a1cHFtfa1ojQ7mk3
diW6Tc2ElHxruwuEUo+zjiPVY9Ztpz95+PkX/mMliz9GPouZWvXjJaZbauSCByS+pfbjC9BHwoEC
JTwykgviNJcda5od9L1KgtAurUc/M3B6va5ky+xwVkbLivKri1e6ZQC13kMtzRQLBeTdiThJ95UL
0StrD2OTVA5wE76Vjad/fm3M8B8Uge2dRQEs74rkwgSkLIOWuT2OYl8bacHrcDXreonBGbQ/WnHw
szt1pdJJD4fsJdBeeDCbsJHwcjc6bHhq+r+dN6+wRMZ2o9niKpXTTS1a8pfH3Xd8NCqNqExuuG7A
ufLjIlVvBPrtk1XrnORAR5g3Z+jYN3u8aWICpberDUCcW5GI1IHOX4opu/Bm+u8akd0sru9TvVr2
9MVgOFk6ffNUV3U3ROiqzfLvoDTTrG/NSDKOI7dhHBeTwrTmnQD5XjXWZSM9j2f7FibkYh45j19K
OiAOARX065I0BQI7YjIv+sAU0ngfmH3gNksRLiWJ+vpbql7yFepsBsviLSFljZXcL7dA+sFWjcWz
lTED/vD3ERLZr95fiEZ14GxbBN1y07t0l1huLikSFHjT/jPFdMqBubqxmHrQsHVyuCwwcuCaK5a2
JmRlcu+gUMa5ZEcSHnzx3/CeBJp7hZ/Umf22HJlz1xdGNWTZYVChsTKUXpTDzR0FfNoREvpFTr4a
VBQKdw0byipoUmBAfhH36sUL8jgZ8m/AOe+clYHm5LmXcJTIeoxgbMzJ48Mh80UfHT2TTKjxWtAb
e3sWGgz1yFQ3TrAY7N8SZCNeQ8H1yWca7qFsSQ21sTlkSmY1uGt/JpW/zjTAJ7ySQMJdG/EDZWib
z5QpPuZpUpqRT59W/A6Pk+M2G4RvLOKGW2tVMjseVVnByBKbHrDYFo6QMTYJgN8dEkhOkemKeTQu
0BBlD59CVvW+FqDdxGatnJkPx0jJqJaoUTbP1AhlK6l0L1/J1QAsH+RRhsrzuaV7nzUVykqFTAeH
fJFq6tReknOxPFYnyuGofhBIqgpW7/35u9T0aQ7TTji5ilypiDg8zCxRhqJLwBwbjhczIaGwiFx0
ci36Rl9JicYHS483ACbQ+0msnQSb6tSeSx1k7kmcBhVF2II8axOBco6/xLrRQWD3fd60ZTwXgZoa
aQQuVTuBHm8xPERJusyGV/FCJDtVj8U15XIW07aWA8kPkBVZM9d+tAm4HKi9zY8ge4xowxTWPjTj
nd6dgUPAGBSqb9K1axiQa/KD/6j/9Fbjg27YTXFdvg0cQjUi+y3PJ94QdhxLW/ocQdNbgcVENUUT
Zhz7mj68voD+GeMkc6I/tfwmuJSybDBcpNmtlkMFNAyjXjkX37ABDjXAUhkXsQgb33N8AKZWIV2C
LdURg8XHJawyhBMyiP2eEdsIPndLcSIFsrPbxaqh0dSV48oWyLzmnnRyf+J0Z0dK8L5/gjcf5gdZ
wjrYRaVM1uHJhbwnY+onPuh4xp4480XSD4nHIOEfxDnqy0KnbhFFgFrjrXxbsCNyJ4xAooaHCQNG
TfxhUrZ3mYFgXiy6NVX0CJ+898tMLnCX/JqyhiK9AIRW32mH3kt0NFrZzOIPTlQZpLVcZv/D/4rL
oBXRqFNiqeTJ5mqEDvMthgV1KSUveQllPIaozeJSJZNHNd42Ogx/1m2D3yo/3eOo/qz0C7MyMbSM
40EZ9v7qz5cchC0eCAWDlhWaH6vds5emRe/NaN14zd6huTJd+v7/bD9GCYQLMFo0K/oHmUtV8Sja
OpdhWko0KdizII5M2Fw9N7J56YOejeuTyk+BvoqOr8dECz71SbAw/s5X7CD384GPHG8DO9yRh/tn
SBaO/qjkKn8fl4qs/6UPU7kw7u4r3B7q1+WzQAgypephAtmfYcHsCuOaIGIHKfSYcsJRBN+jQzsL
9ewJSWR4V3ZM5lx20elVBcBpQfifxlTWf6boCIlqj1qLjTqUHFt5thyOCQSym0ZHL6vcS36paV/C
BZI7HZ9LarBalvA7QWeruXHRCh6Xo6r2QUqeSOm0dZW5hGP064C09n642RFE7O8+7TzrrMGEleas
VCu4lYcKWmgWLBSCesR4+dzhX+sICLWhPTW4rSBZ6tqmbjK27/uDhwFfsi/RRAZKJyEjwHcHmOb+
cNU7DbOxl7Ow1JGM+CpbcWtMPh/55vlYrXHGRNphJTmuNyHyjZrHXjrU2xH+PJc3fCocLQU/V22H
M5vb7RCIizj7A6ktEg8A8UwARmRUhmfVbwREpg56UayXuywtaUdnCPVwq2SWtCGlWB9p0qk5UWFo
jBgDuaR2Tlbwo81HxIyR+BP4+uBt/EARJ6fzDne/eYVaKanETichI7zEiOWCpy4NgHhfz+KgtZRe
nqs4zHoL3chtmVvj+jHTeQNjCWIiflqRkt/X2vDCStnWH+RLxzI3i+joLo17CER3Wl6zj85uMMSj
nzpxOiE4zuHkmCfKG7XO6H4cLx3BCKXrzPrjVSjgcqiB40XKh61+yb6EQbU0Pt6aEhJbx4XMO5qg
GNWwfg/+KcqFasNkgXdvdyrf0joCwFylkeQ08UZTt7VgxAVo5nMsZwvnfc5o7vlVMSbGml7NqSZN
u7JvUBeZkHwjuuCqwsD1HJf4hFO9lI49TeQtomzjSwMRXSaK/LYQqBQvH6azKd974U1bK1dnfvFI
pbgKpTDwkGOu2IjhmSESbXjjWXHINYOcLwIT3vO68H7/pDbNJa2T9S5Y4IGvRWbIJlkaJqUGTwQc
0RlPKvWKevYqX3oVGgsY8uf2RGdQkuDwOeg+xProyw0pyGcJ6cw5KyLBeOEeS9zptFB+wgih2ZGe
BsyA++tCXDGth/uCJZYFTXz1uKXtaEYKGHDt7PdZEp8qYRSs6H657vAJXIUUtiXnFpbb9LsjCf2Z
zRilj6OU//OkhYRyY8ITyPLytpPC96RnJcxxUMpKGZ4zED4r7tuCLGt515fA2JtW1GSZFYh4JXRb
gFh08SZMd4o98pjooFZhpbp1NTT1csScKHj1UqZufdCN7+bCsydZYiOnDsJBeJsJKTR5tdQlxAFP
q+XA9gb/BalBzRVdRsrLuGJHdmhgEu1Zbpn4BVyovb4qIznlpZ1+Xc1p/3/TA51drar5T/1bM+Lp
B3ojTB+aXH+1qjVgIgDn2WpZit5b1XhGH73cr1x5deXpWBy+1wiYukyoNQgqfbb4RPX2BDcCNaUs
Pqg0uOMW7mBbBMZyZ7NggW6hFTqJ99yC2Cr71faYRPgDcyBrBiuua9BhOUIhc7dRD5eRphHUhgBR
tcGA3CvX0l1EGIqDZ/hr4qceNXV0xxPCith1Wa0dAFlLvmVklNpoYGzKNY0gxKUZbVHyEtsgSM2H
b9MNXOdNm8TTyjbv7tEnVaDQTAuVj2LpK+ZhbmeEE+xyYNzRBk2eLYhOYCH3ElNXFCs7mmTK8NMs
pYdG6Id8q2zYtPg4ESqvUk1JFVgHlY5nVHvfavvwt5vCgho6bFR/h97Mv6fgQBE8neWqxPMimA9k
Nkmpl+03a2wUV8LOP2D781e46HpCNphEs5nv4W4Y4J5uAwd1NHrTU5STzuIylNYajdVVPH7fniwU
hiBeobSkKEvJJXYduHWdDe72ILO+xj7ACeVusixtcyLTMW4ee3lNYrP7wrBPzn3F3Llx+UAoXXQD
wG6FoyHujWvNZU9IipggQRYpFa2aQoq7e5da0IZPbJ5s8CRmb2YW1KUepZgojil83jMjf7eYKQwS
bazKtPBWRnNpVryyM+O1OXf3xn6FlqzZL8iYLo/iZZvhvBehDHCjDCDm3sYsmz1cnY3nb4oOEsR8
6O3OJWYzkVXB5Olz+XIgc1NjUUMFcyfYKWF7qRcCLpvtLkC41eXkUGwbPO1/GeYKlIZdNkwyrWI0
wAmxZTB/zM7JN2yyrscxiLYSP+Dz6XNweR4F9jRQ6qiLyoQshtHEOXRJXPZh2XNsL3UTukymijy6
CioZVUWPhDN93M4iaFMUk+GPyPpRGa4qjVYbphUxG9etzLLsytArvZNRBidfeNGfdtZmdk09YZ0g
vxs+SHj4e3lCCeoKGYod7MXEQtb6l4u1/51/DpVEPIST9fhAFxn5diLdzHHxp1F0flKELP25uUPL
5nLDMJpRAuj/bhV+/Txx7HCCUIG0jExn+AySV4FzlKhNtm3EsyTJiJ3Vbq+vafN0Lu4Ztivx4z5e
DYfHEmGJXpzEIfC0w/uwJLxmN3FnuMUqHdlbC7APYYo/tNqdhwmnuFIBvOqlR17cKhA6mwXNrx/2
ftDksGhV0rMbwOZOST2VxUJ9BAn3MEvcaCjAQ1xHJlrFtnQjWKCl+FwGdlvpX95MSEGaX/s3e3gX
+A4LpRufIA4iVQTX1hMWDiXZfPELsXQibdm+U2zLdXkNIWIkMJRjVWa0749mB8UecwgUnpTLn70A
bShu5jiMFMGe+s9snIv1pR/7PeW+j91UcQkQyn3STEgdN3EQyq3SWJm6jS6j1mp02YeRYrIcnPYQ
LA2tsLzEHeQhWAnDtThnlEzOIDAJBw9ZadGwMnuSx8+GPwmirdwleCCMDQ+TCRAkR/2q3UVM270r
nh8Sil3/P5ZEU6jMOHG3I9k8fSgQKSyWXTfnKiobSoEo+LbrazYeFE3+TPzvIqb58sAOKxP4y1fr
6uOy7pYuKdJ0Ay8FHCAWuzGhex1fAf9qEttRxVSFqPdbbCFQ6+4e6JqKiLeqZZQOvIcpNK+DK/a9
Xl7pDmPEE1/43ZMN2ZjYXFXqHgeZW2ZS4MwB97/w4jnbIBUnVhADngMWkQHKzyubrMnvtqq2K9hN
lgkpXmtgOiZFq/vm0ZQ+D5Vb7gL9ORPNfBK+TPoWbjdQcpomGrL2cZ0GtnuhkPSzZBeY5T1hLooZ
zd/b/fjd/f5PFpDiceETy/DUO4j5UiUCNqmAj+cO0cY90y5eo6yDrjrWsv1+ujVCVA22X6RlQGNq
jzGOmTWsv87birrRVpneeLXEqHvFUdeHSCGv/kWVN9PV0r+KUgMOL8tQ1DgV1zyvax9cfx/aBViN
JP610kepEHzIo9H6Gp6Ws69wpg3hCnGQ5vV8lQMutTQSGXZbOnbDCHopAvI=
`protect end_protected
