`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
cuciLzARyO0S0/hD7aRTvmBoCLwFffcj8eTXzo6vgIJs6pHUp8jCvcnQU2C8C8HNyFdFNDcAYRpp
aKTr7oC5mw==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D8Aw4HbouZqClwMiAK/Mk19vsrFb6Ep6CgF0Z+tYuO90CwJECvowYkm0fAbx8jomhtphTlWKfXXN
1+g/17Odke43WrGtOS9TVlHjO8VsFTiBJbt4h2rFjXKOp4fQo+2U+ICj6NcQq6prIrf0lMm70yel
ih11mNSzs7ItA2Q9LTk=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IMLWgfeM7cnrMvR0t9ML1z92jl9LN9oMKu19bvy0xHnVuMKLvQKi6rGjNHsXiOEk2jFPJAc1jxNi
JTdPNh7h/EaJZ1/+ybSggpewZRBbE5nYSZB4r9/ZIFbioNwtFVkptGreZaDpnIVoJriDk4gSDqaN
gAuHEmK6yKdAhGxyXNzyeT+azHnKWg4Bz7c2zsr7IAaEoLKAJ8xumCpayJbSpyGY/7V3y/hyfBcm
ONb4xgoDbpID7lyJnT1aqCwOey4j+Gh65kXJ8d4srrzgaeU6w4vgVIzhzmrPChHy+1+iaxdKPpKD
tzapzt+3LM11yPCuqPRzJXsGb8i3aLIU5tJRZA==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
TB5W6CGk0lXOLlzl5t2B6GJRYbMr/l/pK7K3V4fZ4JF99lGL/Yt10EGBF2Bhn7Q6KoJN6u+WBMhs
Tk3e85EO9sUQoLV38uQ+RLfyAsy8a5e9ddrKe7ORfD73BEbl6kcrZ9kmM3EGA+pj/O2PPwZ6biLe
CsOsYsoK8WAOB95K6uHUtwdxNLVUhMNgsu23mLzb4q8JfN5TO1P/VHgllV0xEZzdokwMMpFtfs21
gCL0AYLfl6zgarP0cqkt9ZG2oZD3iNdpugXvJnIn1N+V3IXPU50noKBffFWL5/m14Vrfw540oNOu
2WE8dTbNNui1RNwWGs/7NbnqzkTYqoULjtItTA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Vloq9RMe2+FUeZofyvLTiOPwyx6xcz0OT2sXCoL+ShOit2ZV8kYEi6nK4cJHljDqyAWMYHWI38f2
dPJA+xCpgW2X1GaZ9lpzeTNjHGU5WC+ajKAN5TaR/d71x1luyHmuF+Ol8ofBwv9kkkq38Yepcu/P
lKEYCqpZEIafYGjf33fOZyssigxG3yyJuDsDIxSmwtt8RAma06W8oG76QUX/43ySeqSK33ir9e6O
9ecb5Ozd2z9/VT3s+Jkfg0ig3mnGOZ2srVIR+AdZLIgDQOaTRYAq3soHd/FNv5Ylkc5T0+U/qhW2
v2O7mdgF1mvh7DqlYyobGYf8/Oy30xjYHIZIYA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
U+4HB+45CXXCQ/Qo8e+pRCfNNUAe5tIeyAGDWOB8P2mW6XdN0rzJfs2QI0dZGzWQXO1x7Hi4+Y6C
feShSDo1CgGBuBy60i7Lh3Hf6VX7HhYOtXa8vL629jkbywVSV2rnKzIxU1OA88GHLP6fY/gFew8D
r3cPBjr9CGa6sTyIDck=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V1s6ZKzW+YeNkF2Dr/ksBClaYc+iELPMA4bhgFWMo0tXDixj2mbXvEpJr9bkGiu00Ff8xwdDYd9P
wsJycbL8o0y1nst3R5itErxRFVGnHiAexe8dmHRrPQyzF+gHpZRCVuBbKVcAL96zWlEelF9HHxv7
hwdw9pi4kiaxQ6p6ZH98Hi4TRXrtQzwhO8k3ClDgb2oiLA8uRs0q8oiJVUveLF/9JWY4o+vKCOFe
3JqVphINQeC+H2tpb6fT97/N71HSkjakDoVyDYNF4Vd/r/EXH0Gzu6yj5fmy3GydcHhfjUsyyfX1
KIidAvpYtS+vzz6jSt6RbFt8KTRio2guFC2K6Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 60576)
`protect data_block
8ZEPPW7gLkpFE9QdJP9dXwz+y+0YXp0T1psxUCjRzmfxTS2G9sJpOZWF8hoSbADZ2HtmsKZzzbm3
bbzMNFlgPjxw7p5pbW86RN638XsT8quL5uU63sMDaKbdnlUbU5s2Z4OFWGtWL7d0pGr0WSdqmKex
7moWFmxwokDlYChtzsPvi6au0SGE+OmDws0YcdtY0/QPpQrtshb8ipM5XmA8mNUNcUNvkgbysMMY
bsjuax1+96coIlfbat7pAHbfvKH4jSKm9U+iGSpWbunhVclEBZGQ/7NcM1CeLQomdMMUkmUThjea
ffh9FBeEkr9MV2cslRScvr13r3CISwHdoJTm+0Q+8gpgHNBdPSS8k3BKYLUYenW8P1H7T0BnR7CL
9SmjLm4ZhFQZKaXrgtcm2IsJmXJPqJbXYtidRWG9yv1/Q4TBxARoZdD8bXD/pI4ZN+nhWj9vLliU
/saquaRjmQi+elHmA7XxYaDAoI48SYFvi0WBMEEFnn+GvFMErw9T9Q5wQna2hb28UcUMb6hAWe6L
BG9X3Up/MDBQKI+d7IWPDLjPyIaros7BxntZcr8Brw5ie24Bza3H40KtjAl64FJX8CJu6rnSvm2Z
FKgRukroIzMhC2C8zgtuB9xqrbUgBdqh/buMRe07k4OcpmQAZxXucoNyGT6wpp0yU/NIXGBDB+tW
XFK1iM6nsQalhLZ2c//i9zz0qJkgWPNk60KFUsM1bQhVd/zmPZw5sF6eedW4SJ+mrjBi0maGMDot
15bXAYy4D0ylERGi0GJ/bFNV6ojGCilXdWbEgvyRRVtPqr2DIAQPbvNYeMlO3thRf0g70cCTux02
ypC64gp688VuiHdmWGImuyie3e1FA+/re2WIqD+CgWymU83lJ/LibdheNUg1k0FqM6c0UxbM5hTL
HrYe3UESP4gv3vpCUNAwQQaBp18Xx8q2Ntpma0LWAJ04Drn1Th3oWCmcyZ/tAGkBXPDfArG/f6YU
YMOA56VtgUXm4XM7MPCIpcHp2LZWZ5Mij3ef9dPJRGIWGc48i30thoO4mACBsRjt9YUfAMtXjImk
uZfh6cXBStD6VuO/T3Bcp3Uf4eWXMbfFY4/jocORyCfsZNCKNLEchxgdpOBg+FppnPeIqJ7HdzOn
0x04DbzpkKpRJMGhtSs2SG+bIFY/Ic790JWJ7y/pZKnix/ePJ+JSkrbbTsfRvdXYvfIaKMHLJetM
e3rloV9zJHD1rPbdQgNlIet+gQbUW7IqC2gPb5yc8MCvxTYmpitnqw3ZK8wCf0OeeLK0XwzaJv2C
6bYTyDpwJ/3nuwA4wZHI0SLpU0hTPrGbizMrc79M5TFc9mdQWOaBJXenhCXbZ6wOiBAe0eCYkPI4
hZcAqOdtUJDTCznkTiqWPsof0/EWLigTiXJKS66lHBOhVS6OjKMKHasGFIj50cYsr0z9wT9N0DcL
5xsa4PI50LVXsKbuvdI4/hjpLe2eX57Mwyc2bur0C9w1GnzgbngKdDK4Yk7ivJV44Ug6f3uKjuM8
RIqkQQYW8LrEwFgLr2TkEHSmqhqW4QG0e1W5u42ebKkIZV4CoXaL0KacgWka4aRGlSN930HzMCmL
BKmWUFp2y/YvHB2svk0oDoUqoSAIr/I3/n+8GcRRNTjhMjWuamhrZZXjRlY9qRn2j7rhgCfCwHOT
iwJXMODcmN1xVAOcXRoWWOFWZfv2oBt0iO083jHSKurwz0VbBP+PLYCXb0zKiL/NPgVTVI7xQL7i
80AYFYg1qcI2+9ExlfwSi7pUj3FerRTbbihyGzFGjeYfO3sQeTNIWtatx6PfBvbk1COpzx9+F1th
L+NEPBNAxXp3zXZPhWnjlX0p2nHaETzDLjCpaDczE+nVmyxC7sgG1IMkjl4+4Y/eaH4rUv3wug3f
Jmc1jnlSErCvHuL0noqJJrX58q49p0LUm7CctYzzEeifyrQ7cFgoVVTeeeCjXQRUNpzuhRt/Oq+/
btRZoqcGc2j/Oepa5XCbF2On6848/BazJntaKxW1SlOZKSGebG4mldjvuuBLfZUNnHtM/RznzRhR
EM5AsR7kan8odqpilQ8B4lbyS57tn/iv3MtUJ6P0O9dg4Ha1rYoB5PEAJ1/r4L/pTQUEr460Rbj4
QvFiDy/kI7HkKn67TWXSQsrzQWuveJCwf8+xiegolCLlevv+yav/c8A+sPNyJ+dlGR2gfgO4w4he
n9XgMUtl07bVunktmdqWCr0bVuH5De38XB7qLGhGX6HLAXXEIAulQvlYSu9Re58mWRmBqXa1G9Wk
4468requ0yHiFZ8A1VZU+BVFp8ftLzz8nJCvdaXqEB3vZ2c/4Z0WvGNDYh5vAU/1BIbPzm62kFz0
gtpjAZkkKQZd+CjD/eU54UtmbTsn2spEkQBppABeFL7DXtkIMI8XTZvgqGugM29tM4caOGK6H0Ia
MHKvXFDvw8VnKjzrplBQH3MZ8dctGQlyE5uUN9Y9H5mWLSlTbnV1z89TfFAaT8kc6FZvTREsjC6Z
FsEO02SmXu0yY+j5iR8fW2iXy68uEUJUQ20Z5S4Kc2U4T9OJ3UAtrxz+VQNQgB52ebvLJLAKHabg
Sv1Hh7koBI9htF6ALbyweTk/wHE5U1NupkK8gxCyWJjpg/oZZJy/x73Qw6hr5Fx984FkzEIXSNz8
eK2YzQGzaUDYE/V99MAJhAsx3x1mQYiItIVItrwK8CsWAL6/820wbTTQhRk0mXk6DKXPR8i8+5UH
Ei0bRGXnUM/kOWgMcYsEbiynLMTBmKVDLKTem2fh7hl4VpWJApnR8+TGeQcNyRZzbAgS27HrQ+1i
iLpGZpHZXwpFpGuADraAkLbrks4GYLtGTyQaQnLA8ss8W7uf6Xg1YYc9nd5aDK21g8pnV7BBwKGD
GnS/I4pnctOHIpcxjfoBkVsKqo5n0Y3RH76kB4bCiHoG5cTc72ZRdCK+i5anxfKbFH9WKy6xHBlA
9tGT1dqX5VMz3Q54e8xlNFNc4ZIyng6S6neohsm5JrvlM5mVyW6aklpzSXujaHH3Aqx9Gb0MvLnx
Z0OAsxs9DOzG1iJKs2oNkqeVpOip4wLo5zq5UktSror9TKL/tWJcf/HRd6lCrJoCtGyrtLQMggZw
OHlOLqAxuAloRumhHOMGVmuS40WXxzD2SlvNksgzFNXn/i4U1icizNo2rQdcyE2WZwDzFfvkDh//
JwyfyBSfu1zJZCwMNZaslV1ACwNfj55t/zHQW6QWEMvbE1AWN34/OgOi3ZY4MuluFhEomLlA1Dpb
/Z9+v/K6NQHXP9+vEJaTHVws6sZuaooX78xIlW8vWcPyCpaP9i2iAw/Knt6Mmmj15Wfni9aGS8mi
R4OammJyoc6O2GAQTqWbwQ8Ogbl6GIeYjChz1qZ+wJcQaU5ZXS+R6kPqCx8DBDq9FS5y9sGgazj4
jiY/CCTWwfFLeWxxbT4cTCTtxgSfoOUfq6JVkCkHUH1i2EmzGMQVz5wnUiEs0lz8uEyhay80EGAo
qt5oEO4/f/2bsMRzVrUAvyhP+dEm5FQ5iCQQ60iaiyMwK8jvrQ5J5IwuOu7OtdhgRgg6d/NngKd8
BRfUFhF26rqdbE166TtHub1ZBCt7yUcz4vlX03a8jLfJuo4IFZZJdPuBGrZOkHwFkimRToIrvo1/
ITNU8SNHV3kXOgzGq5im1RHoX73FDgGR0UPVn+oi24e2eXHjL6uzdMiCFJgA4xjqp0JvFi0hOxGQ
Y/IIBvGlA0fBhoMnq9P7C4CPgcA10LqjwD1u2YiiFsTSYBkXCvBVD8h/xuk5OkET651GoNlYRUN/
0opwh0LHSs94Xtfz9h3OkrRPH4Ew03xVZECBKslnwO3HNzxReuZnJBWfZCk0MB0J6QIROPbKJ5j1
Ke6DtJLgY7Wehv1itgRfSa3PGfDGjHJnOxop0SISe6JqNPnSEe5GkKzHrDY8w2fPAYYblxhJV1Dw
rcG+QVd+i7Qx0o7I4rEZ0mfuVzyUrIz5Lv/1hWy2trXxxDMW8o4kJh+1WvQRFp2Ei6mLhvpJlbck
mcf7aSiC7y6ocR3CesitKKOO38fYg+5WulqAvWZWgj/nouVGLYff0C0CsSaGCowOiBpGyX+p1mQJ
OpEWbwU/Wp8tfyPP4rourNeVlXkgsukcBwFt3MfDaC/c6ajNO0pk4xDc6IVzqtYU2bnGJQzxYWAj
Oc/ePV8U4H5QbkObVvRQgKQUt71OlS6L8/D9gJMNrFBThJDAdDsg/gZFETNugrbnOuh8ovfRHRON
mEDMrmde/tpTMSxVcSqd+iAhVgXg3bVtrPAVeuIWbPrFAADbHp3AmGxcBLgjBzUa9j4ZqvMGKldX
cLcDpVwMJ4xpsd9YOcC4+Rr0TGzzG5KXDUsyId+2N/oKu8UCeOyviyErerrQoJpGY8ZlXyIQgQZm
iBmNnM5l2jo919TSbqMz5Zpf7AcnjK0Br4JecCqIQJm0fSKUDgoOJXMq/4UJKRIA1WydeJ2cBuQ5
lG0KTxF50vdvX6YHHplLqqI6cnNdgDvc+7Z+85e+eBBlb5DOH6XyyS0WUfNAenXDQI+R57q7J6dd
GpkRZvpHgJNZMi6TQRpzdntrW/Xfhqp8lZCCirCdc90dBEIbMyW++oS3+pI5GjwjaYsxttQLZanb
m6ExiwR4f+Pt0n6oEolYw8VHPQn6jjSSdYG5OBZmCfbgAYUim2+SXB0Fg8t7XdRIFFZeJMvABfMm
1zuUzbXmQr0OW8Gt0HTfnn/QC02DWsLzwbBUuOuPpqrAQIF15Pi8SabWUKRtnQ6OIVopVGLfUu2s
3yd00K15OgcYpdYba3Y7lXNovY29whizG+H0rNRNA3uC/M4YmUk0XAmw72rZ4iEhswgJxcbIT0tQ
JOtANrfbsg4gv4TiLFDkE7gP62HmLASf8nJmtQ0FDYLJdyUiBZfRettpLllOW4GQdLsGcwm/SXT0
uNAG7fWY9yzHjgP9NmzBCu6OaGLkqcGLqPM1RHTJyI1lXsflGwwbbyarkS8ddWoC3Raf1Rg6zUMu
S3XW1RuiJmLCYHEwez0XddXv/7CEKflvtG1XoHtqaFIwTmZ3L3EnWvaUrn7ZD+PHQInwxijJWvKe
T0T90cRkf339sgwn94p7GfKQngRiEYTDYTstZjmgDWqHYQmP4OZNKKmCvXFMCSeUz352crTBv0zC
D3fVTOeyvFBUE/eiY7EZxZM6y0+fmkT/be2qFkIxaN7QZhg/9EBguV3deu4jEr67oi9yiSxKjN5c
3rqU4zqzO5d03SWieK3HQ8PhTgTTj6bX0F6b72DAWZ9ZGxQdLBNz5qJiGt1Z5IighKyBeI3BRN0Q
5LPz/rxKUfHI7BtEUuKT3yImz0IFZ4EbUlk7AlBeUar7gvCO6qg38KdwppqrCEqRuLhoooNhGPdD
oeBylNWs+8QWq2aUQjEXZlLF1d06TznE/Wnmi0DDT6kgjvwZGBw5CVvuxgDlfe61wJAVdwIaKCLC
cG0D2itgxJd6v7iETzdNGYNjxgbjZirVu2T+OVvBaCxBRPZS9gB76J3VFYKwezB+rs6qYltDPJPF
VGP9qZPj51JN3Ldwact9GbamHS07vlCgfM9iedeDeyulEcWghkRoMNNv14/puBBfH7+pjzxFEA2s
XPbYFgRnx86a6xNLvcB+wgbHKDmhZzhjF+YB0fJQ65H0QgHj7kzzXKrWSeojHumuoxSVt6JWREVs
4l3oIo0C0rh5umiz3tknmAHRVh2K0hTj8C3yv2dS2ksiEi90fEfXVSjpO78eGNPmhRQgGMMW/ytV
v5GoUzAKE2MSQ8w+2RQiovfaLk4EaNKgSrG4Ybu7+1PAZr1UUTIYHJv+hg2GOZKEbRj64ippONFr
eihjzEkJAsZUMOrU68g5Gkr1sbeuu4aD/vD/1g2OCqMDoaSZ7BnGul57KRi346YIaki9X8v8bwiL
icCogfDTpW7ZNO2NXGbKuBTWhEDbNVh4mcXV9+dNVYcRywfaXogab/R08RjOH7+y4tWU0tJQgVpG
4g0QdBjpOjgL1uY7lFw6MdtGdL3aP/KnXTm1yYh+TyJnqJlz5yyAJqRXtOuYeIGRERd4xOOezVLS
YmS3oI4RhHfKEPJF8y9g9kpRZclzW85dmj7VMOXQ0v0XB24oORi996liTdkaEZ06TjpL4X/BJ97H
N7B/pFQdLkE3RIC5cwOGP27zshuNXaMEZDopkX3eSPKlBgJNLMWIBRVaebPvpnhDaCbWDtdziFvO
L78+BsU0RaaXATr1K0NxssS2FWTRy87IXexpatP/p4UzhZYnc90vVlS9NKAHOe26j71WkYN609d4
2ouTlYxPFNi/WGDPCOcltfKeBF4MXVWrgqlYFY9ibLj1lCxRWGDK7BByjVoM45iE1H66e6qQX7pm
n6u8XH4oqZuUdO0e8t7OVV+Ly4AAqn0ZqOi1Yblkc8HXj1+RmM1L8xD4YyPpz8+eB8AouuZCVmAJ
youk0D9Do/HUr4RQcQFUhAZ2SfEIVgqDUxGm99qwfS/17NbSItvEesM65R7wdj2WM3KNWds5PJZF
qzDwe9SfkzA9VKBHT+TjduEwZy3fy9p3ot84DYNls9B3cNSgNc8oRtd9FA4Cn3MZq6vTeZyD0HDq
7qCtIPAPgoQpa/obWTxg9IYh4ymH4t9UuIN7lSh239cm0/35TU1cQ7EPocafd4gDRaapC+E8gsVc
zXHH3GKGOECgOQVhiyvCBqI9fI0h0dCaNwsEKhbpxMBmeK81Y41mJa3psreyNbRlwMCcuDD/HdY+
wsPgutZcVu75IBT+d9FEhqn3omNLNO6MuEeTlVrD1EXHx/2Y+xWmpvN4SeJSY4O8BrYXeKCDziig
+LwUBRZqiyOuDH8iRwfUbiNS3muBZIujsgrVM2RH3+wj+14olQzMUTW1e3WRLsR9IXhBxUoBsrJy
aOS90ZOD98OiRJGAQHmk62U17K8Iqig726Qdn4lpX07PDaI1FqtJRApgRxlZuqNzcTSIciEFXOIG
6vB3YqhMCVeh8Of5qu1pjsyoIOf8X6J0az8CmjcKnkpw8NuFlqc1Ht/wrPybyYIRzRruKtKjhDu3
sazQAu5rum6tr0MGC4wxS5f7rkm1m4YQq5aIELcN5YpNg8OgRex/DZ2jrcpmkGKa3juz1magDQkc
z2PDEaJDRWNTywyHISAu/ivyPdBlMgWRTZDjONrX0sZgFfWeJ1YSuIWIm/1S7fLwUgm7iLOfyKLM
afw7TtQa0NFG9K+fiuZJWVRlsOoIUjorK4I6nNhE40RrkriYPN+LrXaE05a028ux/YlGJiPqo7Im
2zD0jJPpltzMhhfKw8hFof51bGbQAf9OVXBOHhnRs2oPMhEY8UKJs7JCSMUD560lThawpH5tIOcE
JlSylb/z9vToBx8o1mc80Bibvv7IDzMfbuXI4SwY0ukAduJFT4csitm6bkH8qzK7hb2scYKSjX1U
AI+RmisT9c/6P5pyMNhq6aTZk2MXzgWwg90jnAbOCHllgnQ9HLaXh7JzMDNaqasncVI2Fngx/vWe
TNBW54t5KWA50qxRH5PGLm4Kt2oh/UwcAR3NCis6rfhAyei6WhAelQZmt2z0eqk/y/vASxmvaiCX
wfxVf7ixRxA4FaDucEM1hlP/QkF1Qd6szDsguZeNoJ+EQmNSTWjbAhl58Cq2UsNCoQIHr5U0XoKG
lB0oBQadTxvuouhmU5wztzUrCkcXeLRPz/QPGT4C6Jrk4x0bAPshkm9YT2hHyZX3uTC+OkPImVeI
4yfG2rPMKUsogj8HpBYC0HolgmfPA7SHnjddkR6Ze2Ds/s8bghDBgLOt12GG+cvdZm30xVXQsR/O
bSRUGq18/mEJnqDfT5FCTKYSbE5cmJ4CnsclYndpfbr1XfDa35oe7q8LO0rzPV8/pBAde6508xwj
ucUNncFfh1BiEcHqnZN/c5pB3pTqH7VkEyUsFQcVXqiBh+7+LKQVNEqb3wR7Zh9Q0nhqiB9dz9Zj
oHhfKR3wA3cR/oUdhecMKC35o+cCR/EBvh+MNZwazj25GecyhLPCZb+y97N2bO7Pcxp9yc536bVy
dQAUheaVEl95hEhdTTK1R5IQgciW6FRjeqI01cq/2gu3xtoCa+GrP/kqcVO1P46k3Sxa4GmbAnft
3viN6U4FRtuI06FKgBPPyXWKSForoPFo9simY7OdmxTURsySqrO3mI5wdBSRC3I6QYV9awGd3Wvp
oHvfki/Guyjlf5zqAV7Mr4noR+hKkTmboRehOOH4IPtEYgCHb3gbDG44jVx3SRHmXmyv5wpfjlfa
fxo+leHuWVxK4s3rwdOkKIDvVaP2VTRHiV3o4bM2ll0rRS1afuIu69KFiNZwW2eTWEGxHxlvSgO9
q2mOEEW+jZs/Znsgd3Iwuprk0OUU3m1gxvfRcPW1QLhoDf5dU6HGOPCeecdREFLrAGKjUZKE2g0t
RWQvDlPC9xE2c9eZT03TpUXvMIW+9mAHw0zh0FBP8gSCfQ63wKenqiVLldFq2dqhyDzXzhIoC+Pq
4TwpDIeWTvuTgmcaAEWBASdoXTbPx4xQs1dcczElrJ1zu6y50y5NSQZRSUUCuN3klOMAyhBKArWB
TFDeiqP4cmB9D7SOb4eaQ4+QBDCW2b5px3SQ4p9Fb96BU+GDOdDQhd2HMrgwsYdj5hV2+QfRbAhE
O6WnCPWzT7kjirZW6QbfHT96VKDBwbv6pmF5Uw4PPq0FrGhn2ltB9hOv0jH48o7NsQzdcqt4oHyd
sdyBFFFIdoo0J8FTvRzHbGjbMAGbgxmaI3hgiWvI5iaUVA9/GFdd6dwiwV7lyGuIRs6SJNR3Be4k
IUbKZ3I6Kw4HN3SR6wL7GgkkSCCT3HpDfm0tXqOzs95hESHYa9eUF2VI2Y8kTMDMcCc9sqgvi1rb
opMD8vUVhu4uxAddW8x8VXVV5CF622hVPGZajlbkt43mNvbRkavRDb1hG+URqlyZvvv2cIp8LynU
uaRjmK6haRvUEhW5hZa5y3rEN8Gv+2eUhlpVdJKUpJmJrE8/Y/cxEY52PLZPw0nZI9TrDiL1Jqo+
phsOzcUySow0yPgfKHhboUKxxEbJVqM8J2XuA+lAiNsJ7qGjFgtkK5HREouKmYRmVEWTqtsXDVfp
c95rXOL7W0Cv4PZHTGdEDtGCvRIZwtLVjds81MC7jIIQuNN3HMcog1hj5U5oN0Jf3POi6LoLmB+t
crcGp/1wvig/MNyLGbznuGA42+WZu84p52T0OgSm1mgPpcMWRK8H+IAuegmaviTipsUiKrDM4jNw
CZ0rM4Y/Q2J2Y1yxA31M65wOA2Qv5kNA2kBf+5usLPpZJpRJSM7ZYOLkr51gLzbpXswG8sm7bJwj
PXb6Pc9bVNz6/pzm1Tf3nJYxkWi+Z4HUgc26oS1dxoC2oW0A+9IA9QlnyWcUEdLKdb5KJ3PBTCBC
yI2OBYBKTuFrx0tMUmJYmCe65bY0MdIxLGEsCb7RKxeJb96I+FYWLru7joUsWHqPBtx4uYIzqwgT
2GwylUsH8fr4fuaZMVui+hHO35xginE7MUNLP8rmoiZ1/gm9TR6LQur1Iacdwtcp9qVb/+1+GoDQ
9tzGSj6tZb9PYADZUpfs5vJ+R1USZzeIU7hC9+1ngVr7j9nMXY/h+Ps5Kil6/dzJn2bbn1vMUh4k
HDzEtY8APSxp6CoJ6238/0xnTjFe6MnCYMKmCQazD7RJt+vJeLQvDxcV+bKDJPl2xHDIx1mAdd1v
5PPqTvPGOpm5NEd1n8M9naqrrPmuod0BCmJCs8Ke6zVh1Va0YU/tr1HsY87QkxKp70SUWtC3SZB9
QGyJgJKm/IX1r3RYaSl5Q0r70JN6HwpqeK8gtaqt/3fK5224RSFbj0nk+QAcTcBMpLphaTJkIR6V
NnmHi+DgTV1BnocHLHNBwa0EtZAjfrt+x3uECCb12TUjK9q4ojtOtB7eDaG+yqSbtG1gwthItcBv
C7rBvmc9mT+EMiq/1MayMyi04zk8vq2c3X5ZRYAC5cB7r3b6VOkrPfsm7ZFgeUw+yl2+mJCnDw4E
QiRwXPCrNz8Z+3OzVHyYDg2WdYfakp1JeM/hU+xZsQjnU/WKxjTAC81b2x9KuFGrJGTqcF9N5RLW
L5Si+Yp7bJ8yJigjpfjuWIZmltEj0gwNLUz4mhkEoG79RMnJRvqcgQ1QnU73HNZPjjxkdzJPpWNY
iuSnDdgFBrXOzUTZODf0Mv1Wv/f7rpHqfN6tV1VC7cq3FWmQMyAGPqApQV2H7Ha/5qNAPd7753DC
E3O+3qrkuv4mt+HrlQXIPl0lWLWAdWxDra4BJibR8PtX50GmjX4PynZrVWelOxyGfpEGyoykAh3I
UPISB9uOfxDXpb0MLjA2nW6deJLVT5TtqAEuhGuO5ijFFMvSzsgdk7/F/Po+GH5V+P0icWsloCdq
PJ/UbxbUvlyAE+xPUldQlKvrQAuCmESJCqxJEg+rkQ2LoJDv3Rf+zypI7l/q7dYY+9Bpwcup8wgV
qlx6rXoUGwOBjFFSHOEJNtZ22Xtdn9osvERQOa/aUknFCkDGZkUkA9cNK0ORiXzZExv/YEb3Cb3L
IXLnh2YWJYqbUFOBm0jXOscU4GL1ERkEVOyM+I8z76STeQhZujLJ/keO/GtjGAZxeTyeCyOdWzMH
LkbtUnvmxfPoyelTlzPbQvDSkHwiklxvhID4everi++c0fyGKO0MjWzUHO9PfoeLyjUXvgLHMOuI
gRueAwl8+yHdryiIFxUx+qXhjZbJNIJl4mEaiCrYhrZTscHXhuwaWEC5cQBBq3hp7qMRm9ZCdHNK
iCTUhZYGhxPWvccEKwkQXykQ1qJozpNLixrJOzYk1DSzjopPawZTYei1NOz4JD1GrUJXPwLQuQMe
7U3df6cAdgw7n7yN/XK3mVzgyzHfQxhxQbidQ6Q1z9X0bsZf5Z7zmDVooyuw77Eq+SmaX7Lsacpj
TB6fU54btHp6MEzpUMpKnpTQcyKeoEeFiergI9gMgLo7v9SmsIjCyq4B3y/NrDvgbXedAM9K+i/e
d1q5JQhuyX32r6LotBseeV/lxGKofmXTVUHzG8AdN1ECWEpqC96jlCtB3MSjun4pEUFQlV/DYpLM
MQ7Vw+ZaNY1Dg5ELAKQUcyKtRChkS2qp4zYnGYnkXI0byZjrRHZW/g8IzxbTBlN7xMfh7EuxNt6u
Vhevmcya20lKH7ZDzAdLBEsFxXFcbclps/uIRgIAZEqec+TGVeDu/fAZt8J6vDhF/UGiox7Rc0lk
NT6FoM+Iocu7Sc36e8pgeRM1vmpO/EvCGiPDXl0Ne0okKy7Bhw/htvsIclPmR8yYJ/IC3tKR3bIs
WzOuCREXWqivGjHynwxZDq++8lM2QUbBn7rhfrY3elyAA4u8SfYb2jGJ1dyVnRe5TK7U0L1LSJvq
oa1aUpsrDu9ljz7mC0IojI53UE3dsC9hLrsd+xCjzheN0Arp6o1ItLZ6wOLzc6pMq1Z8aZeTSVKs
pGAeo5oiM4sJvdzKD51DChSDuGs7e8zwlckH/q8ToqhpwfzYdIu0TkjYtL7eTPjTLh2uqVFFpyTx
QQ168yxYikPbwnb+PMXREh6zKNcmWhheFNkxVE+DX5VutCblFy3Vee6yVnd48Y4cffDVjVrAkx+b
Cq61zgI9qfH76VDXlM5JceF8LMqDxFLvEWnDRCu62mli71pNaT3E+Nim4IqQRZXcYWylq5DLUj0r
ybQGLEbA1IsY1DQC8pF0mk2u4GYuviR4WDZC5VYtnio+6ISHurIE2Gx2LrCQDUaiV9wozRb+/gIw
V7AC7l4VYYhOGl7suectpv5FV/PYwsGWCz7Ur9b7rkUk1lwDYw0tsMfEP2NLSOWMnJCoUAaAU0oS
QwYgBBcJ/xYX4jeuVzGHB5Id9nQLJCY4GJzIokzT1dUmn2U3Eqy9Lmijx3Xqmk6OAXXmb/Yt7t5D
vWqAYV1Md6n+b2P4MxehOcGCvli0lOXpV4q26j/gQfMIFc6/avrsckg+ksKJzfdXpK+h6BpkNv+3
JMnd3UfNQG+3Lz8wn4Ri6+IPZYx2/OvRxKQuBnrqNoIV0xhmaF5uxWKDbnGhVaNcF4ig7gdQbaDF
PhSLyBk2Q8jAlZqCI8Qc/npfDoBfkHqGGOLKDOx/IlgE8o0YL5oNB7TjLxA8PZJRECaOWZl0gTlz
9QB+kWviV7WOasS0eqOSsn/AnqAi4m0swOkKEFhyZgMQ2RFQ3UIiwTLeBQ+9mY6KWkrIGai2ivFU
5Vp4xkWNvan2j0uFKIFEPWHocevEC3YB7gXqGzJ/6xQvgzdPimz394oW4ObzGaUumPQp/31HvATo
0gUcAE7IgyFwxdUrOd53d0vVHLUIcAHFB1KxRgKLyuSJnMAjRLGx1iU72ZLenyu7hpTtry6eHUwK
0+vNMdxw1dHQD+isaQ6Curb9rVsCIpzW7lc+f7Z/Nw9zsKkEipGsP8iJiY+KyK7E49/HhBg5HbGx
MBPGP4SjZwcHvZegZnw9u96qXXtTpqdfZI1kpe9G5WfYUK+kYQzmlLv87ZRJx1EtTprAl5de2GA9
lBsHusoENSWbSj1Slj8udW4oEZNnKh6j8hj8tF8Z1ZqyqKVmjD0iefuuMOKRc+6llGl0ryVq4KkK
liMZzsEDScxsp1d+ccuPjBgcpfq8QIvvIZY9DpDewNPItUq+Hpx5d/i0F/ZmNhy+i8G9n0+lcuVV
5xMZrFGyp0Mv5H4F9jXmjWVApMuqyeMZl9R+tczWxu42QkpjyzLURbvzMt3Vn+AjNxF3uGNq9Gtn
yaiEws9mOPy+rJ5X/bWBvayme2FUSHLd8i2bFTQGmrFgWaNQunqZsygZLajqBmBSk22qWinv7Gke
YGdZyKKCHv2mGx3BXYhi0mb2trEbCtZ0DVW5wxpb7NoXAxeWqwDhvtkTjjvC0kYYf07vkFO4Lrui
YjyPcU9yFkTk5EWbwtIsp9QdYOtd1vHrUYSCD50c+9WJ6TgfsbZhRjVefUznje9NPTsNQCKQEAFj
XeESsCIuD46SDbT3xY0wuBzYty68/bjWR1ekCq6Tqq+/g192P6mhFNIai4RdWkRhhxsIa7Q7vP2h
WacWHp10hy8QF34xTRDHiTZaGzBRZyPcmKnDzNGhmgRUDfdGAcsZxCPGE05pPrN1znEZXQVTnAne
5Hqj2xLbDv/m+5uHWTGXRAoHubRoZgz9x/Ybf5ZZ2TviKyBEYKv1bX3FbWsnWbwkGhSC2lpQSJ4J
/TWul4Df+binTxQ6Xkkl1i19R8n8y/jT420FIO7XML9zI+P0xL5QTfTulyddfEULl+FEsAVHtPOi
5z9u/g5fSDPqUxj9biOtkqK5rYh3N5ABLp9Q5rw08Y4oc9Lb0jBvUtBP9EMIlLDteX0yjOn4s9Xx
rLKyxJgsjB/vXP0MNsbKrYqpbJLMEcUXap1mjAlhUiV4B8QPtMaW5e9Y8xzQ0CYT+oYsRgkZyjbN
8V+5aiuh3d7CYiDdNo7j1HQkMjJST49p8CIPa40GdDv458UbW5YYUYJWVEtnQ/MVm1kPbHOuXDZc
is5ep0Z+1e9l4XFRhEwIqI+NDtAdaI5mml+d4+b+w78Kr8dy77XcSXBcm9uaMvMGTeYGTwiXwZV8
jv2kd4ic/a+j1LyxsH8d9MPm1sLBA0upHd4ZBRC50tqkAHqcmzROm+lpZe2eQheJkAFQjVVYeoGM
fsXF3SEKyuoK66ZzH8KSwzDiCyg7M2xqxxqgGh0MPbbFPJIFPSh434SmDeiIiVVTFxU7GwmbWFX0
WIy/sP0mYLJ17b8QpNwXaL3BlY1/MDIYfKOi5UchEJZe2SjH9wKOiqHI+WE1Oa/QRYWyUqE5yDeM
T6kPLI/6AsUAPPY0l7CukLx8OO/wCc7JDPzjzYIakaLrpQ22taSaReFzDrT22IN14LNIORe9pt4w
vFe0fDilytogkAWpgY3hYabn9Au8h7296TEljVfb1ts8iquQ8zPrHL5M0jm1fVULsaNvbcgi3UaX
61t2TjuCZLnQkBUjfn7zSUb90ybjg+4oBWFeMj13p32XMYzrhfbEYEATGs803dvyURxN19pDtvZQ
DoNsp2wpO/Gtgb7idI3WfHcWx5gztCAptLmmxYpZLFNLP+n4zm/mNy4PtK3zuzaJzG4maxCHOJBo
8Xlluf6PezzGYtfGY3kPBLvF5zug9rTpW4M75qZp7YrbnrxF8sERG4k869fyao6zyqwK+63mO1iO
AVE1uuQCcuVbqnNkmcd0dAau3pSFm9DxFr4Yf1yNef1hg+LQE7TZ4MQKQsZQjxXaqpWng7+ZtM7C
jxPAdZSE73yRTIKdWahnXwOp6czvZTwBlWZYSVwbMqibwMJk1nGqCN2Gdt2+y7SdzZILnqeJqAHU
ckmGXPmIE/uJF3DJqHlPSSwLmX0QNt4PKql0831LIwxNHlSvbBzWRO5TDL9SIHnmDNHOt+nThcFg
gYM6tkMaeseWdId5U4fNQCUV6tA9tFaPVk24QewcznZhbRe2HQ7BImZT30EbLPPr1wTDbMlIn8Bh
USyVoXTfiZeLZA3k8mWawKzSBtFGk+fYA6DDluGGgUsUN7EBj+wyZob5rGgkPQWM0tG46mBahdQO
VV9rHOKemj2ByBRYUI4FAY/hMoxCG8n/6nYZUSWAnU895hJe/leEsaLlposnFWOjmFD/ObX7SNOW
6VQr1X6uxKw1aAi4UAjzajsD+4r+5UJBIyoNJaikh/GA4hTvxpJTtVF60VcgKsSJyBzAecINRqUC
mCOzy6gUy13WXkb2H1vnHWgg4GcMykxiZQZt3p4qBCBxUAntRciF2hh2Ry+lqwrXzryzvbNdwZD7
cGaGkK+GV85FpnDfTcLRpLsfJ9m1SdLQPk2X1shVGd+gfO7aNUrQXxul1d3h4Aa4tmlKwICD1Mhk
SwSrYZHk5WXBUOC8nv1BBLjwYxzEPg0X7bOrsx0/OIj8f9x9LoZJPaAGeSM4Tj2grsDIpHtb5Y40
0YlQVCeXY60cCS91Eqc1Ek6KNDng+0Wy4lYMiPU4dQfNYRe9bNu77pN86WyMCoDlPiZk/CetcFNZ
RngodsiDxRkZeEd8QseG+sHrii8SMqrVGEKD/xG7V7d0osTaLX5dlvhxLGXAizgsoL0tu6NVAkHA
A9q62nipZIjsiloVuUj2T7PHDgp+9f58CeGXk4FLMMhVx4cweXaLOc0OW7YaGRZUvn4B+Me1XvE/
sj2K4H9rwQF/5eYFzSRorFJhRyt541K7+CQsBnf/6ZTFCctdvrDocfxx/c58oGbBCzYfafpAZbsh
dgG/xVP5mgHU3C0FdqmnivLj5PZasu7rzIovUeWsXRafRwWN410hvreNrbdZ6UAG99Mt1duZ8xKd
xCy1kex7qC29XWTHmIMBSMzXGV7KAxbYYdyap0RzFecl+eckjs1c20ge8pLBhGLR8SXuUPd/dP5e
mK40fGKFwjtySh87pTz0W6mHaD7meow9g87uj6Gy517QV64T4F0GWjNCxiKs5EeRpqso6DlXR7Bm
+zhj0mBIdpeBmjBJDCT5pIk/JYiDH6YX1CPL3gtGaZjX6Nn9qSvpcd8nw/tqQXjKkLOqvQ2mm9vm
0RY39pwdhqw3wQ0tqedaocCksXWfiSUFFi3uGGQ/QxzEb3UX7XT5uG7XaxAJN71TILPocdiOpRI1
neQuG+/RR6zYIMY/0Nro0Hbk6JSop+tCp2zDe4tdCYQuOTRaDd1QKnSYyeNplV0PdQI7Cm2FLQCT
GajH/e28x0W1RxJPmSttSiILQOgMKTz+jFMWOJnCiwe3ehjLGgEljktxW9y/aKBQ+XN0MIP5PrnV
+1FEakCusvvL00aklqJ0ALryPVUzGBi8ZXLRlMlZcNZe8AZvtSeCCLzjSFd4QvN08h2R6LW8Vkne
6IO7ek1SwG7/MGXXewgFP3dQMJGUpDx7sJc0mKhC2IHKLV5YYUk+W0UyQnZhnVz9cCb5QiTFktF0
Eus/9/efwXpVHRPxxHPvxPOUcAVgY2Ai0lgikd+uLO20VEGf31GoCYQqD90en2la3SNbvJqTGYSC
UZ1QeJEq/nCZGyd9mBfQc6TbqLR2zoU4xbQXx8mDTBajU4tUCaD3QkVSmopYNN5RuYwYrFmDwSMR
sDpIv6vhQqzTvq5uLKoAm6ovAlF4jf9JQB0rniQahXmTe8ElSac69EledYXmCCfk1fXCT/HDFiSk
doZb749vy5rbe/BLD5auh5q5VlEvQZoeykmsxbQPRFbEFZq63J5L1Y6kpSSy3RXb5mV6El/boKo2
LGx6dusmU3UKa32qUsHxvULc/2lWzFlIC2J2mOE6BxLJRSMLYQpTAg0sZHmwisowALADzzl1NXd+
b19p2MZg5GgnNcivhi24gsXG6TnXlEJbR/9VYu5kwLyllNo/5XCuMyiwA6+vB3s7tmeH//zyOupu
uCNkBiE4hXmtTlARkCj02WUKP8lfV8SZ0pZsWANSgoU/pnDoIYbrQ+YC2rlbYk9NdkIDOuxd0MVB
claoHZStjWZuTu+Q9b5JprddPtchu62EXCcDRHTkdt+ndcDfxwAYPnHkTBd9Rb3M4PApTqIKVt/G
wPY5pBYScU4g5Bp1kZzru5D14WkoHQ3YjT2kDq8Rw3+EzloRG/kmrjmOX8Y+e4Ua1q5JN9msbHkr
KRxWmguWJQ6/jBuEDVw+isgnUq/SO7T5PPnr+4cXD4XSBs54hBkn703FfIiiLsTNdngxX1+snGrY
WYbAdGiXTARprpEmft5fMDY/1DK7yXdbayJjIJSv0m8DvFl0Kk7WeehL45Cq7oMVK/XHJMd3F2Q7
Vpv6F0YKN0fbzsuoCrkw1L4GM6eO0gjD6NW8SPeWx4jGgGYuC1sW45CBYYEABlSJcpp/SWfFvSl3
KPjTWp3BDYizRpfPu2PSny36OTuPHarrNZr0GM/e64MOH0pTRyluoO/MGxfigOrpoFtHD32bG05k
XNwS2qbSLMai8ltb8j881oyVcQYmy9cssxY2QI0XW6NbZ3bhai7z1SEWUSaGwP2Eo9vYtOi5FgHC
Gim6QdHBd5o3gAvGGYyixE6vBTHs4QCLR46LSZaz+YdU0qgxdn6bSCXTfW40xAq1tqn6mTP4A22N
sd3k6cxzuPMMogVhnD7LynEjmyCfz6ExcjkYxymcu551awjXvbfSX+DESZtQf6kNfAaETIsR0jUv
3ow3y4p5c2FKTHDlpTmXYSFz0CtgYwDKa5Wq5UDnWmAz7tojkqduGaxGCje2KBFGrYFcxSJm8Ryf
0y5RCF4OEdhtaw2Mldtj4tALrgRR3VhhmBNVoFkSN+fayw3ucauYZ0t3p+7KmOi2+FVpbXYyvuWe
siDYn2nbXxzYipTmbnj+PSfLvsVXj/pF29acuSGqhwIWnexQmLSAk++oZN/WSgnNIyU5tnlC1JI5
7b9In0ihHL7cTSyNWLVe4SUyiGOoq90Dohs29V9Eo2EVmHiRxDu3pfP/OJkB6cVk0f22MSwXj/Qf
PKhu1Ud+PC4cFyxh6IO41de0iSV8CX6J4AVCdECm0FgQ723pJTbJIR8IuNmxAlJ/loPVxeK7krsr
4WWvVeCvxPfju2D5B/tZmsEQ1ICG64XBizv+lCFoTNX41HBYGHAluF/WAXOUtMT6aWH6KKTwHo15
4poVFqNHk8aqjL1Lf+ezJgKnzowz1dMKba92nq4AcvjqPfZjrZ8gDboKs/AY9QuJMYgKLQaLXa6W
EJpS2W7G5bEXB7BAWqKOpKb5O8jFSAQ8mzx11/L9m8Rk8Bh/2seE+2q8HiW4tX/7Aal/EBRczYjb
u5zi+g2uQR5zDTeK9XQB6FfedX9XdRi+LYyFNb6LYktw3NCnqvoTlLqkoNeWm4ApB5MH3A6x2nTx
JS9qar8CBnGqR4O6bjwRLzQcD+D39J450uEFKH/H7vsYoe147nP3YQjLyEbe1dP4lITRhATKzcRf
0EYf6yg+TYwcmM1Ko23ypZVY1XlV5ry7IqW8DJCIFprnScHrZadaaC36wqQuiKppMVwCEZL3D9q1
0ym3CIqSs+KwAFtmoFIER2Vx4Xg5V2+U67iSAc6VSkxOfcqx/N2RKEB6WMR0KXA9uq4j1P/cxa5+
3N7tMLdPZL476VtCha83i7RrJSmc7nTWnOLm1+YuJlXK/WzMUEW9ufb1WISPtxUqC0E9rB0gz6ga
g/NDMi6HzRoWCF2kcd/zOCh5oJCjzl/Rgp9puI0+EHS2MdoRw7/1NkOAYMEp2HMmoHhUbAY5516e
rABmqVEVby6rIhAMlDKns7htE9qtI+vIVdGVX3cblFQe61jQYX7szPJa+nimoQhkoaA7TCLUc882
LLL+ef1IZnxwOiHWhVT9I6/ecxWtsJqCAEyyb2VMrLhusCgIPTqjtxo5gtTRHgmeN2uodsIOgzvh
8K3EtAVkwMGDJctkSAAWxeXz2XGaTbaSaHGF5uwow7TukAdenJeDHxA8SAB2gqm24XwRYplpk4CN
hhNnyx8QzGmllxzwVOyPeGY3QhiiL+LFneFEX/Yp2IStsxFGvgnTbmFit0H+MjeF/N1zQGp0Pfd9
KEiF9vlp34NePUU0OSa9u9Ib9s0INK5pGBXk6UulJGbD0fMoBxS56012GbzEaA0CObUkHu2UMZJj
yYQJNRhygo1bU/snZhlDx2fIinUh321gQpVSLtj39JZ3/hHwy7a86tU4nrZPGspEAAouAQxjJFDf
OfDkEl5EPhS2+JgfBBRyVUIF4RnIaYnZU7YSex4zGKHK0lY1b9urnOezOS95VW2aJiHvgPecWTH7
/vZgb8FAc3QcS3Wql5vxHqZDBwOnhV068oakuYgUyCKdzeqTz2YXVTazQNRGYXAdLylZT7svX62P
x1lrey41FV1LrpXdtZIz81hOKvCCexkNo+N6Qy9SWvHTZyUPfN6Umox9fd0/rUE81xC9zwAzgsbr
S/BoZguyHhyWQGEWxGrH0ql29wwTEzi5a0q0Tkn4p+e9zJT2k3WRrIMxNZzigUDl1Jv4xwNZHG8K
6+wETYdB6pqrgQ7vgYtPjBD3bkmflGHqBHdwVz4og2VJs2S/debAmL1/9+QvJ34xqJudk5o+XcKd
5ZTToJKM1fKQzZmJXcghE/CYt1r8XmvFNDARRc/3vtAN4ylXELXwyjbOAmOfQgHsTQlI0b9Hbgyd
zP79WG7NpUnccOKvs/lLaSnKKHxo3okCohaKtpC1k9zhaKtQwLi47aSEHdRU5xZrbrPwbVfmtiiM
t118umCi1BhxumFci4RtmXwnA9Wp0GENXgidvOMDzCzWa06TnZ7up0dfcBEXCL2VCogtmJxJMKg6
5fj7NcJFnF77dVqBlwoHXgbokg6uVcq8feKgWX+S9dgJC4YQZQifpOo5GZl8O7I5IYUQvQ1Sj1zN
lsctkNtFnWCEw0S+S87ejqeOj1p10uSJtQ/lMEXGmhSaupplFI+CzmISay4euJG2u4h2gvpX/3R1
zqlf5zR3N+B7ZB8+COcj7D6OSov/GE8fGem+yexFB77P35814kJi4/S5Vbjuj7xnY0BdrSNUgd1I
N4/lh/0UsOwChtfpyyDy56da5TTFvuPAeytGs/ONImlFLFHcsvgSAWSy/aQFA4fIaJ2qedPro0UC
XSPRNAN+1ToMI5tSAfg+iy4OBonbRDMIWT29C/ZuZcueRS42FJZIcgTx0yo29H/xwRjEk1b/m3re
ncmjq9tiqOUygSzhqvI1F1OLalX168deWS5P7vk4SQlF88NDzTOP/qDIr3i9ZAFAvfLehCFMgpfA
glX5NEtsswAEBDA+qOhTNLFSmFwYeIJjtviisd0OkB8yJeg75FgeFz6UKoog0xM1mcyDMwRERZJl
s472v7lAJvIiMchN1f/eIMJaY5YnO8ul++2YBBLMA/BZk6f+FJVVDXsurLnIJVbov2A/2EGIAD6H
kfIyOFwt1ja/qq9KlTodyxpWDeWDLUvh1BnTi+G3ZbE/WRzBfmg0fQVqD2WV2zeIc+XlCs7TW8ke
i5onAuzQxsBaWSE/lQ0ePBRID0VBJuPAZDelqmGh/2UlN7BaZDRo01zZG02d+tgPgH6HTz6hC6so
4CUlhurraOa9F76B1v4puCnoXWFi+I2jlwHuzgfihGpx0wyDCJJLy8AWMxl5I0p+7Lp8MS1NLx96
QH+nzqqfeue/FL6S/IqHrjbMH9qlVLOVxX+Cn3vfYz/QWtmRnq/O4bh3YgbUT0NijFSlqxs8mV1t
7k29xGIxpuKha9TYoQVuw0/lbPMxd7PqTOpY/v33vmP9NEaTuR/YXjZ6CXWDnVqFdhcv4uyWghbt
Bc2c6cUUiPSgYaBasPrvLZNIava5VoGxdsUasDwXYS3H91JkCRYMXqz+EgH7mkGjX2dZfPzIe3dH
5DpxeYXuR1aoFEiErBYDrMYhJ489ch4B1JWbllYqsSj/w9cv6KAjoVxES7NtsANVGoYKpWOAml0/
5kNceAcORnyGCKsM4E7VeYyC0iGB0+S780x65ULmH7oRZDWJdVC40nTpYGtP/klqdNVJrqNZt0Zr
U0Y9ZmjR45ghTRCj6cZFxPCYYtM9ebxV8oyx6UuuB+IdI4xXVlAe7s7Iydsxin2Pl0uBrkBRPH4O
7RsiPFs7nMYjBvQ4Z97wE6A+AxRhPWC9ADM1669UXREded1HxZpoagecZc5zk17DJaFwnMjDqrzf
h8iTvbsJ3W+WCBS5PGJE8skJQQNu2bkqSHCK3ThB3yXMU3cQfEkJDb5awNHszmHBvtmaREWh7IQ2
Gh290W2sbkhep04LjWe5530M5g1rxSc+pLT9GNoz8gFGF+Fh1ZDjqR30iYmgRls0vVgukaZOJHqf
Ih7cf/zILRdVvhb2bbwa9TLJ7oCT3EZXaj6cwS2uDHvXW9enXd5g/MgrfsIsLPlxrTRtwVa4V0LT
i+IkZhNma6/U/t4AT1m7YmT9Mq65mpJfDgPG5g026qRUQBFFRVwFxajkjNHs38WEU/EcxIPM1eTS
L/fxsO/iZfSAWmxzi3Qzx4blk/G8Hebiu4blvaotzaISv+jgn6ijU0aise8AsEHHKwQSxUWAXzSp
iVgQa0bfOoxG9mHykYFpgPCmej692kRDEIMVixUyZHuGIYoj1RHbotPGHnCOYID09tHkXaB1gy9L
6cvffCJYMCnEi8SV5FkEgR9do3CKMaF3GgUYzNkg12QOnr6gt0J5ctz+JHOl7OW/9I899YZeFSx+
PbUcdndL1bQ2u68NBZbuXWhYp7/Ffbu88ec579c9b6+cXLeBHMtMr7GI8IHfNMuW68z0sQL8yAAu
2xMKSv5vF2TvxB+9r+eEIw8HE8zJtiQGQLc8JunPyt6+AN6j19Ujh4I0TwfAdp9z51kVo+olzDaY
cQ5ro4fCU+jWPmtRM7fwLFsZWsu6s2029Zfrde8mY6Up6jZfxb65vBOjT0jM07Eu6Vzqo70Zz5cr
Z/h7uXdNlGEazpCyWt84K/vfL+7zFC4UYGygqwFtjOXZna8nifN/148s8RsIC+Zizjcu8KSOQNak
3QXUxzUbQ/W7/n2D79sDl4ktCq2VMJgdPX8jiRwdTRd1aljbN632xLJkxeRaaER89EM68Vrgw8a2
izkEVzHEn3PH8lST28hbJ/qTakftm+Sa4O/OBQeRT11K8G0spz16aa5EOdAEQk+1YHOS1CAW1lAL
16Ac5lgf4TtKW+FNp1xp8YQwAp0R66qNTxhlyYO3JPZi5JqsAE4QHOxTIN/2iiNusp32wgULUuG2
G9HpouGZD9zgVsq7SEtABsDStmh2NYNeKXYxeQfmZ1htQlp8tl6XSDbP+nawS/cSx/9+e46fCjeY
XW5Zn5UvT1UqVsaJZq/gcaMkVrlovWlhiPCUxeLOwjdWpirOSIF8c3I49yZZ19KGkatmHkZTwSAS
4P5nCsMcZEkK08HYtcndWoBJ0USB6EQAGWAb/0s4Rm26t4CjkOthicURAbbtiM4/e2hw6HkrwxBJ
whM4Sz11MWy2TmT5tzz/3UjM+sbG/BqbRbm3ZdKjtiC3kLlpv3oLBmYgT5+QvpDuDQBo7VRzMBpm
3KaYb3izWysauna9rlV6XA/bXPKbpxs0MT7TifgVcHQBojGCixCKeXmuuWvdMX96CevErDj/mk51
LezVOcLR7DbDa1XxmbbD5vrxvFcWJtuNUPQQgVk7MiWBq2EpmPVl8X803Jfthha5NeUOx+mcYuZS
TCeq0w2SNTwloxZusCyyDktXWXK+vld7PSxJ4/4+wPx81ndShK+jPwt2AKeKEPdM6ktGGqCA0oaN
2XaVdCI73OjKiBxMX+QA6WJWYEeOP4e4p5+I7BLnX8WV3v8ptwhUf04Ll53wRyk9Hah1axky/XW4
Sc1oH5qc81ynT7kZ0awQohVA5KXpesjICCzfa2D123JxfPtDKj5wdLuc4Ez1Wf368zDirZlSFSm4
vQzpy2hlF0l+2hKDFhPCL0kcX3TPZ0gLmIGLBDMHDlmqlbv2fn9mp3rzXiqAgBxNh2T7gXhAyfZq
OTKS+xY+NRY85U99wlVrXl/jF2mc9/GFkO7a7BiL99/F+oWWt7sxhedbGiWtRdgu9rLisXODOe6M
UbbGJRDXxhe/KVrh6YL07MB0PZYswoMxJrR0dmvl9UAxmW4xPNyNOF2KzlNY6aih+W93wqDi7hAm
PLkoaRN+11uKNlAqfFZ6SG16HJiUmwv/6GLHv7b+QMzNKlchpPqlJ3wrRnLEswVI+2ezELZ9ddDq
5BO96OlljdTRdhMa99Hbd5t6Xd8/YiFsctgcZwqjFJgQ3UnvOx3Px3Upnsk12TiSrXdsFBWKOpYx
s48ZpdcG3SDlRTnZNR8w/8CFuA6inOcVUQa39vH2A0Hat58JZuTD5F0wxt5ZOGGyEVrkxwmXn7vm
IGgtb5523DEFGl8d7KFLlUHdl8eLJGah5WTvRSbbqcB9GvpbMeAAIgwcgHwwtGDxysR+iDcfhVPu
Bxx3yaVouFXQw319AW2SorR56L6ZbB1h3CP1cOvkcASpeIfqb5KIUCd+GR7RUVk7gzCihskXkHEi
lZr4sFzRnCLzNJiYgMzaF7e8sLIm0lUkyTTyNRNzmV9HFh1u+6MIdJDNW6WMETLrP2xIDgxMNjpN
CHVYGhjJhVzpWfY/Lt2r/VoKfyzgmTJPb/PwvO7/OqKPBf5EuOnzfpAoqWvs3tADSpvtu6DE7MXz
8EcyDDTUs+CXLJfEsr17BiwFus3GgGlZAT5/6RUbHX55jG24VnroThGAd36C1Pmy52Q/2tUXuSPq
PRD9yaWLueSiTnPoR+HKbBhlvKyROgp5t37sKBjoFQnjpoWj8cItMqpavysarPT7PG9+xnbA5i7w
K1q9IfTwU5B0gzY6bpyFhIF7YixhKwnfzw2AaKJapRR9ZU0ORr3LuRAfiNklj+u0Yzp1SvxyW8E9
nT8WXQnQvJpRQlHNXtRyiKzahM7EOgTGfOthyyc4EdC5fJTyiLcwEPZh/VAG6ZoT/zUgCUqd5+VZ
sovhczVvFpY63EPmgDDzsG91LkCD1psUpLrx5IfxDruWSHf49UHR00dvDSxpcz58iIrEW13oe162
mnPZBZzvW646jKqlG3gNHJDlK5wvbamT2zYtsCunzgpXfCfNNFh5bhlg3VIFAPRGWCggDK4r319P
fh8clPnpSVaCtXtcydx8ics9iZlPYLu9bMCXgDL4uwX+ks4OOqeE5gCLsxpphjNwoRf02zJj0PAH
oU+9Q6aQvT+/V0H8IoZ9wwBm6fu1LTj+giuLpbo/CTL+s8xo34xmVd+hASNTKtyu9LbPihEhJUmk
CG3i39FZi2t9bEYQhsUYFS2pTobXz2Tv7QvLDTu/IyK2GTsxc5l9CXgiDdjjGHyqBAkut47IeRfm
Fm+4ekvdlGShbZyXvwzcfwiFiFPn4TaKCHna/SE+Sfv3uQEGMkxjFRzoJsuGVxVNYPQIjUDHEFkW
1m6flIcT212w44KePDgRnEAdqTWCmMout3GwLEi0irOdAiY1IRST5q45IP0DcQGFnn4Ce6FZlvzI
loJTgFPLwT3pF8ee53wpFIO4ktd3Qoiosuc4ytMuxKGf8FUifam0+xraGpKMZILdWuncIbqNn6O2
j7a+RxuqObaI3/S+1re4CdSsvZnCpm2z0I+p78ZsskvYbGkhGQmlLVBeQOPxwkRB2+qR+0sH7hW8
Fgn5GEEWvSqA9CTb21FSMOuaZYsFchJgucAISgEHRx3BjQnrwl5EIs3y+Ut6L4Ys5/NziipojNvq
7odLotHxDSAwJxdupmcWNkbB75H5XyrA0xGw6kF5vAEr82ncJ2M8fOwh4vnLYxANNsRg5+s8D2RH
dkmrDdOR4vJXzNEpVd9yYZiHvdIrAfMvgyV421dioBcyZd1/KReQlWSlIJmU3bnQABUMdu5I2gxI
tmrt16UcBRBDsquCMzY4ya/v1iyuMQXLxV5dXjghQgmCAoKteTgv18msw5FlC+UdnCkWwHsqNTlc
HcS5FkMR+OmhWsvYD84a8dFO8zqWTG7JO8TgGMmf6zcnV0DZUVxGxE8avcIqfz0fcOxoeZF1ui9r
MvWr41gtKb9A3/sybfEVg9P/7Pq6FWwDIcL7BMblBc9OrzW2VpcgryatoJKROuLd6zZwkLM63lUx
rV/G7boTM39tuHQs93RCINKkcZYdtYRF2gm9j5kKb2QDIh6Zikqkk6Zytg+hM4UOOiVFysIckkm2
3RTyD+7/RcYVZzl0qobuWhutagGHjUbdXbWFA3iYuvLrU1LG3CHzGhkyrsdhmO4b1NIeahbXixFT
fAEHuePnJeGEC5myXqNmmcQbOQ5kU0WRlDTZ1K20PGgo94/dePQrhM4Cbnd8SifeoJ3iZWCeQyGO
yhI3Wdc4NSs9+xdvC6qPZGILumFf7WRFxqiiaRoAAC1Lu2dLFkk7FzW1Nq5J3zvXPPJmr625Kf+p
Ksf/k006tioepB0So9BQq64ppZSleYnG+0IS+Omq7TpA/Bs9T3Q7Pv4k++ZiaT3/HvVVpT9qmmjh
JRf05LVefcpeYrV+ylXKOcGo5+rawKuQ5kv10gkskk6JYBuqz7A6BKz5fvnfPDIM6ZLPY3KJPGuP
qPebKnEwQqqUtj2zOXTqHs8nIKH6uQNwj8zAl4HRnkIjyo9/dH3pWV30LoHdyAPYW0duIPiJ/LSR
l62aW8xrb34Mh2GtrO1TfdN6ocildA3BMQg7iLPNoQ0JYGWi65FzVgeEPcP5bI5a398kh0SzA3Ne
QjMPH4TzXmTfE2t0x6CJtqmz3Wm1TsBL2MOUq9byHxel/COjYmWdppQz7/kYr/ICHnRU3ZVbUahs
R7fk2N4w9fJDokgPwkCPcntaMPfAIYL3jB+8IXAiaaUCQhnRc74f/VX9U2UL3fIBmbUnykd9reuW
8J/3oBIjPSRixNJs5728D/Hw8fAjWfM323ftMPKwDZLPhG1tE8IXJhkLnYCDPvzjpSZcT5+VWUhc
YT3LGujIXIEd0emhFgr/IMs9UFerAcC1Z9LOotzKRhojR8ZOZRNw5hitCFFVWp8JmZyekjRvOCR3
Jtj+qbjiw8Qn0305p3SYqSbWUnP1OdmZ0z07BzkCkiLsxo97gvEyJVAm63I90OSqJSCLIMH7yLkH
BkA5HvTD0Qd1bJ9GrPfKodGqsTz0VorxOo0+w97juzitryPuFarjXRlmWtjnNQQEKSx2GRayH3/Y
1jvgSoyl0qqp+HmV3gpXq7WN7+GWotKB0DpcSe5TXLxvMjdDg9zyFBgvfWwTfG1mQGZnQtXyv6CX
/Pkr3ruvpVQkDMO+Luf3E5QbjrWo7sXbd2yxHajSsrDasBu8Uk8Eogkd9Ee4fP/d9QAY6RK7aIm7
J5XsE1r3Xb8j2RZVJbl2H/9Yxy+ibqP778EdpIsVKQ8XsWsiDAM6aboOtSI8VUp1yGsB9CmAUTWC
N6ERqSCNAwbgdwikvrqIFr2QcItr/5AgKHtgbSJLH8y8pR/K5kAFTaXypONTFoj6FlxjFuMHZyyr
TDnqOjYX9YWqA9xautxbTEZ3ZweC2Qhv82KZRzCXIJi1stdm8r4KJZ+Ok20496ogIRVoe3HoLbms
lLJIuFCUx0H38lvmUwwnt8e0oaIeNLfWZKVp6pCidXDYVpTT5BvC5Vn9dPM69Y7HioHoXETY2BRq
Ad6aVrQTzBfA7tOO/rnxp3Ig0toLoQef+GFCPICwWd8a5gShHDK+sJ1i52ZPyR/7exE5e1ZU+ogi
9OivjH2ajJ0dVtWI8ee2UPvXyCsnXYZVb7SMngoeuShjMs054jD9yREAPv0F+BATabVFcWt45BSB
0fQ5LWTu07lgpdeXk4v1tIjdbffZ+oWdQbLXsTPfPVywB0PPx5Jt3jhDTaT4JCUCASMLER1G/V5G
8S0n1vME+VhiPTmJfiyOoNk5us9ZcnsEcLkz/hWzClmO1NFx1gyxvrkkF5eWnw0gSbXqWL/Gh/Cp
NMHntH/4Y8li4MCRFRFW9ihUdBkc1VwzTDvWPZY8neVkFOiMu/D/IZH0Sq1sS7MOxzNDj8uOKmin
3e3UF4Oq6luGmiW9TOvQXxRKSiSj8I5SekoDkr0PrMhvkvQueP+M9Vh4mANBidG9yWDzvwJGKwg6
6VboZTx66Gj0hVNbmt01SLYx611rOGswHr6dGYrt4AiwevEya9XK44aHQpUfJAW76GNIYAvE96uZ
ogEAsPpKL48ZgrRIOIiFOMAj/uMl5qsurwuXHC2ZMJh6FfU+H6Maz80ZEoGHTG7WBSdQi6iSsTaH
o7dqCVw81Wa32eYVn3t9OHU8XGA0WoWm2kvLk9VGheGygayllxPHc1xApJPJ2j3qZd7ooGxv3tJX
7lYwcEnxrj0EYFVCu6QeDWaCHdGDfcxcbgYcztwY6dKmN5+P3zG/4tb6HDQoIOoZevVOF9o6GPHW
S6Il3I9FfixNUhZF+mzPz7+eFniJWvCznszFIs8eAZ1vvoQF0lVD8JLEoT5EGJCigVLhiyEe2HJJ
wBwofi6Ketb2GAkgd1Mc7mDypMkvO9dd1zgJfaFOX0n8Sk3E2reqWWO0hcP4rhaUvEnfESSqTW6Y
W6qVuTWTPVYmn0bc+8ueKyan1zomCmu3VDhcJrBrPV1FWwmhJJIMlsNXy2aPOakgibFD6bwWUnaO
7xnc0AyHp1bOs/BxRzuoiR0nic1c+TTPpBcf/Nta2YBbHXUd1AWU9WgyQLfXe6gKN2lWsD0O0zcC
TgjV2xqvQdMiNStr8t84i4YWbpBlNa9j1Zp60iaEOyouB9ZQnfbci3ULrruDcvXV434wRsg/7x/4
4Cb973WlHZ1J/H+izqXqujjW+nBmCR76i1Lf17Nd5RmiqyCvW/IUTpiGEdziQCynt07TQrzQTQ00
CmJReZN8zwvlT9kYdmTk4/gkoRu57vl6DwNVvxEOVlQ4l3KeTTobsDQDzPA/KvPBzPsKNrJX5tdL
fFkDez8/jO1nKxMA+P9RaZKXFi/Uy880mZzTBmPKRWFJNfdSVmTpfLeOViVa16hIHjF/8yFcInDp
OiNMNI3eHo4SvHhsI773aXf8L1UtSagI0Wtkl5LwRr/N53cK/sYoTp5NqgVU7xwWx5r2Tl1oph3T
uuPLWa86/7c/Hfsg3E9K57srAou0n+V74lUp6g1pHJzGfNX1UHX/NlGT27ghZj6uXnpmf2ufgfeb
hvLI+ZtJc4kbzIFt/k4ziguYrVZ+qPC+pxKxIwoHspaOMCVp6WfJDJgR1TaXpBOX0F3GTBER4coA
9EU1R2zaaZLqy3WnGpsFgGLKQCZ0i6m6HRiMNDJKTMRqFYtVFBm9FMKZQ1dKt7EoiTtgHG3dC2W4
8z0kHZLpWIcm5QP6zAEtPb5CcwxBdWmAdJJu1Ujd+ae0NgDxAHc0bB0NIXxbaVIpgCWqEp/icfKM
QSjJgI3l4LZiD4CH4RVWihZaC1O4Hh/bf8nZRL4cs+eltmpmtzzHZ/iUf5bUteA2jhcWO488mkyF
ZJdXuxZF65iBJAxb7+uck5pkRhzczkNlqOtLcU7CeMGgSdUn+YgURdHodDj4dKzAnRfTtlCW0Q1M
KEiwEalbz8sVRxyZ5iurWXpEyGEnDkzE2MGNep01RRZAWN65RB/Qu7dkeRhedVTZub5DFstEEGDX
a4IWsAHfyjKEerRE7c127QMm8XEWwQGvSQ02FzNrgFURbltMYwDQGbHCh9BuUtHuqTVq6vdp9CpP
I1nR22DaxJ6BlEaauQ0Fi31CYfz834CuGYcHSt2TBj2zHtAzDyGJgr6sDXdRiKvS4P7tRz/eVyfZ
ygL/az25WcK5aDFsnKqxVoCVcd1X33zsOCM701bi5/x+OaK8xZPOFAE28hfHIPzEqt77Qhd6Oqhh
sBLLOIJM7JKDHbOJysuEUR2dUuhzaahqS1ibbhtLl/VtKTlI+YFLqCKDSf+W611/WhmR5eCmlVzU
U3UZ9GbgcSylYL9QQ9kRj27nQ2DdLBz9r/oa6bxG5zQcPi+FbBq8UGy/67eONIW7W1+ATADmj08x
ajs/RP2naKGThRg03OHFqV2JC5TG+mPO6KbyLT/wfS0a0DeWDLk3Itxa2JZFWfuEr+o4reI1IETN
T7aNcTaJ/QLjzweO/FvCbiUkE9yp1BIILJGQPJ9Os3x3CFJfGQl7lriRCzUBUHImG/RMwWD+Zctq
0xJHhacQ9VGigHr9bFC/67BeUF/pEkL4xoe/TDCSHdADkg18w6KmdqFkAbQBJ0hCX4ectky26mhv
Z0zS269fLLJEQGOs81zgqhA1V8JLHzTr8rWsauppgvd8HprzYTEIOF/qa7ntxHfKs4VUL65H9e40
ID2AuL5IUP08ZKCcl5DDryuq9hXsQbBN7OCUc41DHRvQgzp/fidlFHdqh01KAdmeAoyXpEeWS4p0
9GRSXsIVdokuYIfRKg2N4kiGvUYinnlAVlIPOMuJrB85O3XSpJcrTfddc+vHFSVNxInxLhmSh8QD
NMhYcEARw/046ZWsB24gz8i9W2nREcrGArqCh2wo/PAp1xDiGV39m4/AgM0ZMAGtNOB/PRelsGo9
+jN29V5a5xJBfbhC/TSRRMO1PQIkb7y+u5Ffn84eGx68ZsKISuF8rvLngBDxkMwxcLJctkTGmbxr
6za2Ak6xDfcakwF3DuQiW3rxOA0wSlbnwoCfh0NNa+sHsrE1E+qgnvc+zf+T0GKe2835apZ0gYxK
4vErLH6aX85VJ4Q53B+t1UXOgvI2BI6wKnB9avFuINViB86Icn7MCkiAOHcZ4CMMTRekQgcYo2WU
esQHou2mzyG/Cd/9SOAJ46bZjVNtp+lImza89+OpCilALyzHCfwIr6j0q+9v3FwZ1XRpNaSEuJ08
ECdCWquzprybQAr3CNHYIFFLcvNIb95plhGu2zOZcfnHQ6L4VRpp4wTsgHa+BqJy+iWChAfrl30E
3EvlrMUFvW8hR44wElgbY+4NzEc9SPl6BtqL7c4OhEPl04apg6WBLAH7fZfocC9KTAW1dmnQPDvA
iFL+nGG4ftPRGmSEu8mYYBjVz6CECh2KAUv5qsBUGZRZXlb+PpNXuLcqlSo21Y7mccJUz/Kl4xGG
2igasV9BeWYRu1tgT8wjRt5y17+U4FId3ZHUnxPE5Ovykz7/EkkOt41JfuG8ZlkFQyJbyf2dmdcH
ifB25PPasS1EyPYHi8HzCJgT2K1jUcIXyGuiukiC3wmzkWoUuXDhFN3tqi97UVuXqekvGXOSYCAD
xx0Xf2juLWYd2QV3d+kNBn8SyB9/dpEGXH2HN4GaEflILFS5jF7ROv5EDdu9K7gZjjOLBk4YQv57
HPFQ7vpvotzj1+E9igT9j/oKcceKTPaVTSGMdJ+yxD2QEwMX09TA7S12BLe1PGpQUEbespyfS6g/
CDsWY1lFPrPf2dfY90pqksmCrZKeiaD+/eQIN5mehK7+uxsERwS8o97XhExAD5CZDE5FwnMz5a4L
MizQ3+GjlJRecTatMSOor867XyWztTeazNuyRo8LWsplcWTK03jHTMO1k3s7ntzZN58a+UG+Mv6u
6nnyAud+huFAujqPfVcZB8I3OuNyhj4QZKII0AswD7rNuH7hz7SnWPxwaCMGx2YsDL3crPU3mciv
E716k4ddbnzj66NEgTRyclGnWjFYlFI1/mGv8JnSojdJqT4FjUTjJtR2dVElLPvcPSO7nRV8XxGX
8O06hl1ZiDR8k3J9wuZUlIZhvjpG1YwI09eJp6WDTNZ+VA4XEHozwsCu7Hkqeg9yvwL+k19DbsqS
D2uEZ5m1n5EKvqZPrKwDlVFejvV9oEx8MrJBLtXcQcjqCSAra+sXr3o/7ftEkCHQh49P78SHENLr
icyfLG3lRj+/5eZ0Gd2AoTwKqot0UaTOxwqrhPNyKeAltKEh2OToEb+1fqQnAs+q1tiUdjMUZK75
qK+8G/uzbdW8m0AfDGRNolcxPgZrrd1r+dZsPGGSdrlIwSglBqqEJSDWycaxaUzGGwJxW19ycTpT
6VrOgl+AnwEwZsJtVReK6OtvXJtGMPs6+ZdknJ180en6sbGMD5HN3cDy5xr81NbR1BrAcO9Hm/MW
wlB4LIQBxZNeLo68QOBM0SNRyys2xdDkVrX66KJCFBNKv5RB5sM3m/CRUWsFIG+nGSqoe05HRzzy
Cjafojfng+pFBMDCnDOgdoAQBJVlD5vZ3aDNustkWXUf4gUyLbxScUf0mSnXbsSx/9QwtEN7BvwB
FSy0SiCi0Sttvn9A2etgJGWOqyhacTbo8npJ+JV8lUKkX0KlHLmdLfRuO5W5IZcLwSzYquEZcazb
dLzYqAGxfMyZZFr3j64KsrLPwBOyHyCqR6WnE2mDznPQE5kIvaLMDeqgGWhscIHjVTeOI8rvatHt
6RfkyFRs/tu+ajpZrrOEqQ9TD2pnU+zlbYsUoFK2t9glxpkWNifKghVmhsDPgV28z+oOCAucincR
RazBT/X4yyLo++mDhU/s0soSIz3H631F5uUCD5y9kTRyGND2+KpvY3+0GCIPWkJoHM+IEugSrxss
ACN0pTBXBVxCy9KIMRmGgefDttEtMnPMppJQBN1r0PEsLVD1Wj3rfY8iPZlPHW9jegRhOckIZHEI
M2MHn4J6gNqNdiK/rOuMvWIZFb8WPpnzjoumZiydOv5VVPoGJHwuoRiMk6xi5aTLyP+NzhwzAFPW
HwPRNNyqGuKJ8xE0V3YHDrqYzUZwPFPT6+2ifGWxw5ANLK42yXdCs44iF2pX1QRzQ/+5c6URWXvr
/KkDu9XiBSWAGlTLh6xvx42LjmGV5vsgvHbMLgnwpZORxqSj5cSoQMMEFHY7gtAkfASpnWExdW2I
3S06H3QXX3fRP7B7u62dMjPe0KoIUDROMAxK96gGzFRTlhCxDNLQAvgT5CxEvia0EIcCPQOmcBqp
hPQobiwMXKPISjijFEZGyQta8/4xK5U5OD5HatxRStmvu5PknTVC3TOnczKI60ZIknPNikgXzOzB
i1gSbjIZlrAvgV7cQISlUhy5okm422t+QsrEZzWp8cmmg4+HuyMI3JMy0lZ+CdosL3/skhRPgPW1
AF3N4Tm/603f2teJhQ91GIvzAduqoL9K4XscYP8sCitAuVKATrvVUtSWGmxaZaXx6fai/nLYerT8
fC8G5NTds76+0qfWcjO0kmr6ukgG/wgMdjoSPw8KOpZiUnpXRzZckDHTt4cLrewFdbKa+2DoB2vp
t0yOSu+vYvDfewuS+5Yi7BqJoE295vaJhAzcBBTxv50G4SstBU//qU8zVp2FloagigzjcmDJ8zoH
yNLj8BEFxYRMeQ+IcLuExJq0dSnMDdcafyCJKDf8/v/u3htfXBSBWWnYDqGTGRMFB9V19Re91AcR
Q/quP1sI35NoDD+6n4WEsknXCFmU54yDfI9mDp3egalOVngRIktH6338e2uBDHWX4EDdXy78iHFT
fX/Atyg9nVdD0hXDhUok6EG6p487UeWs4BrjvrEdhLrChhKUU6JjpURGlPZGvHkCFUbcaKuFxM++
IGBCgcb/oJFgdOzfjc/1CD6ZZXzP0yylTwkA3eOm7KgZEOXHdeYbqaY4RVTc3AGmUkoEURrONNpx
+GxvbfW5QIgofkrFUSJBNj2dJyF8PmGNK7QofZqUFtzU4MDefUKURPWACz+kEV2VDUiq7Vx5s2Gn
PtNY1CHPI86rdPVTjii62RXowTFBqozLtjzApnoaEzOUfpay+MTYoG60ojxdQIwtySf5mb5YWaV3
fNT+zNICWukWAxZ/JRZQDnE75N2Q/q6Pi+IP4qe/tKYp5Ib0kFr5Yq5Yx2T/CDiypwA8oUv71BIo
IN5r4mEVlvFcPkyVp2KS8yV274ayGnwGvUu2bGwb3fNlypIfE2WuiHTqj/YmhwVhTlnZdZ7NN25Z
OG+4rNv9hUyuRhA1f+w2Vb9kKyc9rIkdQvY8C+TPTbdmpRMP9sY5lmQk7DOfmBMAbRxN5cVbCCrS
um8gLZMlCJB5CVjaBl3BaMrD9MCe4tR2T+Ur6HnOKmH9BUcoYpXuCbQ3LvixQ/dPZU/jtvxA15Fy
wvJpKJKETehA4xxN4rQYiQM9/EtYEjK58ysfC6zqXTjqf4wedHD7VDkfcXeUGIheB2p5WMn6eUHU
JaGOT/UdFeu9P6GKC62rGcABrB5Js+4dDichYZMTocSdvQ/hfPFhfEZ8s/HeJupVtkmp9K0RCPiG
Rub4RhQNEhgYSsS1Qdtw+G7i+gXctKUFcdLsY3Gv+67FJVAzZf1kfJ2L4jEu8vdLowrI99RBmXRp
xoYUDewuz2w7alJCjyF0jrPTiPL/jmAVgjIRJQ9OMDIS4CJ4b6cm0eGcw3Gii5bVLd4x8nVUd19d
U/ABtfqi9OM/FOzOF7M5EwH8UGd0rLjHMft1/rtxfPJC0eecoE41n5Z+G/7KHM7sxYAwneaeXe5t
pdEMbgx61wQTQ2J+LBKhZL1D6qFEm6jUrGN6D3tJgt2k/7b3xkJMy/X0AaSoedtkFudA0Oww/BhE
DlLunFKPxEZBzgJBHjOzfFPVMxYt3+PPW5p8oNx15YHWItec2HNdwBchekm6WArNYFHwZTsGG8y7
vDQhim+K/NHW5Qbr6Tw6fJc284QvP1MgGUj5Da7A5gL1cKbgHT5FTJ+rqONuoKcnHRa720Ab3XUk
X3e01mWtCPogTUI8FuPEIETIZeHLIwlCTIq6rWWVQdmd/o4rYFX0W//FWn3d2oCQc65fq1JO922M
my6++l4+CkTbntdnr8r/HeVImd9XP1oYfzJO0K2GacaChphVt5BJQpAR4DEJOzVFmR3plBrr9Wt+
DsTJkDDXyKalE3d4hiRC/nlgIxXRQqyT5ZFdbubwYC3Nzk2SV5QBzbdnHDKnfvfrHbful3AGZvuq
lK3b1yjkjxWBktzbFp6LyQPV41j4Q4Le8gSD1WMEB6o5eZJl3qFopBS7P9aMeYvv1KF0KvfRgGp6
YYvhCHBWrjQqIF9em6vdnrgtwQgdxUpOw56mI5rVQKs51QgSWK96cOFVa50tlrfRM1RL4cu3fvNf
9FSmUWRi8ntM6Duh/j6cLpCE7NOHp+/oTYJgGnnfNdyPd3ULGo7gdctX83rKwzV0GeyhliM0nB6x
ROpLzeQoGl4vNl31G273l8NaLnhTK2OTjc5bXwIBHm60BpGM6CF1qIiAmte0lLWK3ON3gXRvyU1a
K6v+WkKuISo7WK1q8ZeebcE5x3ghuqMZhOWpALIfOAnOilatoMIpMA3wGTbDqjQzdqw0NUzQ4QJt
qIWhiNbhy8aBeUK/kO5gZIuVP+uXPv8FMXp5zbOurxkR+OkqjB0a+2TCMpafRIHEV+sJqByuAAPI
AHc6544m+0yJyQxFxGJX1iyhBZCHh2IX/HRp+zpQS7VCkZNgIhZEZMu7QXOkRHwhmMdifpk1WZF8
oZpeY4ddw5L7HfBljMmmed4plNbGa4Eu7YfYsbCIQiOgQZAxUAGYhn7/LRIvKuncaLmZNN1SNFdk
b6+ip3FD4AWk9nKScomQ6afF4XWqKF0vsQOLU0N5uegpykBadjqcc24HPIqG2MUFce6/NzbFR5sh
0dr+EXe+sYPCLNkCnZlR6AWoJfWEvphOWF6+hMDa/oA7c1QWZb9wp+ah3PDtN4HQE06t6b8qW0dO
osHHaKJocZ68hJPUzO7HJ4fzSIYfR0puM3t1BvU0jadKtPYzw8+Rs20cb8YMarmtDW1FXlMjtfkm
z5hO01YtG3oBUXSWY9CC53IjK1MjHoHcyR3HkDdWebjij7hn5UG5llGy5X7mbbOwJi/b95UYc+Ou
A+fGN7NNQFoqppDMVSq5wri/0ZY3qMiu4OFq4jBMyb/PUml3CaRxdZflXD/3/LHfn7Rwm0ymJhlU
gFgG0l6dBFZJTELWXZZs3Tu8UiQh9zjBYsojfPpVsmztq9aBaGIdIzVu6S2yOrlWK8ofjyx7sKvX
N5Hi3gbydF9X8fdDXk6d3KmCGFKtSACbJM4dhT55cAiYWISug7m4WuB+3IzGE/6yARmO83XRrosb
C3pK7qYtPA6nK1jGzrkMqW2iIj4aRdNOiDCcQMfNnl4DP61mbBJxm6zlpvM/A50IIBNzLmgPDNFO
6Zw+nuQvVk3H3H6XpD461OT7SycgvKC5qHqOqU5CbeZuom7QfiwDIcfWCDhoW6+k2P3P6Ov/KmZq
BRuZOzSgq8MFGlaj/zKQXzU4iztYxKuxuta6zKgWTo3TUHFqLsq7+hmEW0kZEMUC2fHxteykEQ/i
mgOxhKatG7e7sxYixCiJjPbjA1Hy9fbnsJemUpnkN5TsS2Q6qgnep/t+WXzfCtMvks9YeBIhqV3Z
rlf2AXjUva6mXiATBnXApyumNGgz3nqPMgR5dLYBoYilyJqMSH7HuiXfXI6eLiZCF9Rw5LCrnmLY
432JTvxF2/UhEQvgUikESX5OGVNr4mZG2hB6OgsAZ6y8pMp3nzmZZ3Iw8YP5iinHXphw41NPvIps
ogzj4QQarYq8LAuMH7pc6Nf7hzEuLXjvNqAiSoczMnpBe4cTBzMTDG9MAMyyPGnqPIhZep0zYYjB
E9p8vvYYDyFST7Q9synfYseYNnmi7nlH/rTDnQwffp82RYfqojGOgzy+Nuw0/1QZidMXdS6sVuJl
9z5Ly+ihRBcS45Ar2Vd7bnLBm7q+jW4or/MSxsA3wvZ2x9m12JokYw9NYmcKWTDqk7wCLqosp8Ul
GtlWVfcfrVlJiKsTBGsF13+l6zrz3DNyBunxReVihTCHJXX3njBueUvdFGg5In+Mhmf33EX77NYv
t1oYZYOvO81hLpIcFENhP3HFyMuhail2D9kmZE5LG8hsBlXK5jjZTaRBdbSJ8UOx5Tp6eoAkwqDP
K7IucC5igGcJF7BjFtY6xPDSE9VpOXuzx8tsEO94/oSI5d4+nriCPgXz7RlmSAS7cJnKvkHc8tRa
KDvIMx5zRzj6KZ93z5rlzmSbJxRpvGuxpmX3xyx4cQyYuIBtozz3hXgYLUgkHccsbCNp7/njMkmH
HV2MVKyTzsg9glRzzQV6IYJNQApvcVbXdULqQY4/NZmmdfhzOcZY/bv/nsFMJRIwk7kF1VpVdEkj
tjK8Ozr7Eia6Ds5ql5Ep/wv+0iSFW2U6/rbIpNs7/OglYkgK7SDZiQMjAazYscgVAiWtyRvWHqjX
LDHPgNOAkqJ9DCw0q5cwFQxbRBu1ufU1+KAepPEl8tkSRN7ok6L8+8DiSw48J3ktrm+zqm7+23JR
7Kc18dmckNmxVW5JpGQVLF8W6pkJ5x44FPnyv7oazMYIKkpJ+piqhO6aQmXKH/GXm/aF1GlUnjMB
m4QasreSZGV3tmXUIjxFwp9oxtYCu4kOkfPybi2I5+Ev17FmcGhv+H/UapxSj53g4xwJhxSfnMS5
e7VaLV2rI8favXYagVSnHhVakSFU7H8Iv46fP5GzGLL/9Re7Kh66KDNXPYyEiprPv4fOpf0xB+Gq
05Y9VYJ3amhCtOVTXmgf4np22S+aoedi0O+v2jhJrIQtb7XRk9A5hiwP4Vw/MRj6hSDUZ6YCiBBo
zPA3XanAUE8LhmyBVYBQeL1ZHA8Cd4gQSN3jt8oUszCeX3/fTqFGSyWBVLb0ZkD8YJriNwbFImSJ
i1wwPSZN4/CVzogCWiOmWk6NfvdgRN7SBw8BEbBZ6TnpIwyM3yDh2C1JtYpgw8EPTGp2y7Sf27EN
9A0pXlwLesibnFN+PZ8qvQgm7/6YlJOsl3dydYvM0aDMoxNVrkGPWCgzOAqKw+DgG8iHhMNxsZSU
OPS2sG4LaxVTaoqYQzst7I0OgdBlCY9KRV8X/hvmoPWEz6bTqelAst3Zx29azoGlZlE1jMUHzqsz
oT3XAPd3pUzL10tXZKTbEYhwOnTVjei6qNfZIQjphXSYvLbUJ/G0O0fqec6/ETvoNApqvW9XG5fI
/4kiWmtM0Y6OuRPkjEF0QF2TGWMQc3tIFnLvOFwYyTHUzLUNT+N8BPqRde5t8xiPD2NrqtfetQ8X
dD4LDuKJFfDjfCqJlaVtgG29r+nHEY8UEhVpLacmU5SSzTmJB9AHO8OLCdbRYhYruK4SWLAylSG8
Cn92GCEQ13rf7HLSR8gZ+MDoyHXVRbfrxKYO8WbcXlhRbpENydskDQLFfRaSHVjgn7eOwbxPmszh
uXiLNwxBU1PzM3364TRsM5K+wGfzMOqyXAkK0AnqORbT3ET306VV6ojPlbutpRQh/l7HN4pBEL3U
aCnS5So0LgwwBQMRYGpuNNlnXxDcml5D7Hs8VtzE7/kaBceK+v7DNbHGR0xv03A1znm96TOcyO9W
jK3m3f9H8W6hjD92rf7kqnRoYD5v3K+X0wiTXoAsNr0zARzajnOGuYcXbmZmvL1ONd9ukLaGfVpL
tFmCsHgjfl2ony8p5CzryD2u08Q87MZIBN0jt8s/gxZVxg/j7YgzCh3cY/WRe9b97e6snb/Eevuc
5cfYmBCLs+wcIz/QJeWsyCguYIU/fAatz2Mk3jBLZ/sRgZVmZ6y/VaGt6KDKRFugFDm2Sc31+6mg
5JiQ6i7NHIzXP2cwuMbDaFQv5l94RzpDtkS50fKbKonh+tCLF6YBCnkwDkMIDlLLIvX66Nhvh+rZ
Rf9m0RbtvSasVFy/Cl3wX+bs6qeky5WMBMDdkhDZuM9A3OhAW2Lrj5Ol+pvSBOe3VGvvjkbGnv2q
iOXNfolsO1/lqf4E0XqlNbiProxpuEodG/VrfFyk5TrvTbWPvLpMgM3ciIedOQWW9kvrQE+wY/if
XCbWvITzipbNhadhzf4GvIX8MbpnFPzbrhzIHnLehFf5CCxc7CatAWGXKnVq9yH+G1pa/0bbKafj
Xr9g4gkvtmgu+8qL+U8yXadozpzJRHyJqxCe+gpsXu+mdePjIbsGFwWr2XF7TOzwQC9qglxuOIqy
47iDUWQw3B3GucFE6riZGukAt4l7vVmW6RXIx45qRsYMuOx/kWs89rQq2mRMgzVFJJf1o1PKrtRm
bph3OVpyMM8v9RyDUhA2hfHPA4SShZv1R7TMkPmJted4ILRXcgAIsDMjEwtkXgIeIvq/vaCppJPK
O04F7Q4JkryZlJXQtf5mdymoVuaRsTLMj0QYXPD2juqMDL6OAY8IALniYXTdbsDk03hKj0sc7usp
YuK0ZwVXWbyltgHiAqm0pU3Vt3V9zO7PMOFlPh05YBmccVDeB62SzbuEXT9UbhYa61jrtaGaBvVn
NXcZGGAh+CA1wsLpc0HvqoJ3s6/X5nY71gXFETIvGJKklKKJgN1PwGXCYhEefDUL3jOlNUDnGD3I
iEWTmiHj0Qlpi/QGaBHLpjwPCQ464XvofYV50efVM5++Y9We8qkTRf8KlP5a9ovOwwmGdBF5UNaw
A8asGdcq12pdpxnn4qh+JyuZ13WZaik8L1WkTPywF5TTJAr+Uu6SJTELv51InZvi7Gv+ZE079doL
BSOuHGHcEflj3sKXVG4syeIJzXR477NdQh26r92sEwTv8OSKYrxFXMguiDH+n1C/cE2V8kO7M7de
snr98IbofVsJZiauh5uT+NJiU8rneYU6JbymIDdwSmfOIBNdtTmpKwsGv848HnJuCx9sVQVwJmHu
D4a0GxHQgNZdFYMqP12VPzy7FRmMcMd1VOIvy/9rkXvOqc+GDoAYyZYfzY2G8P6T0ixGZ2CpM4/r
dwj+g33dZqhfLiTsSIWT1hR08pkdCEyti7Wva8zs05rPAyrExfd8dtGQ73are/kAlmZbGOqXPwvm
11A3VpqIzezT3nBHepYeRrSy46G0bPKCkw8j1/rkyaz5m/NmFT+7L5drVtJRmruZWYP2jmOV41Gm
Sl9v6EeYMqZ4elz1USB9BeKScTqKjuKU2YxCrLbOT8CbYNBmlVebnTneuXeOEY0oosCfCZ+48pj9
D/X/zyy/nJYLfFX8Lx82VjbKBhUe0OZxi732aQr97YCvW+fbouWcBqYUVTw5ivYM08cTK9O5NW7s
KtYXPxaGPDi+KCnm2/8Qdc9N+zt7/K0lx7+B39zgzwp9LoUeJtX0WXH76BOHbVwUnXJ815EQLqLo
uWjDpYdr1kkr966PMJpMVyDN2+CX1rS/jAs5qNX32qvwl+7gbpyX9wTbWHlXsxzOp6Y1sz5zDfSt
EfIGmf8lsqXvOEWxeXzyu1LNJjB92TpprQjY7XAfLloHvN1nT6g7D0alKOMXL5uE0oSM96gD2fuU
fIADlV11awFETu98SvcDl9PxtYKCniK84wahhHWOpP3YKYwQ/bZawcc3phdTZ8LKxRLLSJ8zUJvX
anNm/hccYYyoPQCeDTUkKROnzr8gDVxfdjQbh8jqw6U7o9pYfz1FvV6uRlKOmjUk3aNsPLOs5Kyq
qWg+yl8KvrAvUahl+hFy028nxpQ4tGoRVWGF3RbMi57kpCuO4cj0gdlCCcl9kMUeQrinTSjAOYD+
vIa0sfsdtfdKJzL9j0i9ZVJJwYQ5VH0zBlxNcPh+G35dWp5uueQqjSacFh0F6+MZZU7KQLmtLwkP
CKcNmcVOSqCFnNLDV4ubpin5A21BESkgpQle9+euzGm8dFZe6voKfzaecGQFH2Bs2aHVJyqVGk3n
Grdp32ucdtJ6Dlbud0gtP4a7et+ZtnuTvN0PuL09sc90p/BVBC0+qaibTUCv387NNF2/S8f3dRDp
O4Ul9S//+MUQTndVnh4Ip8/FMQ94mP+z4Q3lWY5uQ4d++9AZ35Rio66KzvrbJgMFxfHN9imL8yT1
C9Uf3WxUlfuZbEd3I/ARtS1ZMr8xId715TY18BiMkGhRDGA3/4OHQ6c3RyUKUzJr01fhWrcacfqR
w+H04hnS4ydTia0TRcz3gHTeNcb6RIJrAfi1KCtw91M3r/ftAtfQhtK9b6z9jhocrxj3/tQWOA9i
7dSPMTJgMMtpP//4sleps4Il6c46Du015l/JD6SPcIPWRrNp7SHAkhGRMl9zXDsXuw8MHQgKAUow
aW9tOR3CGgdfPFdxQq2p5jZ2Vz7/aG5uV+rvfhAmA1owXtDgZ869wLh4Dmkw6vepGoUE3Mo1tXat
kY5DEURTQSy7ZioqgYikZYJtnDSWJxwu2Wt8xS7GhDXU1bxTAdXdHRqwZyNJZTEwAmHlUDuVAL9t
g3Ka54OD2xfAxR76Vj2+o63cZ8jI5qTJuNGf44WSd4sYS5+KzY+0bFvT5+R3XZdmT4zcWPatR+6W
IgiEUekI5wAQW9jqBFDDYJZ9D/7PYZ6J5DF0ARAws6dus2wSfX/UhYVCt2nyiV1X1ttqywWYDeLQ
v5hof6H/IalR4tnV4mX2XI8Xy66toLmfaSphn4jEtRTvJIjYMVhzdu+e02S9QBwuyj7j+WUzU9nH
ASgtBDRet09GqeH55scEmpK3mecRr8AmFM3soqO0EFjsli3gofDCdpscxkWpkeREXSXLfg83lABF
MeQfISz5b88F0ZsYuxghxx5VPRcDvOTqIwjBD5UoX1803Wld2txg22APiPYHVw8CCctOC90Yi3Tj
H1E49hfHVncbMSJOrkgthNlvsX+tmRBYGiNpO3E4/m+zeJDOl4XnnjK9EVqrapiHVeaDTW367ZZP
ngu4yP1lhO7uOAv+gt7oIEgD5DkeFvfgmPnmc+rWJW8kegAw4jFfqEe0jGZCoONBZtBGD9BOvguj
l66l1xsMRPdnpVaLXog2e50m4p24+e70Bm9d+xIMnupwYDh3QCXNIJ7BV6Tz9Sge+SodzwAu43kD
pSN71fVWk4olFJL8XSiBTKZo8pic280UAstW/akTHBs0zPgNz6wj13NcuDE7Fsldg2APOxoSABLa
Cy1ed0oSIvYKco/5t79Wz+eB3bhXI1L3iTeTWBnJmbuWkrZbKRFB/H2mQfDRSEikFae6FItTcalz
HdVBr7u8bREb/GZkv9rJvmaqsf0iuTwbfU51OPxwQkRHOeee9xdxyHe4knetVgIQOo8i06yxvEUD
CXBUnhy1Lu2pqM6QCJHSk7jwguL6in+GcRYuGnTWRMDHkfd9BDLE34vSaTbpzC4jdLJSdlBYrWiA
JL5aYIc6piCrDcFJDsuV5PdUqPw5MQbTr1GONQRdTfdkz4HW3cZ0GtEssyphF2449uAeQZpjaXsP
M350iM2WXhY7LHQrMMe24mH7skNntw055u6ZlTL5c6I7fqq6Jz+aDkTUC9Z4hPibrJGcVywhMf2H
aEJXy7Nfd+LIxZ9NXxgOCvq769+cH6vjxYpEGwAUZgT584PHkG5CqN72ZUoMqv7EukAnhrj1SSzD
WYEkTH2KvgBWJKkZtBq6DOe/HEVsuMBLYuo58Rpczfv8CjupfFD3mWlqvgieboS+P/iGGDB6ku8D
EIGQ3LRiPU0BOG2+Qf5lvFNrQxD4aLxdzhVHBg5Jmk+rDFsfXhNQTyQO0lXU4M8M+UWJwKDtValp
dXaGbB127FZ8SNBjvwhkENY1WboadKCYfFS2XnJz09674AH2ZpJlPVw9ZR9yFEBpoFH7C+yr6Jwi
Y/sIALYDOB7ZikvFpMBLF+pecq4tl2n34hLYh/Or95Y9QMn8R17FA5oV96ITXIhWHQk8URRVUdsQ
FM42jHPrUYxEE/uMd2EUAl/IgIxMGOBl2CEI5gYVJXwfS8waeDTn9lN+x4iOHeUZmlq2dPndFH02
MXA3VL4Com8D5oZTVglvqBV9ub/PsMOL15LiXbd1i7mrXCGtI5o0nme1acGPzEzG8TlaTjHHmRvs
bVdzrbpw9c5jKStgiz47ZvdKiFPYKm5j3QHXfgkCm2KYBrasMGgsLpNNbcy+10mIqll1Oh0TZOO8
VGVZh9rC1a+WCNohPB6sUg7ZqaroiwEIEShxezDqTKwhMuh9l+sScrf1NsPd1cf+k3+SytysD6QY
+H6RwBerfa2pMAPJO/GLOFSJfnJxMQXjMHcbiB3Zg5dToYlANNqq+NX9RS3vc4WB0NWp4gwdD3jR
d2ePfC6MPZia5KFvnqGA92gM9Z780fuIOcSIB+XT599pLYob0y7H1+84h8RGFCsp+geRC2I/RZbR
QIi8f45hmrpKvNyTjOflx3Ml9ypFsyoMIJRuEj316+7jU+P5yAGn/z9FWAYY2e8P3s5xuN/qvJ49
5AMwHpUIN6H17wT11lvTyFhN06z4pDlspZk217sbEqpXYc9a3NN2zjo5GtAtpzC+0x54vOe8GBwb
u8F3kK0NqbYaCYy2drI4SmLNEXGKyc5FFr6bcGUb8fjyhUj/IPLMjQUqtWwAN3qU3fMr8SALjl29
YtA4coOZApXX9vFy6j4w6RENrfYb4OK3lYOy1pydNFNejq16bWTAnQciBrFahF331BIsM9iAl2kD
ZcsdCrxR/ZvxtDOx+bcQvzRPzLXklXA4Wb9gmaUU1kh+gwFAjTMtmb5rbTzZAqHLBao4p1huM7ru
F3neeV8C5/H619SEDT20nla6kuhMN/EYcZy09l/u2/EXpvsTAVc8FclkJWskhUyLfVLeRtaebJt2
xYoyWvFGllMsJ9NJGwrl1zV7KDH1HVfFUQwOhglkdUMp+APf4tFTnDgo+ACP3c2Nw88cfaAKbImW
iSgK9ik1sFPhy2RxyxGyiAM5Egrg/1cCLXkKx3A01FECXWbtnhyPv1wb8lZBH1tekDXwJrdvX3lR
44d+vKVMoOYdW2obE1HhVKlraIj9aJtxBhuH/mlsovZq8eKRPQdVSqziW0vUd/UGXm5dGFuuR00e
sZf9GqA6gZOZriJEn32CTZnI1sKbtyc9rp4bW7uHy/2dKwT+I2nhmRu3kbMmZuURc+7DDHHN4oTa
U/X0rWj7UAd1gdkWqufe1av+iQ2YeqYi5T8r6zw9BggDeL9Owov+z5vshX0UGu9DQbMrXKT3GZ9H
nAPIo7tLNr2mJok2R6d8LymuXXZTUmF1P+UrD+USGYIee9MrKhLw0GXhLQ/aHl4s1iqN6tdMIiir
36Hm2qAt0cH8qSCjt0XTircmKgFChwNdeN/PeYIZpCNIkQPFc0Z756WP8vGeyu28TD0p+TFonzF4
NGNAkedWYV/W138lKYS/42kLmpANFQURcxCt9w1GoHOW2siQATlI3qgyd92by0RuZDbM+WbYZJb8
41DU4rQNqB+f0mbVdF5DbF0AeXP6WioQugGtLqIb7vSC8UJcdRvhMWbNqHiX2PjqIQ4h3tYOK5Xr
v49HY1wHtwv5xOXmfOy1gHWdyNOBU4bW1UjJUxB5dPvXtlKlNbFNY0J+DTtlzmzfChYJoGBXe7TQ
dKDojl/Pq4LJNly9IdS853CES4jXbhb0baV6wWIpf2Vs5ey/WZvlVTlqJsjjeAtn6nN8CD3BvlAK
DvhR6Zu8ksJvf3dBefwieIXRDacOxCx7WcKyFFSmxV4NV4DYQ6M5qy3VxJndNC+T6bHxWJ0nSp+S
soT3es+PB+N0F3V2/Qeg9H/HQO57CbhgfhZSbHXnjcdaQKfjjlUPcSWRNgktNpjtt59oRPIcZKAJ
qyTL50sBcjMgSeDbdenc6z/QIpmTBo5+meWV37DExfNj7lPCl9ZkYLCxeZaT9+uhn+/GbbsTOp3L
IosJ01kvjTYN19fIbKJMl2qC7WYBFXlAdENQCtXyyMX114gD6ZeVFOFLLAQ4rBRaE8K8UDCDOSHa
qNtvZ5t49uRWcMdOdB+rw84UjjbUgrbRsblQqZiE/b+Crl7HxE1hZA6V1Ace8+Y6OXvVXPjIJk3H
9/brVPnqRAafxP8gKjKmHSnwS59oUj53B6JdURXWtN6oxiV3dsvOjpz+CHMyNfu7C9A23Ogxaed5
SkOB+W/gqFY9DMc3UzbGfGEXlZK/VOrj49fQxanE8urGUDSqeKXFtAYEduteri6x+2xeKn+7zSpm
5w8Ln0y1QQD+vhCm6Zdljdml39HQm9qJbMlE9kosIHJPkturXYNoVp8voVf6EnbJaYOxhQ+paj8M
jwY25npoHjkkKdYqAAsv9jQPP67cDV8wYNb8pXa4+rHBRYGTgAiLc0qQgD3GJcMSGtO70iNAjgKf
gBUGa5H5+voOM6owwJmqiWjkxChRWZZCSWr+ug9NlUT+pmsWF8KLDR2QADkGhLVrp4dnQSxM1Zy4
ZclEl8kvJ0xCsgPfC66SSvTWHI/SBS73WSgoul+vNfbrSjef+LtvzMw1IKvd1up9JzYCFv5b9Hou
eo+EHYDvWYy7t/Xb1w6YexPu9Y+lQtMvuJdUaq/v+hdPugB+VgssFP3CBRNxLvoCYLfmLfG1AXSt
sDgShRRakwJ5nEIL10s95bjNIFC8J4aV+q95cWQTOhZ9ggmj/e3bFrwpfoIvJQtM4JF7i+EEiaLf
BIKUVZPOO6yvgaHFmEOHoCHMBW+8rw3hcwv1ny24Zv0URAujQuX3C4Ce9d95ArNttS+xMHeRnpPf
iMaGFOFHDEY1lQ4Dwmgn5U8rkWBY8O+yeIzQ3xxHg0tGVYmL3oOx8U8tPHxbrQADmo/YJcRNwq6C
7MNggCwjynzR01+leY/p3hjjdS3IK+gmnCTs5SFD1OoIymobE0dK+eSzgkBd/qw1hN9cfxoRBOLV
e67mvm+ELCUx5KIBi+B+UM118yaR/wiUWJ0bI0+0C3+sa6z8sccDO/M4lmdu/mGUmYJ4chCrfDUM
4EF/Uf6LStbtBR8tA4JOSVW9nOvBtn+/iGRt5cYLKjQt2a4jYq0O3QV5WtNaWHAf7DgHoiD16Ogf
ogsnfj5PSuiOyfB7fZ6QPYrKkgm/KGG3bHk4CPu9ERoLzXURGm8ticDiaQxpHfsD3rNXa+AXWhww
woOFNHAw/75QgYb0I+r4gksJ6RuLWsGCiTlWa3fCi12J2JnFd7wBLUbM5cwBHtN2p2Pn0i9CmyUM
0BsBSHTUPdMKf/g5VUUi1gm7WTWsBh/40Q1SOEY4R1vhkmivyVsLAAj24kHbqbbtwaRzF1etAShf
amosP74PqWJXtIDN9ur+6u0jLtqamlhejXF8knM9FOix475FpeucN+nTGu+aeW/NzHab8g5skY4e
owHlksD5SjrwZfliEj04XloZDK8N1eS+pVtxZstNjvWhFGPtZCaP1igOffQhd5H9W+9OAzGRRiAj
CwFIS5NF844LOdZH9FIJhjp5yTFcX1rnXiX+wM9aBODvT12ku5TvLuA4A7wrWYsv+Ic+/jEoZlFo
D2GyyL3uy6ENyfZVl8FXG+4LVnKZ/l3VjTdXdISeJdIN6GIKU6XXAmTF0vLd0xmondNcJ2L7WVKt
rr0EKQMpTotmNYv0j+bPZ0lEH7sg/46GaFK3PlJxf100KXoq2/UbA5GitjGiWLMaqh3xhxsvORzs
gx+jw6+/UtxX3y18cexKjpzhe5SJuFL3Cct7Np7fZNVt0zks2gEpDjS/yrGzToCUKcRoQaEsW57n
7nOxyuU4vtJre+Vi8xsB7bGEOeeTaKUDMZyGGpwB7weHZGckvYhtl0yOJqiOJsKK3Aos4fL5fqeu
ptC0PBqc+MuoIznOjDBwPLS6JiqHOLJB0yWmHAHZ8lIRLO7+Zn9dzr0RzEuwtw9Gbq/ybkWCALOu
UtYV7f457MUWk6ypIpDpIuSh2aaa4XYbzZ/8QY5AYuhgSHcNjdvRlBx2AkyT8pJ/ClG89HV9IiP8
14tcYWaWf+7EeXNp7dmv/FJQ1RxOWKlb2gGcaf9GdzLQb1VAJ/vegvaTMBWjC5tskMcaQquKoNui
nvqDYmjDoWrXDMGNxAYHmKcuPX/Kn7WF3zFDgfHJ5fFh6mfM4N3Doe7QkYWg6s36nsIzBivxyEe6
LGgCcuvt+mwwSYSD8gFAsUclFVLEtughbNo4rebvVpuqXQF0hnsl2CU8njPIE2/zXlQGdn01Xdo9
4hMuPPyb8nrmTyb6M4x43X6ULUxq0y/jQSWLFDb8N9vKekfcUHDdzchs5nw5/5bQPQJL82hBHFmV
59SvOwaF8wZNE1Fc9wMToW71lkfaucP0ydzCTBiHo05dLPAYrZatclVu8ncqc0dxO7bUl23JxVwe
kJTTQGHV0R/WjmGljMK8vMyvhXIWWTuVtFb0VDzWPYphaMkJoLBFe+AmcB08QD+KWe6wZZHf+bM+
dDUd0FTnaVgANdeq3d2kAJ4cah8mDB7ks+7Wav5P4MMHCA4iQ6ojDLRTxFtnVEz+VWDbVg9rIrnp
4DZCvDa9VVb89m6g2D+03Ux6R3XS0WzPzd478mmnCvT5uUzLj6SSCQSaF8qXkGRu9zq+nXxeNcPj
E25diPMDjfJSvChpsqmhpBbGU9ERnShfzmmw2g8uZZ3LpoDfLWzeNihYJw/VcgNnNKS38yMrK974
7R9wY6CZXsp+Ui6+yy6wMMmN1W3hLfYfoZQ/vjH+t0wQ8zz+l449VVWFmy2HY7GAK7VoyjtghCCT
Y+Rle5mNP05xlXNBBq58qMzWiwKrHf2w5qjFlirQlWy3TxpOrmN2Sgyr7m/Vh+1r99ionj3RjCvs
q8Wfqr5qpWrk9ErcRqufE9klFBFcnOQxAzJrFKimebab+vU90U2sm/ftU0pZn0yAkIAXWS5VgqNi
KHChfWQQPA+cHc/F7isPCNwY25m2dRLBvPczU5We/iNYG2czlOPrgTJxBzd8YejNxIZ8eSaqawVT
ZxpaKL7JAItyySY6C1y8Vr6yTwdETZaHKIzVfT1siXRvEDq17OXnFEuqssGg82ScysOqIV+7dPKw
2UKgNERA24HcUUyx4CgKpb9/Yqf6v2IHeAMc9kEkoJuR8vsPZtR6A0eRgrkFvarfETNiYpHz89od
jFzZEXixfIyxV1uA+W/Rp6yPSoi78j+/GC+WqIi0ZR0Wf+qvm/S2iNbdbFqfc8U6OIfo1+1EVeAp
E00cDDFOAMi1FamyA5TMh5gEU42Ims7pIUyHizMNWcmzMfhrKXwkqqqP05wTGLuAVpFsKRj4BC50
Jj2uJEqiD8xmaZqsU1AJo0XrHmkrGyOa1p8YqeNmdQGU6R+6TZVk/CpXQ5KkVBCJ32gVTwEt5DU9
V7EbTCS+MOeM6+S7/rwagaa42AnHOEV2/Ph2C5/vAv7Z7j4eCq8QSdWW3UaurpuRv7hXFLF82bHn
Ewo76hyNy/rNA8hRloh8VNvLX0qAoeQHqME/OynHSbFOQFNaKwZnsyNfQDaU1s+gOQUBhWu964Ay
/FyCj29T68Gn6pFXZ7DndVHY0ncOXllfEnbmnt5475r2lq7JwIjzRAvRvDkh7jDr6pbc6rBE2fyk
qGW+/p2Ztao/RR9Eq2h1kYmJhAvXXmYrC/eWYUOyP5J19HKVykwdaF0N87b/kzr/YG49asNjkir+
ljnp2kTHDOhUyl204W4kbXrptq4G130vYgMvtEB8z+wljoYzOzmp89uRF3e0a2gQgRCBafheUveN
ySSHhn0v15Aj7d8o56MZ4H67YsyLaHAWYhK2kMsvcNH6TibxjXlxoauOfQRyJu6XfI7X7/QeGVMu
mR1vkzKhnQ1x+mGvWJj0EOBFTVtfcHLUrI4tFjOGX2bMVMnNSZefTxghNbHNL22PYZgg0uOnuMO3
FXrqivfG0PpFEdOdsz6BDt6HGg5rCxCELOYhjl1aThiDjy0iRx/FUD8vFxMtZ0GQ+t7lTS4VGV2a
hD27V7HPCUatauJ6Un97Jcyhqd2bNrPfuYrWV0XEHNBmZG7rUZF4eAXHJqWIqACahRNp7y42Ze4M
iGUIDa2MU1svUbUkgPwBWe11IC2VXJy6EZIQdohyO56TWcn+Wf69uKgTsLrOUIl7Kx2KE2ZbQmZ9
JP2TgfqtI7Qr+Bcrobv9PY2uq0lWGSDl2Jp8lz7hcDhzsFqPFj8tvdssME604dKfQ6HJQGKatrnU
K+Z7lCUjEwTAOi//zBL5Ucipra4ZjTccHqjlS7Km4tX1ra1wuSKNEL25Sdd4lx+7UNZgN5QiRp5H
nuSPh6UAkFhYnl3U2+E9YVKxgafZKZx2zB+y1Ts9uyWPFDDSdgpptqPa6UCvo8wNfbwPydYAP80v
ggXtxmX2azd/phfqVfXvRCw0Ej2sBiYYv8AMkn78at4d3qnTIoKSrOeLytFG6VSo0YMXz1Al7Jei
a5SxrKGBFaav+V0yBANUV1ifQyM3nHQvnTwAUxk84zyORPggOWmvB0PPPX6/G5TIYCKdunfIVG5k
Ubz7MayeFzPqYTLuW74F1z6qxZrDYhrAKyMzImsrrjrdfTVx8fLafcbL5vfkBMVjRdmtfKkSkpUv
cfGyvP6dFO5XZOTa6XbVXYWRnUk4aB6wnX2H25+eDImnOrzOt6eXS6pUtI8uY+dFazE1uz8n5WG2
1QLKsxfFL+hDwDtjr443vE+ljSt5cC1OzpPSbwWIfGPW9xryjvrOtALDZEI7vbYxY2SChoU/SKSd
s+XeXdKMB1FAOgfU8Y9CFopayKua0is8U0XWCqOq6EEyG3q3H5sTDmKRcKFFtwMAYkusaIeQqLdd
UdZjMQrnoEopTpgt9m61Rppwd/6bisX0/J3eSBCF4exHChei3MJKKKLliVBEHP5ajPbBXxeVwfPe
eP3+5cAv7VbeujUxyVKJQjNkFBkhLIZ7Q7AK+goVHaCItO1mSM8++mSs1zH6vlwznNsgagOkW4qX
YF6I6H5S+O2aVa1tNS7s1w0a/UCjaiZmLP45ixZ56sRUOBksOayHl43S/MKnFdotTEGBxcRDdWlJ
xLMou0j0X2I223PqCL+vQQ0OmJOMCBXntdvxs1qD4xrmaHfkfNpAH2jeqsSOE90WDNpAKBMUdtfm
cTPzy9i3C3bfDGYhEXHKWgW70Q9mDS1bcR1oKzBgNMZKWmGu8ws9nMKWepp1TOzf1qNt6vWInIGX
pJzOLI8gs91og7TsrHS9V0DvemYPNM7K6PV2axlONNdNnCSUcCoItvO9S6zbhbTtTDdtavc+LBwe
dBxe+HPuFoeyqI3wjadFRAdAha45sLF1zRMZqKc2sE7/VZD9Z6T26CnlL8eix2YWaF7695Ji0PyS
bqaH5V+uknkWvP6N6k5inX+DHbQeycqPh2t+vCCFMJIOHYJ4uVFT7u6wd9EKHeP3QlUP2DSq736f
K0sdlyNNR4L96Y2LgNOl+syLBTkF1JxMyq8ut6NCwzsr/TbAAMZh1xrZupauo60vuxmhnuxW8J6S
SX6reGsJBP2A/KYNRp4SJTR0CSsmaEl5sHmsfCGfWlHeIerTC0ZPaBCNoPVGsb5iherzAy3ecwYb
OrzM5EgoXF8YSR5I7h/NOfiWAfwHKXYwABVjYy3vScqEfiQGzilZcwn/EBdNoGh6DkqqcQRP/q69
SyKo+TYr/IMhC8IL8Takz3+IdNJUrHfomZbfUc/NPDRARyWv33eeM1O5Dh6wDJ+2cThNgexsqVuV
i0Q2RTwUd+oTFRFQ48QOWCXrOcZmsr9QXXn6qM19vhdCn3fmRCZXe+CQX+1lYYfAk2jHyUfjIosy
h3sfET8Cl/y8ynpOavQTs0XB3jjJNNtPjYd7l+TL707wZNzwtpWQ+u/7jhgnFD6+vDNWuAgWpmpv
tX6/891pAhgHAdRM++c8y+ehcLIfJYvIrsQrtiQK3gzN02qRM7L4BWV7mzmPoi9JI9h3ZCBJ42sc
BRp0jP8Zfv9nyyXpnMU4dPxfZMxMfJgJgqSAZGYiMjoJI2+CEaLGd7pievXpv+A7MiHGCJnpKqpP
ex378E9XaX4jtkH39TauLg/ZsewWKnJJvRj3o04HAPE+sbMOhKSATZc5b9cMbBtuJr7C0pVWnwTC
JuuCi3UVLpoAYKZpuQlB1fr6pY1whlqI1BEAJhCiRBGexBJASugv62Azb7/iC0VtpVeXiK0yCVew
N8SkdJekZj/jsad82iF7YaHQQBsHcec91e6JcrU3nPsbF2ideKY1fUkNXln1V5v3f9q/oawGY7sf
6tclwpd8WIXzVZye+UXuKiQjOANDVaAnyMsIgJnZuDruHfi+m3TEYtkka03fU2ooaggX0OBbnv3X
tADw9uGXfRwrJVhXkxYToaLa5np0ya8poq9DvcE8qVacxkCPEM8nd1Mt+RLvbMTpMUXjTDRKZV64
LqQLkQZAi45HMKsM2lj81tUPL42lXeSxeWkWWf6B5DZhQmg89FvQzJyp5sHq/ucE6+YRI3oxjWBl
l+QF3ELBEHhn6w8tVQvY0gDzC2WWvg3/OhGwmITUlh6WNqmREL+OCVEkjggxiYvCaantwCT/eEZW
9A+fRgc+GNTpKSaF5b3/OsEbBSB8DfXF0tNitH7oA4Qs3caPHM6tsEdnzzoCb8/+Wx1MSg89r6Vd
DHFMEP58IqqzqAkt9nguI+ThqFRNgToz2/HG7i4g1C/rPnoSSHBa7TtUwBXZdMjSw30M/WlmSDof
1ANbBp3os0FzRTqMFy4N1YGo+4E/VN554BQSCAQtOz3wfYUiGknzg6617tB9khQjIxSAdZVw5kG4
lJkApyPeXc1RSHOIIoQwbZLZI8UO1qp+csbakcQEOGhfpyPYCK2fEVvRGvRXhS3FYLRA9ewtg5u/
kWr3OqjHanmc0EYKd1dn9v8BaYOeJTymxA9+ejevKnFoNGaVH44ARsp0+Ba+JZX6K7/X8nfoNzPg
UkrBDHNFhHR5mLOnu/KgEnYWZlWYtO9AigDIge3W10Tpe+hW3ExcLrGNMd40FRgbpIJKp20vj8Ge
59S8pFhEqly54AgUe9A6gW0jgKzOGqUs8fsG3D/hYTWIjzBos2s3AD2HkjQ4QYgqHs4Pnr5f1I8K
pJaY3yH2wrw9pOzs8l7gD6WRmiwsmn3a+ZZc/68ku82XqWxt6VZ5ejZ4r//EfNK39qk0AlAZ104C
9NpJjbBGDtyw+x0RVwXNvbgaEmsRWz5MnZd7WqzPhAsvvfZMZbqui+GknlhBReQ327bDb19sz5Hn
C3HSWwMWeSOP5a+lrVjeGVQRV/RJWPpXLgl181EVK0dDcvT1U3SF0VxDpuYjK20zateyKskrp1U/
31+bCZkttnI+idjND7f1Iw1qD7FSun7KWq9kIOXDNqpYKFD7zNn6wCCnWlM7Edk7/9cZR+cdEah8
ard9pbgIy+uyKcmRIrymLpg/uX8Q0M/uGyjOvOwBSkaJPz3aV7nkK28caZBIhQCvliIRj8DsHEJv
KR9avFJeVTiMpWl4TaP4X9465KdY35P/1NhrRsM5Qj8AoudBFrdys7YNcVcu2eSVliSIqfCOLtUB
66CRNbDtqYzm+pAQmQnxO6FhCHJ1pILGaOZrHtWDl4BY7Ku5fbSxDYHYxYl8rJmeKjuYhVIuIMAI
jkkPWViPT+OYsXyj8Db0GyeTfr/LBTeO4UOEkyVcmblElJHlaSktWEZxcn4KkDu83NqNKBldaDPP
gwDed7toNijB9SCO2rZtVW4d6tOigfmTLfwLQ1Hl3ZA6zwfkGbgz3fed9sPpZLovZQ/KIZowjwHW
DVDnLG8P4CnrFOEKjXBtApmQBO+soJX8C45WphmFJWn5s/WpLgRImIrzSUIk1qin+dK1YCK914Q8
Gz6WRGfe1SE8cIsNEFo6dRs9M7O0zUJNlo2x4EXqK2EJfLIEXT+XsFKuNUxgfvTI5vVelTMjCpOE
BaeR6zl4Y1QamHYAJDchDVGH+Ue5XeUjfMaS7UDOglEWG5j9rdsu48F12+7SYGzxA5XkAJJg6DPa
SYsWyVVWoHqhW1BZPW8j3sylXRCjm8+mfZgcIJyRrNaGgkNXkYWrivf94H7g0ECAAH1xcFT57Zbb
5J006p7v1cTYqFUzPxZOgGczIawtLGiuc5kCuC4lQIazkzvAD49QuW96YWWc5sDEiMOQZp3B85DC
ZIlevg43des0jz/bi/6UhkWImxSBhITPuV1W/EMjuigS8ol2T5iqQa10S/wtEkXUthltBb0AWeev
qzRGOYf+JXTqBmwoQBlpu6kSJUvrR+hmO0wj9xfOVqe7qiH0HASsto6kTLljS7Uqy7L2J66zHwHd
9sYyvXwgjrx5Iv1bmJW7HK3X39HrT3r/CmAF9ah/LpayrKrNmSDOw/yYMf4D1pBDlILu3/nILkTZ
+cKBm1C2aLtiEELdCdQ4IyB/IrUugDhlVcQD9/MfTv1fWF98OpZpb7LO4A1f3QXy+OfTrKJIW6B4
O+WNntsiSPS+2elDQtX8FJOitn1eQ94YSkmd9206Gix+wCfTxRdieIedQ/0U5ZtOwUJv1ymUxRjU
pbbe73h2k6hQGMy6LSBO9gTqIROy7LOOBPI12RrghTR7/V2kFDWkQK8EqHEQkjlnWkiG+ArrzVvi
lTx4FQLEUvMHfr2fzlDjWPssyZO6MbR4m5v49i9uB5RtNmW/ahU9NbmVL1cRXxj+1SHqciI0mWty
F55wR8VOokPjU6rxOjrc4m10bk/oOOfHWJwWL2Z+zkh1e3JUZhJR6P9lc2agjEA1VpSdYhz0nMd7
4Pk1rS/X+gp/+FEpgbyo8QPWw/5gnenFATLX4w5YQ4skDc2hvbTIfDnscU7Jwc6BysPFAqmx5iel
wSI1MAI0DAsym2QsGEikpHuCmJyvqwLpTeCuW5Oh+pO2SA6NMmH27kaiE38pYntLnsVvvM4NuTlx
7JJXu+eYA+vQNpGAiGnHQjaHxnHclNpz21iizKkk8Pp5Lto0JiLHR5OsiEpInHSuK3T0Eq4oIHDI
1b7i9uEkZU/Ib4eBdo+B0M063iGH82iATM6VFVmeKc34kvkRkROhSxlm+XwB8KZAyMs0Fq/It3km
Mq7Q/AWqqY/rJqtK/Qqx7DO5JREMMXMmyndJ6x42M6P28WQ3h8mESs0glCeralOpZNLhz1rqlUQl
cCCh2M5DsaZRjJNj24XrPAOH02KBWrDTTNHRzP7jOB/DGF40QlbFbKwTDtU13jdCLrMBVNzKZwwt
Ix8ALvPebtQxSI9qR2v9l1Y6Li/QDFlvcDFeseXC7KaUQccbZGbZfuT4iUEHzR+ZRdDZwIJoA3kH
EvYm+DaMoQ59DPeCCLyGv/gmwCZjZqlyayshPUYUVHhpeA11CgNJofi7dHZTged1JF8FCRY30heH
ScNW2COJN58Anfz8M0TbE/bL/PCAwsBbQgRSh2fS3SslSrsso0gRe0v+UDjW+UyOuK/pp3+t8LRy
MHdj/NMiQSXLIasRPy/aH7vFm5cyxNPWCDulNrhjRMRtO3/PBlyYj9pwBwzFuU6kAs81HfN30ZCr
75X/kDj0dAb3ZLSRJ3+91yxZ4JP+/rU6rI7+LzTWMQAE7TNrlNLSHDMKV4KPUojIKdBLbN7baTpG
faPGXxaM3904bSIMbZHKeaYavYmIAGmWFygn4jP8C+YmsV2y3fe/+BkOhg03jRLXH+HfI7hc/x5T
g8kEQ5vsXD9SHe9P303oMnfd7NBS0p5tFZoJLRFs6F1v+i8imhXVRuRAwDoIj12csC9z7zS1/PPd
T27IsM/eq+oCfbhCBlOZZfPsZ+q2/xbhuoBQ3dvkdhCOojyktB/xB4mLGTldL3wYd8aFbXs6ICcf
M9ElRm+wBGdmYGibzKwIBHGTAmLllH4Wu8gPpQrsvs5vx0L3hcH/wwTHr292msSWwVCJp3BChMWT
zQZPqNyr84zwHZp07v/KizxtKiOryk53CXCdOAk4w1dB2Xf5ZDIk0vMla9B7r+k3MWDUAT1V57LH
KIAeoUIkEaPAnf9yZlkuktuG1+/vLom8zou3+MfyW4BCOO/XxN0NjWb1FQLC8HjjEPE5aq0aQqLU
JVWHlgNXzX6pqvxomnbBNvJ398aK2omOXCGv0hY7q1zwndTtozkZBVckLTwbHz83KCW7D/OJPS9G
yAq4cJ6ffI1s/Sa4CqjJWiTrBkcbUZ1jeIinfo3LXD+dtssAYhUTzvItDvz3+gH01sULV7HdOUA7
ntZbwKvvWJ3D3bF8+H/m0QLOG+rnM/t/u9b2rXVZVjy1vduM2p2km9vP8X/7OPIl2rHDlOfM0SbF
Jr0yjAp3y/Rtvds0cUt/VlFg2RVW8moINaUQlftQ0qRjZISjRdLAkS2QqVcQOs7GNsrMZGlUlqWT
8h4GCwl8SIfMqBDM4HSzbPgZyw4UM3+NUhBY+RmkGBFTtbKppz7nCGTzdjmO+BBgMD3kHf+WGdq1
fJ3V7mYKvG7LSFQIJ81PUY3Q3+rrsMmf6e0rZVdxmkgGXtkNdYjZl0l9l5aMBUwFBxtonO2QcOy3
jaDtg5xyuDr4+BovC0TEfdg1/8DkUwNT1lZn1baK42mR9Im+SNSu795CEXSFfRDdPLB75/rn3Mer
l1Vu6CdsbMQWgYqTIrEQiAZno5c4jfmK1pT7/8ngd/r1brvLbyIlZMGM+xm6eh6lmpUhyzVeCKyk
L7CJ39hU600kDgXhopYbukzez8hvDevJb2sXRQuTIuv8PRby2mtaqD1U3M1FfWSQYrUZWlzNAbp6
TXtmH73+GBt/6TJc2kqwE1vvkHOBacRdN4YidUbJGxTBfcXbZRC9qztSTkAktz474hAmOZmo3lbd
L9FqFvzVrnLXtNQPLWruUamgycLAVlEtyItg6HAzOiWWys1LL1eZmPCpq18v44ipOJV8LxVvACpE
u87/K8Id0vIuXPRifHUtmlIEUchRrWNPD90AECXFErb5/W+bN/uhrbY4yy+TpfQPu4eDOTYlLIsk
zvMMtyRz3Ko+1eoeiOg2SaBUfBs75ZHhkIlnYAfb+tr3dUgLmErQLcC0YE39ZsUp4wAZuXYzKybf
7+rQJ4X4LQqZ5/I87k9yz2Wkoa6V4VUHous3vB1syrHk1lAwUADlY0qaiGuiPhTJJSCBYgyvpw0z
tBbbui+DE0+t8vh/MIKAz2h7o5LlaGAdgBjW2ZosO/jVhxJAuTfM06dryz5amQJDAvyvLmM47iY5
uRFsdqhDaPrlBIk+rTQcPZ0KF1Oyaxb3UvI0AXrfzlo5bUYeGPTu92UY3841J/UuIL9GsfbTY2Lq
XkCD6jOtPvqZs6J4ldviw5SYlZQlQyYm95qLlD5xqRrGbiCWyjLTBwIaoiHPejj/0yq9vjz1Pyc2
PH+Ih0W/xqScdHNlGR6hWA+kFlvN4wOAi/UuFQaqrIhZnroiQTFzyvmuSJqUIic16+OlVRQgiEdB
fOCd1Qi0vNYIdBR5Haz8O62UIkjf9mD0iAmMi/uJWBJEjVh3IkeLxd4TkgURberiD6W1+jcsq4qr
SXMJ2k+lBwpirNo2wLUhzgWRAgF54wVvicgIwNwMLs9Ge+zzJ9Jx0+A/J+Jj2hs3jAQGe0mHVlpn
6hD8kCrCkiZpr0zgolUE4M7W7B7ME97Ez5cqZAc5Uir+ctXlGZWaMV3nd1Dk4gn8EUef9hquPSX1
mDn6SYmNLTs6ORbCWjAoOHWQ0YcpI190ZMveXJQtGgEpzg7aCLbcu3EJ5TH4dYVwk1Cqzhe/BIC3
cqLD8sueVDF3aI1URIHzoM8MVuuFTwfcjFYSx+noz8LSE+CN7TOzJCorwfPCInNWohvjsZquHetj
h+E+n3yEa8e1gJbn5VO/VFN/KjHp/WQ50qC2LHTlzPUJS0v3Q3L8PeOClGfNUDYWzfAadpsnccry
L3cukea0tryfFEI8bAG6laYpVkevU2C+Zid6b4KwLLiS1kQjp2xaXlxFtmU1wvqc/rre7BpBpvO+
j/kdhkUlydkE2OI1yegrRMIc3632NYrPebhXaAz84dEDHXl82OwlmySjaFCeLbZc5bW2MVV5vVL1
w1SX/fyUZJjJvlrICLfWSHmD/LAHAKsj2SLkqRk2Yf/QCiHngBr6vwKrZXFth7ijta+CgBNlXy8G
yTSnG79pJvVdBFlkmu7j3tF1j1XoG0eZvnOKZoMvw+0NNcKSbf1rIWoF5vD/7bcpgvU2Ing5hG9M
Uz2ho5/cKEsOQX3xafcydxja1KS5ZxEq1prvocY0yh8951RI0vsXbxzAvX0ZB79WzDJxzB06I5c/
fY1v2QhoZJewg5NrxnGF380UIUZJ+Tk61QvM8w2/E7qyB++muyiYnRtlkqFAyPxduAUZv1ZzdUZq
mPXOvWlDq1oeKbV0LBwa3ANAdGFXfuWplPwFLc5cIqLmcLoUno0II4pdlpClCAKzxgc5jyHcKnDH
dRLQQsajX7MzuQV5s/Uca/4vu4Spr/RdBbsqadWmXG8nCGadFZqJVLwLl2qFGnd7uSnYZsjKXPth
ByJWcGv4oylEesfp+tSFwOkHgjr7Dvn7EHzWRNq1x9k2KSYXl6Kh2YsGfmxU9DdtOyrUK2RTRNDt
M2MZB4ms8IA1i7kNKRaBY0sQgDbZAHtVT7isLbMQLN+cWjQ267kCCOnmURZCO1PUf/bqzaHnW6Ed
/56z7NqCbFfSyrr6CWhbVoXzedTABXUDyxINTiSFgTNngaWjnC2Ox09azGVuvedlD36KTfG6pcBU
Zfoq+Z0eqpajuhvUl3mqs4fI9FoLaeXLYRI2JbbAOoojr21q0qGg3vvvkq8gN/nPdo+mJYClJZ3Z
dKGdfRrCjkeTFeP0AnaUYo5cU0UwRyR6mmRZGjoFUZZrqageTWnyUNszefouEozTcpLSAIxlw5Pf
Fgk24oS9/f3qLzI9hPSUeNofmaH+iYtClvW9qVnaKdyWTRA1Iot93+WmW2fTZJ+rRoX97YCydLJw
XNi7UiS+y+wicc/a58/d8cv4EHORr2v2ZIhnyuifkt149FZiPz7wlJb62Qv9VIw9otpAneTPUA77
piphUz2zpiPWft28pncSil24Rk02gmjcFRt8DZhNYKoCUDjHps3etBH8xBs8+VOMVd31gPpNraYW
f2jEUfHR5sfcsIuoRdCX6kJMWSeFDUIegSVfv1Sf6J9KmZCJqbsPiFwOvvPJv64OQTbBPDJVNCYQ
LibUX1fj8aPzp2n+0bfhhVqB871ih4eOkUxbL1vz7K53LKTmU9v/gQXaixhrU68XoprJHDj67JyO
McfOQ35IomKnN1FV0x9gskwnsiYzGYch/ZqMVb4eRBvio+Xf+afgROJsedYkqUX9Qj1mfIv1QmDU
MMIweme1+2cIx9WkbwBLhcWBJlu96qcpjlq4rvKy1lkB6kn5ThLEC/LZQ3caiIn0GC2MPFR6YYd8
ba7RsxZAio3Af/XceIAmwR+uVm3Pd+Iy4a1TYbtrzM3LC7cN/FyGBfwtXGYZFSN5O6j5zZcYvteI
iOrZhF3kXpzCtC9Td7NhbZEezmCX9m44tZpKwkk2Q893sfLY9Sit8jh6zeSvB2SOpa/Iq+UJdr3l
kHqhtWuySXP/vCL4HsKDPKnmLW5HX+6dIj/ieIjayLmKsRjz0LBT8D0N2ovlGusUsFrLA/Kz2S1/
ogyoRl7GmQtVM4pVHR/0DtBc4OmxXQ4uJVJEL7kuDosLQwC6jwR/G4zOOAOzC+vssVnJw4X3rgK/
0uxejflxSStIn+4X2KBE/7LVHgfmlPgEnc3GPrI+9YUGEQ2AyThzgge/tMypnWGklqX/v6e/yi3W
mbwAWVFe4CMRjj++zgQwH4P+Yn8D7/MEAioFKgNw/7D97P8oeQbquD+CZeN4SDlK1qyijoHGGSZD
W6puGhS59iGAhtok6N5fnA728ojZdn0VVnTS52PX3JaZu3hXoli5/TsFTnoaWJN360t1yuWRs4lT
XZSAt7G8dq2VOIhPOmBmzB3g3I6Ow+gDRKe1u16JB5j/DmPXS1wwC5geXDxGy0Y8jUV6dd0bL7sf
QQCb6fm63ZvzwVuQHCtbNq+MGjTQDfZBQ32qzDeP8xXqbSgkrT3VQqFi6kOQ2IsGkfVgTv/Hg89g
TnAzuBNU52DAz1ifLU6RSBmpv2jnccCmm79qiOW0AA0yzaQsI0yOjXLB6c76wwzenf4Aj2KNyI1f
T4DepNqdZFLDQC+3TAQVQs56HqZ/rePOVyyLuLtKMK+hFvswJx05pYctoq89oo0tuyA88d3mViNb
i5WFx9E4VC63h42U1Hb3xnp7lM+q2U/q7jaID82UUTWUtTpZkNCzHiIeK70d9P+AZs1Kf/QOXlA8
1fkuOn02jWtpotD1uIhd64bfZvXW0D1xVivl4kwKrQZI0xsJh3JcDtPeGtyKEcej4hlep82/h9Z4
aHd2+axC7jgStIv57A/lkfcCGYAV/E8v7XNiFN4lECIv33k2o9yLtt10vev6RS0beqU0GrPdsavZ
Y9UTtxEvwGakOd795E3K8B182vF+aiPs2DBRX/Rph8uYGP1Vq+sA9N/9y/YKOaoJay8JRldbX3jA
YEl/L3str55+RrG7NDZpqaRJALP8mXAokKjMEYPKJt3dAmgzjYwBEQkO3dgyhHA5SfUAq56zSdU0
iUNNiIKREEYLpB0uByzJALnUQoarfsyORyFoQU/DdQvTPaQRBgpM0VKg9QLqnGxAai9wpoVdRB2d
BYTj/ZVXwqT+04m/DSzTAOqfEFpv5lVQoHTCUa2LGCUG7Wdf6RMk/vqMRhg3iOYFy0fsmtZTddAQ
6x5I4tA6NdTTrQBY1Vp/VRw+1l8/uib6e6UhVNftH9ajvzCEGsgja1rn+4y1Q3N00l541nJjx20f
IvvoaOVyu7McDEk5XKbwgtptXcSb75m4gDgtEoNsucsHl3j5u7GtctEajEg1P1P2UlTh9VhypSK9
tabR1eCom/a4TTrTr9krGdVTn8AZPKhKU44OIcEBjcPk8UydjJKFoywO4WK95rSq5f7Dayj1GTAN
ACcK/tr+TrMkYNziZo2fM6iAUOxAJ4vzfZ30JZq/9Oam3WSJ5DDkaYlpW7riWWvSVA2XFVp0BOTg
pW0yycfuPSMwhczlPiMmLRUwzfRffg6ayWH2jPo8o6oRiHUtRpNaInjodWv2QkHj+6mQkX4CeNSC
tmlYa7YVX23cWXTnwPY8PrTMhKn9UywNMPnZx0TLYuXYpKRBf5ncsIEPMpnjmSKY5bar8QoU5bP/
ahFRCdVGQ/Yr36UnCfWJCqFQAfJBVycs75CLuxM8Hk07Asi6SO6lUWbhYuZqhK6e60Uc0pK9IbML
JRVAlUmMAnDiF//DZWv/aL7Zo5icGRHpp72BlT/no+FlpzTfYFRtqVW/6aQlG0KwvU6OX8Qe4y2N
Fm3LbEubkfGG8YiSdcau+qSL9Q8F9KokwaRMzl7c8eaKZOH8GjmbP5Vt3c6YShPa/KG6VADVxbFK
dlnhxcd3+Ev5m3LyCf82eMF/RNXHZWD67A4+OJ+q9vqmA6TM9qIMRRG2K9xDeBttXCVkxd67iew6
B4pNpBTfctOwmLCv2LmF5foNWmp3JzrHJs9BVSVNGibIw+ai6YyhQlVDSesehtqfDbn8n37SO+FW
y0GyIUGTEgKER+DLmYhAU/mdH0IATq6hvViOuUaTbSvLGnP70BdI72kmXHt2Cs2n7cu9xmQzolaS
idK+iv/+ZYnBhpwKFOm6NZP6+PZe3D+4SWUVfY6egLXIxQHGhQKyTuIhX5usat4+IFdxiSEv9Zih
nQcofQcqBuBtarYPZysXsBREJvOX0WKwpFqMumEwoH7NTXjP9Mmev1WxOSr58L09c8zb8f2Q+sVL
U5fM538ScLIaYUCGAtlfHZlRY2Xwk8/AAyRPFcxy62yyvXK+Vvx5hfhciEeElxGyT3oJoWUgfEvi
os97zGRkIvOlMpeOYhjPnFPIQu4IDbwrSdkXZ391wpgVQEJTbr357r3rjQJIjLpHJ9G0ExOP/bg3
E5/CxZWtLmrg+FsbNlz+3MYVNoaQMgFzqqPup/MBNaa+qb2wBiDsbGvqunkMa6RiKgqbVaRarllq
adRC6ikWm8wUBzValwfesmL+YnZ7uQnDbxzqlFIPBgwmLNuFhe/BxkarhlGsSj//8exrcEFPM60Z
dtKSLTQq24gXEanTvEs2bJn0FALzJuST5gfiZEwfWTzd/3++XIHGUHZ4D2n9inIt2kq3/HjOM99I
zG1BhoKv5qEMg2tB+nwnvpABNkfNcYM2T50akOvOYZ6mLd9eUcq6XXxVOZ7RPuXvCQ2zXrAbfMJk
iwb+RXVvuoAgWETRn+W66ituBlMGcislTwSx58fjiQ+8qLqFmK1gkWx8KLvfa5/DhlizpZ/VmmP1
RmniUDz7Ad4Gx9lgP0rsDX7YmTuUxP3pdLQd7V7oeVR65HYTCr5kVPrWYINA31h9UTgo1Gt0UZET
qQY1gGIZAizDRb2EIwaT2DozgsNaF137rq9dntN2UcTAT3voEJs1WKAkiiMSduTzFAs7UP+ESmwk
jt9Bd4xleNrhpufgzhANvXPwon1yU9UX4mcquB+Egnx+fQC1q9lkHalfUuoEchVyHJsKIO+Ogplj
PXKhxwb9CpLodTDrDqX5s6kA7CKnUnaSEUoZ8P1HtqOBC0AcDxdqYUtt84o3xCwfTYqDbWiIIziC
5cIdX59OIAGi+4DAsUvOfodYXgQn6LV62E6kinCiP3jeo29jFKvpYPIVRJU4lRzeMm8ltJp/L5dM
2UTvYiEPjzdtxKf5qU7W9U5FsjF3TL2wTdx/pGH7MVMDaPfo15RHhQgMLn41RDF0Zi3JIkjeiYNw
+0/fJkCQ2ZeMMNF8uCFU7smP57fTcq4Ae3vQMUsg8V15aUMKpgKK/W4DR4K2aV+84WQE4MiNs6wM
8SK86l6RevfzhzjAwzVpojX9AmKHkWcwTyc1cnHv0asD036zGo7PBnLKhonWFZwTwA3iBl23h31k
9Ho71XaK7K9Gk/Am4LH7MWwXI+6/8hwwuPy8tCsXDTyC2Pi/WqJr4++fs7AfBNTFmpVDTMDZisYj
iCig2viDJMXh3eONIbZ0ZZcvNhKv61CY9VAX3SLf29xAmWXdl27jQiBQpLEZWo7MaEiVdVWpj3W+
5+vzqb+BeETO0tqj6SHH201ChkYguP7MdifOKYdqLCqq2apXCZcvSz/N44o5S/IMExpN1xcsqaqG
UqK2vJVgExRTqC3WCaiux2jorT6Cr2ULgvYvVoOOWvG++jf2uB1Z/hcppgW2NzFLdQQ2Uie0lrfj
TfaZq2qBktAF5F2OE/YhgUXQB0dRrLXJlCeNCBJbKiujlOq5C/xSOsrwoMoNexSEhyLm7I+tc02A
wdCkMnpipr2Z0ghS7gdcGUESd4w9nOonxosGLXWww9RIqxFvrIFWnOD2osdCJ/y680tf8xeMZAVZ
r2zgKINOXCCl97MrawhkherFhnGxPJl8RpVsaM4y5nzo009tqXpZwg6akG4++Z689Y1NctDk8eqF
L5QnEcFzanbiDNQHG1tUKMeKBHOIn8RKztg+CjnJN2pz5XgXx2WmeYm38DHCcJoszlMK6q6ziP1a
nzMPsUnbmS38js7x7CsBgKYwMV1wj+6zSIexi46jiiItnDo1/FZNtTmkOJ9dQPEBy8QAw+Lk+P1i
pyje/g+K7LYcvQjDpxHJNpqgIXCljJ6NjQjyH2eHI6BhMDBRJiTFcijshe7x9SawR/ENVQCLOU+R
g6EfdbZUnp/HVzIGiQ4HG6CT+Q97pgvsn+28TrB0apW0ypl36hEGiiRzyKd31p2Pur3unLA/Je/5
ud3WI9hoYyYF7aPCFvcjnNlswCAFQJgUfrKQrrVrq6PnL4ewvX4dYb3wBQ+7ki1ku8ciApskhDqd
srwdCj5OAtsyyta6doAukeD3asztuDzKdriIXkyHXuQBgnDBSCJCst1D8LfDvKeZHwv2pm96pI95
c8ymtjbWf3NDzB+2WhERqzLutMCMH03qXTjYtyAmRkoqSLYfNWsqRi5zKhSujw1LHOWtFCdFhuhB
BqpEK6YhQz2gdYFt31tMG5YGR2D1fyWMBjSemG39dbBWs6Odb0G2KjjRyb3JVlRLYcR2f6ipRBCy
h57cygbMVWAeq8DpYQOYIk9rWXt9q0D1hR1s+uj6A0xewDrizKaUndtRWLpXxjQUaxPiL352nVE2
1AmpyL6cdy2ffipjktBMRTnxrYoJHoErQG5H3MCKyJUBsU1w/MJ/5poOW0bwf0Y+dnBcszFVwD/2
kS2KH2mwKcFTwwNL94bUosBviN7WjWBBk/CZobDcTX7OuoYgF3rw7hXGB6V3utyXmK06Bz/KkT/K
ZVo9z4Kwkzgnp8+C936/GKUYVKjyCVnLest961hTm53cgB6ecTi9uAZ89xDHyEpbQ8eZEEhg3Oyh
fGL8o0aJuujm7Fm/0gwc0zzkyJ2DB1gE2tk1tqyliHSGONJATtR7DUQfRpW3QK1bUfBpUQ2MAMGP
DOYOvmmLmYYJ6ZXVLVhH8xIhuygC3DGEvO7cnMG727rIszH2JB8yUNf/YKJ9+3pYoYprVYZ/zofh
3mteNzWLUEqos5EUHZmDrPsYmqc00znyGu5FYUZ7/mpZDB7xQj2cBJwAuzc/tf3H2kBLk85zlsF0
+F4Xow6EWfiqyS7aA0NjG3r3u3xiOjzSXUYb8XPqS3t6WHbyu7cKqt40eoGxCNgJZIxGzq7EgRCL
ILkwXtIYr8sx9f402XDJGNIG1TWXtxuGlTwA7EHv/mrRqecvneGLol065xz/69boaDJvj2CMa1ib
POp8dxoJQpR33SQttQ5853ixyj+iBIi06HyqrAoBET/vjajsiqjjdpWSSuDvXQlk8JLHYL37V5gV
ZGwVA/V0bkGLdYwLBZl6r4GbXXEUaHZphwSrGqXUh5MP46bTpudJDmlqbSUUTiy8O6uVaEnLseXZ
aawFJYUL01TPTf1klc7Oe6I+4M0X7qpmygrF2RJkaUZwsWzAZnYXE80R5x47nis4h/tDrBNoItHT
UE+7r1SVMVFmlYaV4RiHRQVwPu3XSXHwnjE9TwqwbiOAGWyrCdDdqvip8Uwef7P6g+vxzA4cPomQ
wKt1IoNkx6f6eD2d6u+wnRCvdHB69fnUu6Wp/ozCTZTF4sjCTXG4vSI76UDyow6Kn9UsvMop9LHt
uCg3/k7BC6/fwQnjJA/ob82svc693wdUFB0q/dyXsPvB6uIXGIyz1pDuTMrszeAQdqLsoxKzLuZH
AkO5bQoDthl+sLhumjfhuVj2vAmaKFx5EVHDoi3XcdeWtHW7Tbub9ftwCRr8v8xgpquNbwC/GHmr
VZSURaUwl6c8nkBOpArflh1QUgHpdZXWp7hyOEqnTig4cuY1B094sW7Z9bsvhNzOlZ77QQuouoQK
wxsVMdNhpjP6nFp6L7lQhIGxFHMTrHxf6fMG8VpnZgqgy5li615yJKToep+MjULvcTAktlXkBwmH
ONCX4GqAFsjfJQiCI8fv9kgNV8cHqBsdQtJvbb5snKOWUTAXiVcy1rQlml1KpVq27TgrCE8tdIoN
T3vK+ZI+l7F6Xb21F0KEVtof6l+FA/N2uemgL3Qp4gGYh76g+A3jDHEUTtZAiXD1EJ+x05zRJB35
i7PKdU04+eQ4opY+hnpXmtm2x5DzB989dR9yavuHQ1kUYa++U0h44KDB/JnyC2cR0VDHz2iNwPxH
ZNhywJBhh15ls4t6n2IiHL5ny2bH3bOri0tEtEfuvt2B6z4/iP85VMlNi+nkasIH2RC2/k3ve/W/
wLJM3m9taomUJ/gSbiD4YU0kVijAzxt92Qa7Xism4dyzBgBgWwGVJHHFcO4bEEidOE91TG2ZnG2q
2jWidf1Tp//w66hVBze2WpR00C1Ch/iS/NZ920aYXAQsCTogZYuw+aPqGPwQxVW6DbVOU1cRf4bh
32qspgKW70QjTvL+4jvZIYja0ybwN26fzNOtbyc1blvaFKveZQzbFf3nvhX2P4AaBh/5LObsN+hB
uVYO2/4/Ie+rqQbMUv5OpltKfMlhE7AiCIBtjIQ6Hcn2yQLgUiZeVHj+VdEL1lPVTtF0Rl2TKI6F
UIfA3r+Wf3S5bqXAp6wIMSWzUdNYzPx7bzGcdV1hBFgS9oEXjfbPlifJfh3r+tKIfGkI8tKbsVu9
j9tfHyBmAou3Bi3h47fMI1XVMDe361OblQOrPXHs+xnqZxPY/m/80DSLTTlkAedoWksx0qHabkw9
2LIhLxXNxuSqInz+YomnRc4gGkEXuGPaIWuCGD7XVLJmLON4SsLFCfydbmnZb9IIIviHitX2Q+dW
nn0YJYH/SQRIvelny18qh9bbN/Srdf1vcfz7/vzyBlyGbvioZqYtbdO8Cguo/BQBFiBCJWZvnRDe
VnqgqqiGe6VJBn6MBGBvOEUAg4V3GS7+NGbP2TzENFyBHZ7PMvWQ3nAduLuqt2RQ44+lrGORdYEB
1svgQTOTyIn1HZ+8R9/UIMNEOgF7K7fVrQof/lvE8dZAHeA90OXtsUm4QbAavJv4eXPP+BdIFu1C
KXOY8zd8aBky/TDs0Ly3UQvNYwGn/5hnHwRblH6LbBo6poH1Qrv9m5Jkv7lDUQgd8NVisRDP7a+H
PT3Gev5I7k4vMEgbjitP5aNrBncThwgqHUyRJTU2wXgBScMhBb7pHX/NJZSxzAl64NM5253LuJLI
MT9PFiWrSmlEp93Zt8x37NoB7Wul0u1631ZDBDhsgaPH4pbooeioSsL9FMTDimY60KtLZg0oro1w
czLWvy5sTVZz3iXk8u6bAf3vz9+N9UM/LBeiJNv9AeANlzp46oKJ1Y144AWtB5vyusgRvHWcYUKA
HrQSK7gY3wfze3TBA8jbikDQNYtZxBw838ceSdnG+PM6DQKze7I755yL7jDatf8TCzWDJ6tIFhKs
BV5hkF2oRFDkyMcaEjK0ixKz2Q4jENF5nMD8/p9IreoQvzplJcPVaXZT/AyGfz53/zAY2yvW3f+0
CTxaw6Qm9xOX/A43yUICqLwsRra6H4SHUaOptdxIh846qD70xi3rhRLyfMaKue5PeGD3MqhZuFMC
pHaRaLT09e1MHfahRX7CZmdEgPOwwgPRRv+X/N4ZlMQVkuVkRkHSt3Meex0bRT0lo4/CDTE9Iuru
MBKQZDvtC0BLPS5v0h1C1ybatWSgU4zrSrIOaDetFRXVdw7+VQfseyfaswXPC8ZVOteZ5NY0zcPM
DjAiah+CxQywO9mSv+rHcpF5c9aP4iA11QPWghBMhW+eLWZFX9tT9k2xWbtnZY38I2L+S0mAXHbh
rTRAQ5g9oK0SAVo0wK9ZzpBE+vJONP5cBrdvSBEG/P0XopJTbopd59Q3sO/kKvOjybPE4uMVXL9/
Ud/syTBxWBpc1H8qBauitisTseBYyMzaGlLTHMH9TPSymm0Cp4DLvTTtINF15sIqC0zF397nc+7m
QYyazwNT2UbWbYy0Kqe6MeqNBGky+eAdtUike5OteklC0+JxgEuZ2KNhSd5Xjgi1ivSv6yYnhdeI
2dp2Md99ipRYHr/bn68LMZhPGvEOSxwlpn49S8OFO7Y+qCXn5RrM1EQI8cep/rCN2jncD0S9IToY
NVhAJ8kIVk8cBwlnswVabXjRsm4qDohPzE/WcV/zltWSY9DFRsKOVICEI4xt2oWPs/AjpYk4WL0+
D/KxvJ0Stxpveb/mEeVTnjEA3Rg6VWxgN72r9nnr0M1PplQiELyvtPktbJ7Hm8LFIp11pcyi9Qlh
5TL9mOkGzi1qQpaZKcekV/huXBZqxJobTBAUFR7nQ6mqMbJxOwbR8FzhlqepjhyiVSc0zWQJmyDt
73c2VMjrcH7pr/hVcFny29VOsfKwOQf4oOFIden80dRUDhVQ0xHh6p3NKMi3uoZk4Sv5jEVWzbxL
O8GIFeJzD1i6Wj27Th7hkayyBr278eias19KyTsoQc+nPkWs0pRcCPAujyXHZ66Vr0+eCvwApVrN
WKOXpk+9S/TxbIlnVhYGYUfqq/ToOXQiUO2KB1DYTMEDx0G+UPLzSg6Zsu4JCZ3nZmSLKDXh54Al
zZO1YIaBY5ZP/xh91Bugh1xjsiMdEWAMyhWyXgqn7tXbb5yVC5n0qFw5K9QPNw2lP/cFZlpeEB+G
4Ff63t+FHk8lCLzwoMJABD/9YYrY8qMRaZcekzBt/RGhvecvMrOsrr0twDY4KBBKV+EbIlpvZAsj
p0nzsraIbO4EW6D/lh4lYS5FmsSYDmYupHpkeW/yW4nmrtuuIyyJPO98uCc+tBkZkWVMfoMSNdL5
+GDevDti98AA4vIfXFqTmQhWP7YzDOrOqk5jWQNNV8oz2hKFCPkQS3MrJn+j+wYg+FE99x4GOth8
HapNCvObdzaK8LqzAGfYwSrhf24LzaS3jVYFzo3x+Oic/o6blrDqChpZtWJ64YyQ2w+agN3ZTUv/
SRo+eGj98s1Qfp7JoTAWI9IfrEOWE9ekZ1RG+KlKLUR6TbMAShvTVNcWJ1E1EIbZCwhweK0zfKEZ
5ws/kvm5MB7+MI10kJsN5J7+LnPPdEYOgy/JcfAiTxFcii/ha5mDfoOEeUmfCkDfmUAgt6/9+vV2
FK4AutPfDzXtTSfxxk2HmbWoOGV5DYCb0FhEaBuVjV7gVtvi3vlLLQxd7SWZGLdprdDQ/PKtfiLm
Ewcow8XxGFaBOCnOEPzMgt6K0Wy8SZ7Pjk4Qr/LPr9SDly2Q8R309NdYh9BVoEworP/WextFAhp+
BIBV/Y9lmXr9MndLWRRE5c21W2rXpq/sfGqOVMK4/UsPyAj+j3g+GL4KUiqoErYS+otoobQx2KL4
x9kVBk3KODqnmJ3sjb/T2kqh8rqren3m/cpRfTbgMpTlDZsPzds5Yrk2pHvPPA+v4rTXtPGQTlwn
hZ7PaXC5ZpeSSA069vlKP0B1N6xzu56FfO7fMWnscJGXZT3Fq55Uk/h6JgdygYhv0bADwG4fABlZ
Z9AC7kSzDcNfG0JWeGHo0f7gcqEsvPj9n0Uje3ZXWuBvpBOVRv+Hd9wIoUU5UKLY2xpiTX2mDgsP
LcGAcXHtg7/gb8CKBD5zUcVL/unBMeOqhsceh3Kg+jV5Sdcb7awCpsmYAIOSlkRiqf8D/RwsGJXG
oyzGo7Rw5VX/p84aCFAITDDBP8fPT2w2TspWqex38uvupM/Fuskx3fhvTdgPpBJFcSEuut48Yh4J
RekFpWEETici1NqZLdXsr3i+a8olGmaztxPcLtVTC3MuQymFd/8+1HsvjfYDO8SQWl6KdejuBqcM
aydt3QLnI7xOkaocUHxfKEs6CdY/mAqSi9nH2RZB+6ZYPq3dfgwgb1QL2eItQPAHQYH4C8FtcUtR
/wVsjmY494exr6xaGrpvReMA9MSJSCssT00oah4hinr5YGzw+T3828Fyhj+GEDfEoH3U7PBQcw6R
QvP7NhpgfpBfqZlpumIQJhCwv3M9zB940oZhZL8NcoyiabRczlA1TntZS8g1avMJ0uXRLFbi969v
Jz/XJZQY1duX9YMSkVD92lpb4QSY4wTDrrAjwVesrxh65WV0SkxwsanaGN2bjY9Y4HWyKolQ1FRu
gctEQ8pVPyellPMoTd1umQ0TF3BI8cs34mKcuYFfjkySJ6IKJ1Z7AVBLNGHpGRvA1U1egIq2NAOR
+yMTYSDaiuDUYdkYabAWMrCaUDIAM13KhiRXoV+oKVJIWpz/kPNtGUZGHvKzWJk5CpXucxS65nbT
Ls2LfpG/I+/9O0KOhj7hrRLSLufZvZ/HrZm2zWRIMQpRKzFS8+drlGoAzIWRErk49pbhWUJtZCdL
9SrL5lh0ofNswY5TD+ng8+Y750stuvWRlUPhiFh4sY1lVa7Yze+wb6ejKnv5boK2rRzhW+5cx6xQ
EPO5yztM+xb/YEFzI8/mGOsFwjpfJtdfOcZZiuYxAD6FWgGmbKa0NHWBqBp6y+hOfkDXb72rwtLb
z9qY70PXqUnxOrU0LRmbkimtAeyAs/vsmf4jFqSGMoGO1eebLFEpzFNWpihhF0zkj1GXD3B9IBPI
IWRHbQsXXI7C8OebGQUftVomjnCfogUEOoZRl2am5BSZu8xuYkz0lBtm8w9xJd/ykVKZmDmAokkD
7DmvBA0le2aWfudvldbODgmCsBYhmJofLaENc/lwxxdg2+rPTKtLVQjjmtS+YExBYMhErQBdu25C
I/6A5LsBLvsWmEPY9JHPfFFv2ce+6ad2ZySi3CE4npcUebHNWvAWhfDu5W60MPhOTLECQaM8PXgH
9yKz4dyKB9ENLkubCKyqXVrsoEpk0OLW1QE0JevCEzmeRJBuzUSctxaIoO8dA8AVNkGtdmqguYAk
+uKDHJYNnvv1KDT+lOGvZhoi15QcQri5IMFuPwqyM9EbLrWoVVdMEwqkeLC5cWtr4JmzMvQyV+yb
n72+U7HP3NumFxx1bzJPout0X+ubpedJp7U+ydeuJ9fbVDmVdx9tML95gpBoTMrUBuwzq61nAerM
GxacRTXTB22wcEuF0bmCUaZ7aw51vcZztIXXrd/Xy9jGAvMY5bCnkka7adLmH9j2EWz12fGvflvs
NrsWoGGtCxQKxtp7fF7Vjb6jpprNUdTdOW40Gvxtwj+TX+mHFlZtVMjD/uD7+/E4ri+G8JOH9Atd
pGKLMpWK5M0BjQFNmC9FptUgCc5fY7gUEYd3VTUr8vruoo4fRTt/8r9qoYEM5nNOVG9n/e2ajv08
foRLVB8PLbIkCMCoN2EVXQaviXa16Mu2LqPXcXf34hZ3fCMiwGmppEaDEWSjS9kJi0KiujnlkQIO
FRHvlpEQArYc0/D4SAgU6K4UfyNlDp+fFtqyLsR28jJVpmeQ6YWbNGcARp6LMZQT9DVD2/d7bfGd
qQBzOYS2x8UmsIA33Znh2Cf34T8B2hKFjpKzM5fsqhm17D/SMZ5gcs+SpFsnDzHHvqb+Na4j4nHS
xCL0VzT955NkadP98jPq1KgNXXHNB12AxKhTBUkmcZ5svrMCQugR/uwl8yRjnbsDC4wBKBKG7qYM
NSga3jFk20CoDD7jeq8lytYXP95M/lhWXICgQiN0l3aVl72WC6rgaYbZRN/vpFVhEL5O2BvRllV0
SeMwiXCOD4z+4r+zkAmu1hrRg4ReTYt14Kf7d+qG8wcBC1PXBRvW6SkBm0TMDJS4HcFrk3TXf0KP
kuJ3RMw6T9FY9rNfk00kFle3B7xlFJAUf4tnPiuGan6MTvorHQz7PtKqCmgWBlmn+RATV8bqYydZ
X4fF1K/v/oyozaR5yVbq5dLYDeVZE65P3AAsaiubwf/EhIlWawCf4nCQSOkyoifUw1m2MVDDview
my06P9hfjZK9wugpaTyX0w1EE99DT4QiamrFjK49Af9Pl7wTAjxnwsOEvZwjHCHLnpBG351hHi4j
oILEz3CNspcVcPS4Xi/sg66/5r3kn+HJLFBZ4vdmpn0RBdpiRqiXa7lGyApO+tAdyngYiXgsLRvf
UNqzajQDCdG/4XLlFYYkxtVXL3omBaszGvLG0Oob8uIGLMYyAJUwFcvoJWILDgbIgeyV3mfagXyX
Un7ItTuEnxrNmDYliKxcC/FHnF5CUjTFxXFsyhHLAcrq5BR5nBUK/kjzOpdusgp+zHQ1i5/2eDrG
N9uL+7SLnTtmtq1Gima72avYFDp0W/Mvztabuwqo7xFwEuvQsNXpBMMTccHZ717qawVKOMbZVjKk
MiguIDdwsME1jq20B7e6yOPJa9Ax3aFohyA3E1Z7g4Fe42ThhWOotX7fd5ce1XaUf78initXcR1i
lABzUtW/TlqAsdodRXbZQNLl3O2bdBke0cVBc+bbYgIlR4KTw1FniXYwHVGmSm9/6nXTxQ6LqKUG
DbEq2w4/R/Fp/F36NhdX7njAOfPG8PEpvXu3jcfrnPK7x9WRa2aFXMqIMs6mj7fIw+ApCPVhbtC2
FgfHXhv/WgyqWb8XecQu0HMxz0xKf5wifcrXQRtI1HNs/tPabpRHSxFuyoYJS79WP0q/ek8J3nY1
x6KYfHz0xPoNxPPu9XNc1rhrzknU5SAQA0qkYHc3Z8/rvQeKwLz3BqktTCMER07lvXpAtngYSfJc
VTpMEqZlMDTCGbtc8h5wbnAn2y2Bvl/+SbKBw7RK1fskUujBCAEHuwQAtttdbvWFW4VkvClomLRy
B1hqJXUK/xwL+5TS9GnMpNZWniuBV8F9H4Lmyn5zUyaAPU5V7ET99l4Uqeaw0L42+sM2FZ1XVLqS
HqY6Jp7Dhv72l/Nhcit5Pr49nct84gVN32C6UpRpYlN/uKRcD5NDTnrDFEBk7tc6zJtjCa/faMjy
gN2loOcNb4OAXKO27siUtl0dNEvxAJoSB4UxZgWeZ2OB0+0hiJEFyGACtbCGH5JIp0Q4/L1kouIy
40kIjcDy1q+9nwDqRjLR2RiEA/JuOcRT9kboqNggRxb+e5XVvrM784+k5peilqaml+EXTzUKlL5d
L2z5ljMiky+2q+QtP1FjGAEBhY/186nGmCeB+3zNvEToOI6ASj4elJmUtrjxFm/TJzEFgwkerYg8
RDgbdEKpLie8EmbxyLCv6mhg+WOIplIz34CxpENZaClW2fLwX/6nm99j5nrFveXQMC0w+9enuUQ2
1/3z1H4TOtUS42ZMdcfJXDxkRyMx+KLm6JVchfkvHvnR6k5CHuxtWJp157vHzgoChqs3zydFTZqE
D08YMPhiDmUXEhi1RBgbURDfQJTaQk6hcf7Gfg6HN7kH7KzTkBzvk2tAWsfxnp85MyI+lACaoirz
7GAenmthXFctmCSREcqSntVMAzA45l6VsTBKvz8ei7iHTn0uWJEFWtBSmMiXItjV8piGRU6XWzax
bfyRm0hQWmNsq+L2M3kYBSnpAJWGosBIT+nCt3qUcSVTVlGSBwsaQ0Eh2vvg/1HrOkC6tBdtnGeo
DaNeop21p77J6N/I/U232MxlcJHd1PqL6Ppx0aRmzpqqcNJOPmsxwGFElqYW4myxCurj4WNRjPvd
+RzFOVhgv6wbGEE5FAidmq2jro1MWvqAWsJ2yvd6Ja1gX2ZEGbiwJCWb+Bhj4tA3q7H14c1FN24I
V7zA/noLZlh29KfgXC+g4oCBXOGe64hFxrpENz1fEausMK4YqinVabv2BdOfvY/HKf/BrJz/P2zm
30tQKtg29Zmv6SphVyUpuja+StlEJoUvZb1DcQ1d2hKinN72D7ScfeeyRJ1IBjYms/jaAXCsuUUE
jgAIo1rORolUaGKPgPE3z/zmsvywtblp1ZYGY0qSU3kmEpUtBFIvDcBHtNvVv+YTw8OHND4atYZ4
fb/UBMFTDa5Co6Tq102LtrC8xj18Rl5AqXrvoS+8/LxK3a6DeVek6nbUgeOsA8mvpxTUSkVERjLU
s3REwRplwSWVfBHcoLnbApk6fkVBdyMiZk0BSoV6rQPXirGevvXo6w+oT7bH0YEhwI1aROx6lZMP
RxzEzcsZPIyQmGzMvM47upQ8nYYUI7EyWRCQhWy1iAshB74YqTgQIoW+OP5gqHt3bmTsnjKFxlFG
aaA+Xeh46lOD9tnFaF+0hisXJRcyBjbPqyBVWQb8tfPpOYilv8QhzNRsoyZObsDLonVrttxVVUHA
gBC1W+ZgaFz9FJXUpXtAP4cnxbCJBdHlTdwiTh8RxL5NQtaZXb6Qo5IL3fHvG8JV5C58iGKJB4eu
cK2iTQiIr2wzqverqBtt/566KlgUKCYa7WazHLBkRT47VE7hA9mtKLUelFm4LFosXoD9vfRRJYF2
izpm+hK1dz9y2rRBwjXd2RnoaxUZQyVZ3e2dQynz7fmpJegwawKvsPQx8F1TRQIDuc/oKxzz4CiD
SMnOMFN3dwywsVG9geAGeUCUHiiocnrbSZu7xSDeNe4gmkGQb2jkBxoiN6atd1WQgg2AYpzVl6zl
vuvQ5pyZayGyy4TiIN38hHRtoL1MiBIKGU7KOQuO8irj0ieqZFzmtSCyQtOD+CC5pwrrIWpNOQbr
r06X7ypBpn8honfck/oKWOjUXPfwmbpLOARNRGj0FCB4K5UOIo0M83KsAhb3ylJPEUvaO9y75p5I
Y/1HhcIozCQDYOnZKfC62f1jyd7x2P6P0mv/Gy09X3rhuIh6AW5+kua0sn9PSNL0VqNuL4lNdXnI
YBh9r/vXD/H+vL587w5TLe7hU7wNYHqdD9go9SkCgu/88/z1lS53Y/zAQLy8hUT6HTjjNcidTCG7
UO5nFX2C+cZl8HWePTpWLsrRMmVoeHGHuicutiAdP9SyKNe1Bp/ot7QoJ5ZGVv9IJ/R/eU88RhyM
iQceNxVpIslKVVU+cVEnzeAP4YQkEurtDlpAdcBPafR1Yo51dCV3cSJ4NLmfhoHEgpU78y6Vhin4
yAQmrCQihf+EOMtSbBcNke+554R9TGo+kfyln+hdMaU6NbMvqETQxUfLYmiIQ5G3tgP5iLdtZT9/
uIING5aYh/TK/iJheMIo0WxD+nrRpO9n9tqMswKyXQLmdMT+GjhqA+kSMMNRFVrmWxSGGOXzDwOp
WhTKBb/J0RfmFHwFleV5Jqx4+nISDnrETOYJ+sEIxPWX04GT0evUNVz3EdyvSpKdqwEoLyg+Xngc
REaDklN5khVXziWDvioPzXmvbXSrqKBKUjYvHMbjku90Qw9lwR1Gx+wD4+zXeOxpbRWljaeGDLeU
1apN3QHrliiL+Wl5+O/5OLIBBIZfAAJBXkiWvN+HyVkeGp2l9uQnCNDnBTA5RBECtYfcseJ4KCYi
qFR8NW8Wljbs4jqusURulxugmAuuul+BuUD6hLqtYXGJEa1i3m9TNyUK4eStACX0LBFJh5emX5f6
Lkva+mWeDHbuJNrd9P6xlLHVAwHbG+T5GS7gtHQkNNT51ukuvLd/Tmsng6pfsIJJJCEuLkqF0330
v/Nri2Lvqv3cYvBKVJTouMSSCgm3McZhTmObVqNq05GxptDq2IEpjPrt3Th5RaPzNIfw1B6EHdmY
aHoor77mbkVz6sWcbpIoyxYhX8tDNm/HKitQ1fht6i7bd9ayCK1ly799OVpjv6fI6vtqOaJPH3Pb
uF2LoNUQjh0AsBEONG8zVMmxG9ang1o5I6soyhWkwO2sW09pnwZhR3NQKa9Zg1GL7w4ywgGHTnPC
mKqmdb8Cr3j9GHKuXOKX8K5N5ZisZ2a947fuhwejrnOmRCu6SGu4yb99rKU5j8UVQIVYck2t7A0s
gLWdhOTLC0ESi9SqXntBOg04131f8CnL54D6HrTjat0Ev2jTLpZV6jRyImarLfFpvnXu2U156r/O
vpd7pleQiWdI/GW/34+rCOeccUXMiWA4IaAeYW1AtWv/G2q///beeyxg1PNAOFACrob2KKuQRYfX
VdgIN2qc6I2qzVKgTgS7IRjOJQCyyv7+9ZtQj8SqsKcqwYdTPPO9j0MIdlmk3jhlUwG/EpxM6OGS
X3Zgiqi+JcYxYAkI1CNyPreMrK0sPPcW6zj1LByKDYS7ukSEt5aAM1rgj7XEkL6hcXmE1zF9WrMY
eBzxSMoZ7GbFQSCcS2P/QabB+r3Yiwzb17RjejjA+opzkuqeWkg2RqfswrvnH1LdFfCJmoDd3gLx
Cy9WwwvBbemX39701S0gS2gdS9dqKdI/POQ6+OEDNXxxkucXQPHpaUNRIX6pjvX5G986i5DPfP0I
oPctRkC5weoKHaAIL3fTkphkiIKFplrWNud1hXmR/HBLWXz9loBdY3bggXYWjpDCqrnoVcyOTJTw
db0757xyoZxkUp3usLn4X8Z1v5b/quhqjrhM++nbJjpI0gFO7cKtE/jFvVqEIb77HA9qLPMrjRd9
zNU7d2r+oV4a5nUtI/8xF2Wb+pkBVIuIb5FBrnKgF9yBMSReHX/lKaaZFBVrluZLBGgWhrbZW7GU
5pE33qhyKXjORsedty+QZAhQ855ggih8IdIeGDdeAjJFmqver1INPKeJ9Gs3ymH5wam2Qy9Zsauo
Fu/Yi426v3uXbkmzZKQZg+hJMu1Sv3uw57LeVpIrlNa+BZZWNt+xubko7xk62qsNJrKcgiybmMz8
dq6WkV7fXe/M87wbHIcnaFi/dOjl5nZRnAPz6qiNqOUVCqW2TlLdbpxpbRhXkZKaWZvdkK9SSiBv
3vm/yH0MfGnIy+aKbVkadiihXMG0tLTAiiU2PLWr8ozQdngxuoZ+VC+Y6apua3CuVjD9pQXsHznd
6E/90eHKCR1EITep0oopQZ2UupABhNzHTRX+7vpoAK7ME6TmIvWPxhydifYTftRqlvkEaoo0hdWv
sYvDEvSBGCXd9aGx8yN1afMg0u3gVxRFQkPbfBRNdgaO+hPDMzAIWuaefOBXBdTWE6P81Pes9sYd
MmltQm58hsqojEZGtzVRXAcC+/hUOaTQGmYtmzHD9sSAJvRqaeiajqvCQACpJ+/XHlR4LTf5mVUx
DPLQLniTxmJSZe3aO3ONWP0ILwMD1NKmcT48p5XI7nySxp3S22Ko3+deVntIesT0AH7h5/ztXfbw
rh3lqlEJebtmF8SJrJc/5EjzfqWOgKFR6KbkAtYc1YihHE+Zq0HyQ8+LLB+yEYuYMF2bsUowrRWs
9FD8eC5GpFXPnjkuEfRoC7wEmuXeKE4zjE+OA/wp7I4LbpTbgHKBt0R7RRWKb7NyMRSVHHWC7KPS
kTCGDJz62h+kG5koMEKpb0u1db1jqwDtSbo/+4O+9lSUVQ53B4ZUqM9ImgZtopDIVW33uN5dcChx
ORhA5ws0opkUcrKFCj90RwKjqLmA6hehVEm7nvBpxtFH64AVFO1ob7rNuTo7XV9mrcyYixfkIOR6
9aIAFKeVBeN+lhoH2Cj23m2leCfO/pRQREm2rncBKeZkFJk5xhAqf/b2IspE6zwbiqTu0HoYI1+G
+nPTlGGp6dFhVuSFiYZx2JewgAIEsUN+5uNIG6Vesr+Ob8f9vD2zKO1slisg9th4QJfFtyPkPWzV
lGv1p7sNKUM9OSIGdTyVTJhW7KQTufyHmF+c73rxQ5xAVCTAjDq2E4JdvcX6VHbwZ1LwXI8DMA0f
qEbbKA4J/0jkffXz2E0ElqTnYHEk4IDf6slNL/MRzXZUsmWFgb3DtJu4Bw5fJx+ah1S3YpgOu7wL
CoW3YKw3/J6gpqyrwUcibYamA/M2H2RGqVuSboiektv6ezBqDxfNt35vxARPVrwurs+z3bZr5Dv8
odqu9Zz72vGyQLiF5+IrC08VLCGFImWwQepVpBc21LMoobJiACkXO0p5hkBeaYu7D7EC/PCwoI0S
Swl9NKIJ8q0NGKwQGw6IwziBxSDZOoTd6ZA7QIhjGgjeUHT141TWJ5yo/I82oKqXZ972Jc8T8h/5
w/1YarzLi4A2TCV74eqK15nGdaEFdfqlxo7tWQOlhmJgQqbaNfcdG4PsaspLAJC8WZJPkr3zvwiY
5NUuHItI4EfGfPQnognePMSdYqoN36tsz2+L2djFvV4h3wr7tsFdbMcv/aW/J84XlRtXF0jR6zDy
g1GEXOCHFYO/b9uLG4rp+eWGdZ4nWfKD6CAwFac70smjd8Uu3hSgRZkKNjIKfaj8z0Fn/FNtV98S
99hX4g+Hg7B3AJ59rovHSx9E9fDRGoEd2XAJXO7I/H5UUBZVNA64lUkLm6R9wxAMLuhvHmwII/jR
9texDl93zO2+SEOiUaZQyLJsF4b5dyWkVpAAfRAIrkPcENjPrzHszFrzbD5w4XszMXTu4JkfcmLg
GTWjVSDhyeo0wns8UKtC2gWXlp9Y7OjcBLKdOMPTBMhsdL3BSdMm/juJi8VXiFY0OZnAb+kPNMZn
MyD2MCPgrZ0T4Q6TmS5YI0EMUGI71wuAs8a8EDvzuBP/3NRb4F8EEdGKBne2rVs+rcwEQeTEjmrN
8tuRu4VPaCxmeYoware0GM0KNzOkllxTQdVDPevUHA7UiA2ypatDmXDf00GViH0nImGylxrgieYB
GNZzGakY1eenr/W1WkmFP4Kqe5Qr+rH9MkJuLnJajrld+88YiW8cCa1mlLpmSOwdJx16+k1mHuOm
s9zkb37f8cEzYjqv5oaF9WCGJ98kIWS1JSCFioDbqlvDQiPD4YUIpg883NezTa+lnwSl3BRFJxGS
oBZ3FKin+KmmoZeSmap24UMIkcRHE7TQPEBgLVTvPzTQM7zPfHY90gNNUJ24DhrG9xMvFVKypSO2
V462SMcjZ5CQ696BfVelO9hGyVpLvg5t7nndT6vqUTzNwZAWet00fR36qoSh9ZX90V/NYAktEPJK
8knE4Fzpyf5NKlU489IMZ4CDqvqkX++FtKdtodIXCXgj5aQKoPzA9nXGyCGSQ/DbGC/HB7NK4Et5
KWGMjf/XeTDHdxQzjqFk40+A865Os3/7jEH2I2UWkN0BpV0s/hKHWH6ePwVVgtCYW78QyZDZWM+2
WC9QPcXbKTEZmSTqzIWjxljptUOa7Yn/jrR6HthfepAVS2poAgKaHpkt8cNkUrFGCpATEgVJisQD
T1a8zf7XJ0jZjev+zpBtg0YrNEKAlVTgYAW4hVZg/DD/dZDWUR/rgPBwnTBlpLDKZGcfQ6IW4gjm
F59CSxKDkbGOnQbNhwfOhcI/XGScOnEG10ZCcY7V94V0f/FcMqqO1teJvdj+VehcrgkJd7bawD6V
pZc8m2oCtG63f8d76UV/9LNnKVScRZIx1IPqb2q5Qs3CG5oaWGQZfqBJuKjlFcNyl2/jFTz4Rxiv
lEaXmNuKBM7+8dVJiS0vpNGk91X2a4K2kAcwO3gIlipI+mO5Q5OZgUVLc1Cp3NWV9bJWtyGN3Vpm
BSjXY5+TiuazQaIMw8YR0CS04qHbXWHcZpWjhQiOJ9W4SUl/NH0OMGO/ProtRwJn3d2KihLwPDyl
ZHGlBSwDtabWzgjb0GcWWz/NBNHPorHMifUaH8xOcfATdnaF9Q2tDaILWLPdYB16rvRnRA87phRo
4gqiY8pv9lAWsr7LqsoFQQdSrO+FiqlKtPS1AaTTd6Si+Mvqqbv5VEjo3jbGUeGH3Z42T3oNaZVs
4SOwSa94VvPTGN2738ZvpAApBJK1lh3hp8eUJkqHz4iTwPFJ/dZ6JCiV3htfJlQPNeXz6pdw1pIN
dTyrTQyHP6EAZ5MPXJ1WGMvLzCd9SHrd+TeRCtQdhSJ/7FEb20Qeyn9jjUC7X8v00uByAaAbuYzr
NNcTCYn9mYgueB9amyK91E7yn3qdj1TEgXlAZe+1UySY2PJqCF0ZrvVcCYD3/QCFuEj/SVRsehNu
0/rft7nsBOLcudz9V1fLgMPnOXDJhoUBK+HqKHSMG+kbe7HDTvdC+Z3iApCstWVh7hABoLj+3gLj
YmFpW1jgQpqqou6b7kRKyRpAVJrMXReobn2OXpOB0hBmHqG7reQenyz89hPq+SA4FP91REtYbZwW
Y2yRnxfP7RbmVn4K46uJNSn7eMCEZSqs/4pgC8dQqSIgi1U4rZIh4yPSqeM6IQfpXn6vl9f1M98z
aeXVkb4cSR1ZzkPgQlRbexSHg3HlG3IyYA6OonYK6HJGH43+z8Xf74zkWWgTbPe2r1LFTN/fQ/KJ
Ejt+JfKjtNLSG/QPSrjkpJUcSQ5RCKifSOnYGdP1Ij26ntEIxuE+uUnzanVVmM0+iQRlbjRJr+xA
DSMoFVXeBGj4piUNQnaaOAc+PGDVpq5TovXT96BO4qdNbe4ir/JfyPiZbFafgU68QY+AcLb2Ds/S
4r5zxkbeB+ZekniDJ2RZPgF/KLMBQ+Lr4IPZjKq0N9M/iLoFTyurhodnC+0NJG55aIlPlPUkIpSl
ANJbJFce8P3tnIPwdXaqyxzd7MRLrJlZNh6X1eRvaFfn5S1kOcSwzb0gPtR3fmsFu1SrY4CyKi/Q
KILW/PLRYduJqEGLkbxKmdlNIbua3F8XhUWueDrYteLUzRc/CsLjidpxOW4lc9eTubrOg9BEbCjY
3lWWSIbCkz64mhsG3wc/0X+Pb7MSrM15F0ZAOMKrXGiEnuP/EGXO2MFCy7qzvqSWUi4Wg3xh+vQN
FrFi+Q9OcceK7p5aBzvos5sH+TqSmGRP4Fk6d3pdLFTkFB83Di814YBB2qUdKHviKzQHmXZ2iKDb
YKS9j4J4M+sQOagmfz1i2JT/7t/54sYsQYlAYsZHjGAT1PGK6sLqpHz5f0rCJUgvFMIMon5uJU8k
oc0Pn7EGY/2Jel1pv4t5Sj5TIwr+t3fMR1UBnBG6t+VLQD19pVRSGgTgm1ni3j9oL4UdOZvWKpfG
XrVO0LbEh3uSYYs6abWidWqvTbitt+K5AM+kOnRcas4ZM47C7kA8xSLfxYF1WRXXdofYZfsS3eVT
MwGr7Vz4IiKreXDM61RvqdMv8q3pV7NL96gzrnffmtsoFqXSICjlyHlVi9a8B5WfhAvJo2U5db5Q
oZGNah5CRW7oNaExl1sNGUzX5jjAZc9K3gRzWhvvntnKUQQ4DUdf+j/gANwJJS8vCm7vZQ/cGmPU
IsgGZWGOOgh2pddSFVmnRrYEF8qliiMZJbv7RUaObcEPokbKlSoMDnWA7vPDRobnPO05ds3DkHUr
eLbOQNicXKGtK4lOVeqqKWccdt7rUQUh1IuFY4OJmirFFPszT8ucuwDToE7073fyPFCWT8ATyNbl
hAu3AK54Fv1lV1MWakqpiTKX0ysi7AIzLFrMUDUdHxZrQv/xN3Ca5cKAEpJlQ4kG7Lxqw+VFOnuO
0jB8x3TtpXbBh1wR2lBovFdSUPlY7BHm0dH9GnDY85ImRe2I+1rffnpI+JJgfNk1dXpt1brZ6UYy
GzawNbYg+AHEX8fVOOhgtH+qRB8axpUphDmjQ3BnX6L8X793RnbPIji4AzToVZz4fcjZtCmiVqbh
JSny8AMPl+V+NNnq/Duj08gRXuih3QlluXn2gE0RHLY8NfeOvfNkykR6/bNifT/vABaybqDL5Dll
XSqSdSrLWVHiWJPaBC1b3ps3nZM9omEVq1xJUe6BrafT0Ogean3QuYIPVEaxBGokPdDJTEjx9kCT
12UetQJ7onxbhHDavTEU2OfOhF3EK52bterAxH+XLEfalYSBZjAmTIbvmMyFX1/WUKzR0Pxu7S+A
vTtcohH7MhiNfxAycac8Ucxc+q1Ztq4By9QkpMmfykabys+LTf0uexiZClUzO8l6/iANlECCx+M8
1v5bEyBoV58u/vCZgawrqz5qUSFjK+BQBY0qHOhOK6uCGM57K3Ob3TARjY/A7gwnN2eJg542Nx0N
cBKpNSqHKgJ5BP8Z6xiSidKj65psDAYmuuwprIHb1Z5e8vgy6Mw+sV3rx4GJosXRmX9y2i7u46Ai
jdNWtb9fPsFXFiGb6MFhNX5dXFWMqrL/Gx6BfMjc4x0+81ydv1pxSz4R9veWLbL0DpZAt1Eb7e1k
Mn405RosztL2XEa6MeXXMx5ZhJbZRGnvHo1YiIvKhWEO/6iHSWq4dQD47AlmTjgHA4GDFGeVv2nt
MyUODp+oD/Fo47Dw2CDLbdBm3JQbVWu87/i37J0FRbIJwUFw+HI2Apy40JSzbQjrDOa0Ztmc3p27
VcboNk9rTAngfCeibDZaIPFwIHsfFZoJ3zdkPExIy7Z8x5Fo2k2gekoetPpEL5qzTGo/n6LkviQ8
VkpieIcdOC+S0ivjGKYnlJ3j/1YQqxLeeEuoB2YprDy7qDty7fB4i5E4DAqK9/sHUyCSpv2sv4Sr
jwCQCOn+lHOLQhYSWBkqLtB1t9y/nSjXav7YioEvtm69Ibzt1rM5bx9uyn84l9PMGuKl2sg9l5At
PuJHkb3TMo67RTqOqSPMj03LKTHCCeBAiSflaogKYyPF82X2CjtWMG64v3P1VzbQ1mjwq3gI1j+R
vr1A72AlCCSkrvX1+C1MFjIf9+3DjAJ7aFkNXC077na4IIV3cUMo6fiSor/Zj2d/4PFn0rzhYEjc
RAMtgTrrOBgWLFE24DrUgBXHjgiEpbL6uk2MCmX6BdlZfzBZaW6j7U77Yb+TSO9O44VO4pjMCL1e
W4eRGkj8f14O6QJelPgoQu9d5c0UzkOt7LiqqCECse3M9M5lriOr3ohhBouepZ4QKtmzlEGPK7Bg
rUbfkRLBOoA3hCe5kkGYqIPl2g8F02vcay0QWoKuMPPvxIEbVIBD4rCgBd4N4b+RzlT+B1lobq+f
t4MwNYCJHqzyp2DHL6N2rD/xYPOr7nWzsFfCT35hc/hvgHT45VY41KbF7THfWnK4RkEVzCPXcVo3
biVpE3U0zemBXPs8kcN7yTT3gteZVCI4zSKXv8KQnUXvlb+iXdtRxvD9N6mP8z68iq6pM1hOONDb
dgfeJVttvbSxCvJYwND47qBM95shfhhseCcKBTzbUryJEpEXdnIWPyAL+n3j+hIDBBBNAN+lJHSN
u2Fh7r5SiAC97cUrAMp/itt5SNB6jxHozdDbnQZHOpe/7QWXQG8bmv422+AiZ+qnw5midZ5zclcs
TqJpjzF3BYJ9cbbPXM3D4A9jzcQPLXEKHH9IdsAO2O2rKe1lUujFTIxaQYB/T7lrE2dx+Uogoxp7
pjAR5ovYmnMeofyncd16Or2ufxSqHTLtWIwqOcwpPlZmhimh+iGYjO44bEdTQ95TXztY3WCI4Kai
xKInQiFQEqAYWtJuURO6HrzYxud6bBWLZYSQUJlV19If0iTU8CWfYoSHvwuQdOftuFjgymJSm61T
D9FprjdRymXQruIzSj6EgWfdtXnp3Azvs4wAlojfsXBDF8wM3oWfrP6VQ8kfoaI7UVNuGv/KMjtf
P0nf445XO59ju9a928WgwhXFtfyMIaVKO6awFcj3owirthi+9wxtGOBb5TRbE4pzY5YQHXqBVh5u
st6Z8E+k2bEDIN91BfswTqf8FvoOQZCInN+YOzl4amOhXwzRVlC0AOlye7nXzFHVU0//PXgJluP4
EkSIrR+dC4FlJb7JHtnnnofVlwTTs+LybZWHNMSEB6PRXrAejXowLU5WaYEuFTEysWjX2Gdlchm0
iBW83bo1HaJfiruyK/WbusiihXba1X/SKkePfsbn/Bk/FtffsDE5EeVZCihzQKUIdLzTj0wpO+Bf
+Y0SqHyWieFiJGee4wgm00UjsVqE4ldC1rZPthS3gqTRifkFxcY0NGkoKEiwaGX1HtNoF156cNv5
IDxKvlDeN2Us+gQCystYj9ApmF8Nb3nCJt4S85x4no9tR7A6JgH6Smkx4PWU9m4dlW0JjwLf9GZc
CvKvey2pXB1pTGpKJN1UMCK7pzEM9tcl9tIcsjr8i+kyjAbbMu8lPWAdhAkwn1VNs4ahoYFJ9+7+
jFllw3dHAJtLNY0bRpnEakBNDMoVz6Eb2BISXh1fvUBi8dogRCcPhF4GAFWAnw8frWPyqzOlHESE
PXl2Yc/QzCUNU5Gs1VkM1syGWuCG7tKSlatrAtNQMbluTy5ZYu6yYcCv3yTqspTogjfcVpMpWIv0
qNPwhMkUkYAxU3XvTjOBQIO+LDJnasxMtqePCcXm1V7ovQYFTb5nWvjujPnzB4dn/+ze9Nv2g/PG
E8zJKerOR8FuLkJ0hv/gzWBoIco/fxoBfX2FrStXT5A5CTo4ZSgW0rTb5NCSqZx4ZwNWBUnxJDmm
734K03RUYnANcuitjyvBl6VdqvU4p/c8N1Yq0RQF8H6vWT+PBpIZcC3Yab9w5ZZEzTZnmohJz/Wm
K+nKigsBg45S27Fwox+hfPBpmePxMaPh62Xx2UzZcMdyIHmg6L1By+li
`protect end_protected
