`timescale 1ns / 1ps

module Kyber512_DEC_KEM_tb;

reg  clk = 0;           
reg  rst_n=1;
reg  enable=0;
reg [5888-1 : 0] i_Ct = 0;
reg [13056-1 : 0] i_SK=0;
wire Cal_flag;
wire Verify_fail;
wire Decryption_Done;
wire [256 -1 : 0]  o_SharedSecret;
wire  [2:0] cstate_flag;

Kyber512_DEC_KEM T0(
clk,
rst_n,
enable,
i_Ct,
i_SK,
Cal_flag,
Verify_fail,
Decryption_Done,
o_SharedSecret,
cstate_flag
);

always #5 clk= ~clk;
 
initial begin
#10 rst_n = 0;
#20 rst_n = 1;
#16 
    i_Ct = 5888'h53a6c349b0fc6bf598fa0cd1b39bcb852bee024e8b627c073fe8f1bba960ae881bceb38fb50de3dc7a297b36bb8ca3e4c3540f77bb1da0c4a1aec0d1ea36da754cf5f20071eae75f309b40539ef84ddaaa89f637b315950b543897ee23458af0b39d48e060f0c900ce9d70c67be7e4ce6b67e1e7c3d8efc2a707e430735127b14f34c1f48063a71f4adb0c1a90026dae4a1deb0b4b4230d3f5b6524c67d32d2d85ce2d76686c6455dca375410a9ef4c9a56a87cf73fd1eecc74cb48b1e30498d2f94eba053d6016816986bd4df6f3d118f4e6fb3df39cf484697ceb22db56fdbfa389a4fe2ad14fe504bd36b09ae2da2b92f6171eec0b0c8877516442867eed8c49517b71387968a4fbec672a5d7faeef5e9c1d7145ccbe9ca0677e7fedfec8489d99f371d63731e52e6409ab7abe01aa8874313897668198db9caeada0cc65589682fbdf905b5aa3db57636f74c3afbfca20dfa9a4d55213e4e0b3f7236e3130735d3e8beec0d676c9145999e91c7b36387b83daa652b370b4a9f3da3a35e047511c3b9b8470b5d98d0f51ab3d260c8f4a8145e7487fc849bced69bf23595a9773b9da405584c86d14e56273dd9e1361310ddff7e05337961b2925d160037c8800b2539a7ab2a1e70d8419fd194951cd3c5dbc7c8b22aec7ee183f55151472ddf974e717678dab58d56e671aec533fc52d283f5936c933aa8299cb559d419b3a45fd3d88306b91d6cbf3cd625705f4602b341dcc2d005d62f32013da789dafae8ca800571cd7105e23e30e1dd95173c81f2acfd1dd4c5f84c037aaf6f219086cde9a1fd0c1885edde022fa35e0ddef4819105ebe0b9775aa210006d87e32f4025e238ddea692556b80f3717fc7a086a1d3f8566cb61b794e2d1b9323a135a58e713d408e27ed2725ed019da4a2b9552d183400f0af0f2b08f03d32e7fd5200356a0635cccc6a6d2a6302c3072c664a1bed039d5b3b9211302225da1c93ad06261bde3397ae9e3b996f2400a1ac4e0d280883880f9d55a76f37ac038cfd6341c;
    i_SK = 13056'h462396f6b21ff625b96b4b1f5c3a38b3c80708f33bcc1784bedb48bee0253b426cfb95618712ce9825a53b5cc87c8143afc46b40627b4c4bbd2e382cec457e48a7130c8412c2605c475915bf08476de4b8aa70298ab99def9386c1f11253c398c6d0adf9d97e2264a026e40211b59a26a23f16102a220a6f2bf27a14015f6f3261e274758cccb757a406005317a050c22d399f994974aa7313edfbba4608371613985481b0aec89edd6002754b18e275b97af8b4adc682b573b9a568732423b20df418da0a0f6908663be9833eda1269127702e97db82bb11de22cc0765e26cab60d256cbb27221315c2c1d75f56e6aa4c08cc8345a16b6800e330756cec0267c02d1de1ca3ca8738156c88ed6ae90f8429b5aad8c5a53fe2687d2074fdb18b1241a489e8550abaa7b559acc6ab4b5396c821b854305caa66a478039cc2cf7365f56a344d1f09aa73a667a15ce71b210d9b930403a38a2a10cdef39b9e8960ad463313b7ab3d723a715c1d729b79b46b7bcedb31b92b77864ac9146c15a89bafe1601fcc8328e657a6ebbabef8115986dc87f17234baa3885e33a185688b915883ec4809c5c9691b95a08179a48577c1724aa1bcf664d5ea49c69a727cda3e31e71e67257e65e847df5947abe2967573ac2d6159f96699ae16a55f654e8fe00bea6791135aa045d851d0d73cd159be5c00041b1033af18500cc62b8dc636bed70e4dd4981e378820eb73a7d3bc69a42dcb9103ec8bb8020763ba76b48211806529553da6487539894722443672bc7ec31646158ca66343e2e69bd638cc4a3c711e3775ce88b4968a2cdbb772a0d9af6aa39168550074a6582da19366f61be174034472182d900c0598369a6c656d30c99557aaf6e43023f417bc4a2d8e2944c4e6010152bf28eb2119a90467aa185706396f933722f19373d3431b017b794a19b98b3990188bcc7142cd23a75a28a95d2c25aaf7c2dfd8ba06e47066940c1fa55655dab9beb686428c72e90070f81a6bfb6345766151ffc059ea64255fb24aa3e47cfc01300f43911ae393e6d7a89e1c228f3b55d70b9d9d4b5cc00671ad0b69f173be9dc32739492abe003294559268c5bdc3a6b9842b0a248131d9f12cc45876eff53969865c71c20a9ef652b13b126df81d79093862c9ce0e219f70a31a98779cd9ac39f1c672b6b924e50897a69cba4d88c117520b7bc388362c989bfa861f847220cacfee508c3056910b0118bf50523c894101d78a771b0a90d7419c382f35c8206f24b8877b37cd1a3031c29b3645be3edb8f351b0382265347a3122e895b459502cb649e0e117b092723d5188f4a327a556c03c6a7a292aab801e7babfa8070b2c9f7fbb130818973129674acccf03450edcf0b4fb19b8c2fca6b75bc930d25e30234833c19b827630437662a6e792388a7501a155738a2c1a68a8830568013532b7678419337328ba97f3073df5d2766f843d7ee93f3457a97050827eec83aca636aae1a73601ae25754a95c93c79c4c86cb093cb6073a7689870b20afb23b069576db687b4ad36019d395911d640a78345f6770b167b08fccca294b65c615bc7bfc2ce5628a23d0262be61b5b19b1a94e21869bb146e1b0e3300c8ff81af9fc5b9676495d14784a6fc20f3e266146a9aff72c9273375f2a31199f1ccd09246cf86cc7a4b37092a99bf899bb5527bd03692bdb545ba999c4d692c7cab8974312530763c18e0533ffcc4e0eb21e0a4bb1ac49f9cd207b764661b9a0207bc1e870c1477b38052b329507a8be971847065acaa512343b57314bb4ddcccb51f172ef8c77bdab2627db19d4b203b79d0876d705741b5c2dc425bd05b02f7e74684d552f95c7348c586aee50079e58bc7498b06f11c91e3300869cd37dcafcfa65a93c0a458d0433c0c2e6a6648147756075c040b0149318567353146e4878d2772cb6f2a00aada5ebcec3c4b635079436edbfb38a9b2c006c39609bc6fc6a1a5eb0531d636429171a4255a6a6a4cccfd47746881c9636821e60860c109809c8580d21b5905f788cb79cd85d237a863b8add20f6a18a039a96ae6e57fd9334c5c11a3f83569deec2697978ba30b7671c61ecb491982904c53247812a2140e0721df402ee9aa150791205ae2c60710a9e7e2a75aaa4fabec268330b020a5a5b72f9bc85c0a13b9d041586fd583feb12afd5a402dd33b43543f5fa4eb436c8d016a76538ffd5d46619e1ffadf2b8b2af8d0193ed673e45eb479de5f42cbc6d33e2a2ea6c9c476fc4937b013c993a793d6c0ab9960695ba838f649da539ca3d0bac5ba881dd35c59719670004692d675b83c98db6a0e55800bafeb7e70491bf4;
    enable = 1;
    
#10 enable = 0;
        end


initial begin
#700000 $stop;
        end


endmodule