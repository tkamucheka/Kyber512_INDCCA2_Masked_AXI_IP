`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KZt/vRSZJlz5Y7gHTfP62cYXk2+BKpLy7K7ZfAycXlz1SUjTRB42J9Q7i+LtEG3bl9INdhhmpRUI
+fL2l4Ov6Q==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YqaQJhZj9idY8zD2Arjw915EBdPqsXI7iaUov2r8QConrhljtdd4rQnggLFPgUDvhC4fwlkHIbwn
DJgmKN9npYPhUIqlluL9Q9OMg4D4yXYwdVafzicPpT7j7hqzfEotuBVz9HoK9Ezr4EYUSa8A8U2N
FjxloEIFLGxm4zQZqyQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
I5suKyQBL92Mrf0qbOzq6L4hnWCMTuxJp+lkL8HjPBWkq7Osz8x00lQAvPK134QBF1pts7gtMVbH
EPRBa2wwtqIfy4UEvAcp1fHjzhVSD9G6T68hSwq1eBv5dk4iwOamxs6IlLVtbOpopX6CfGjIiA77
6aGAUdAwAQUK/EODizvXgq1wmzocrJ1yIS9AFnesQoOTjep1qtLVPABVTCZbT9dT5oP0nIQm+ENH
zFAHWrYC6qxVutY82PTK0T55WmivfsJkIIh4/FV2nMnp9qjvvRqS3KUev98WcsZbhRQgPkGKY44l
HTF9X+wXwg0L9xXEAvvCHww4oxYkvxUVST6K0A==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PhsAxzQ2BZRgVMxSUvzXsnbhQ4PZhBGy2u5EbndK8zRJomyx9gNL5AWZDX9ARuupb6LM6oEXx2mg
B7C3AVmOog4P79NfTKDWgZj7LlafIU3xcBbFMcF/TLNiLiw7zRk/bFQwz9yladLTzodFYKYOM+TD
YNPkceYiDkJib7fS4hGz0/JH09YoPz32p4Nkn7LJ9ZtDnyIPZThaz47BPpxbI6ih/coaJDsWAZSU
w1ceir/fUtgLy7Zs9hdjQpfCDnHlPSiJL6Bj0Tlcr3vaY22ipOUCyLwXTLyZtZlqtS3XPE9R0Lwq
beke82XE2nrYRoaSilE7I9+WQwpNWRdvSBbwpw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZLMJivw8rhEuOSPQPyQGI3xB9jHTtTO2boyaT19cZLjvjfxYgzO+z/lsLYww3GJAyzXz3slLpdUI
Cao8z0bJsDncu3HtQEcDIZnwJTeyShne/MayL6Rx81BZxdINlrcjE6ITwbQiVkMS3d2Pdv/P4Lc6
rvlEilSqQZYS2iXADZiqRA6ERu1S2SB829cLLbpMJjGDxGpBiUntxxXpxePv6f1eh3Ap8662VR9y
oB5bvTs5JIKy6aLtEnFDh6vyzlMen/xCBTKntIG7b9OkVoOagogcfg3ux+ZpL27ApP5+nXMzRYR6
At7bWVu9fEjzXnY73w8pddic/aQV6QAtKZ1oYA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Q+kE0mp4HuY3bfZ1LCFbRha1HkWf/rtKHYF8uonMwCVMmtIjEiJUDD7XOqpvkcSo4PUmuZT5hNpl
zK0zTNnzdSj60HVhTGdC4105xF8W3qNcB9JqaFWVMGWlRLgTPHaSw3Q9O1IHgIzvPDarFzvIOgLQ
DgXRnwZBgel+kITpFRk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
snebycTfAaO5qoTQJu9YxMcrgKrhKXbAoGQY2xDQa0X6yXiZEudTdlWfBTlkDQbKiXrIpVAx8SAF
+3bjqqGqA24i371mLa3J+iFZ9buODS4RnicaSEGNdIpBxAWljrdO5HzGEgq7hM5D4QG2ERVpHofj
E0m2OuQZqHSA5fYV5RvUZvDKcKwSTRE9gICPFi61yPE3LOiXfzx8FfaMUeS79rORytjI8sPdK7kg
WPujZZeXCsq9LzTyK9L2qlc1HIYfKjjWH4jZKYvxAhwgf2bIV9w4J2T/hdhj9Uw0ode+dFc4t2pF
v0XkOHZ2cRzm1kk7BXQIxRqwFoCI/ZlRKb/7BA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74240)
`protect data_block
UL0Dtn1KwtGZK39kGQStVnH6Fv05mXH4KVSwdJL+d94cDwKyx4BGTNnKARYwanbruMLy594PD/+U
y9NSkm/no7IVd2LbxubYYzYZS4T6GBI7M99GYP5j2TlubciwOWZSma589vvrjpYIMnrWzmsc1rdc
/tfWdd35X92MDPO35I+km0BaCS8yb0z9slob0JCik9rKOp8YLlpzY5LjaGO2CCtXE36kUHo5wBT4
Pqk7DpuMjT1GYhZGxffgQzx2HZN1zlrpvoAzkGb+WlFokVmBW3rVb3AiAye73KMj+R1rrBBbhphQ
NLSE8Vg2Ytd55tGndjHtMYkH8RZqNr8ergJPYKOUTOqrH7RWRNaNiy5K2v5bLdN+CaFI3He1Qsjb
NvCNsbdkFf1JQADMpKQMQmTdsY36oU955x+FHG/vp6JW2NuWZpaIyzyBa0J4052mIR2o9j7mfK25
48uN12K7+RWTYD+Rxi79GV9uj8VP1ALk2P9prCN60xVdiJ3FajJqB2LLYEbnfS8xSAylsKJccyGm
1wyVo/mYdk7KZLVaaFWyhD0yfbSPaX4Iix2BV4WSwYViVQ7chXcpa50QBsnGFr1jWKNWF21i3e1J
l0U25yF6zzrr68/2UP6D9hzG3yc2PAUiIc+cKmSGHM3tVK+5yEw3o7/71EH1KvA3dtbVhAXOFm8K
JCnKjVceVx/HFFe8pgJYfDN+8jic7P6cnPnDj5Btxqu8+E9WbWHjEzKU3knUYsmZvJ5FAInNl7xc
+mrXcKC2ejlAwUPTakrROeTMNfcWjycelg64PBkwl01BDQ+Tt4zfNI4BOYCRZKJB81PCd/C+JHar
himdXx4M7UPVRh6D/qUkjcFU4zy8OqYrVaxAjXAn7J6vCLOvr80V9EA+d402glX822T9vgascY6I
KnguKDv0TuOj6gZ7hTw6kkuCdnoOYj+ewmPTV8LTJXe+rHP07KRjQe0sApR0NBfmkkVsvagBTB1v
+EVnOoWIv1U+TmnhDTwlMLQYitGykGLacizhlc5ZB5Y/cVD2RSnGDpZc27ale8J2Oq5r710D47/u
BeDleqfbJWrlv36oo8Fw9V08E2BfqNu2jb7cpjBuH6to4HX4RuSW2hyX3USqOaOy/zcO0ptZgz1j
vGOGZb3qxH/Qpph4+e8UljVQmP2G4NRuSaswNWGD870FvQeBcrpOlg8wIsOY6xSKYF+vETIHX4GV
LD6w1KDMz2nQatN7rZrLy4IF+u9JAeqem0sko/3H4jMyFA5AbDzcTdgLMc6m/N9v4BD0dIXZ55Gv
g22saXZ9awoOGQ7eKXlx1ue8LMSohII2OD55ZNgpJ+xdkcqROCnIgj8St9uZki3RTy9KO2N4DK6m
t0N/32HQ0gtOmOBZOP1MAsXWRG1R96+pD6SYOo8Ea5AuZC11cZIuKT1IYZUtbsbtGDiMd0nvToF7
70SmBv6/w+/M0GDs08faBr+kubqm5Pjea4pifbr1kBRPl+x85PrstlYrwoySjzZNaGwdtDcecliM
xHJp9g8q3yEG43EGyanUowp+TFr730GdnfOcPK6bR+tQxT5Zwu6yJR3PLyLPqyZrZ6xjy1GRxWof
xOCYIs30iMmNVqftEsR/7skSpGTkYZskbTaa2g1GFCGDWnAmd2LCUmrT92PBv3QNPdHtCVZVAff4
pkLw/v3zxJVhhiDhE8VQhpqkK1GxdlogzcuYkqKrLdWrX4fcGojqDisYrVAaAoqU/+r3jQDHGudD
rXtIqjw7RL1fuJrs153Q39B0zghaDNWYLAWFCdjtCU14NxwnvTVwJQvY6SsQwDpqX1oOevnxrcN+
wANvpuFf8LTOeeI8mBYoKj/EPKGqD9tervOG7ul31ht1sMq5C08e/yE3+ZXnkRwGeDEDr3uXdAGN
8B26+oSzArnEDzLItzrcDaHWSJmk5WTjsQHd+mUBnLpoEtZJ/QsOlWG+taudvJCFkO6UOSIqGoh+
WiSwgYQfeaCQGC7RUVtBMihtYRckx5/wHDDsOeJEuYa/5Dk0A4/JcndxFJQXq2bSSOgujMzUdLT3
yrOVwt1JomLHhKuCrJjdA5E2QEvPreWO6MoAHGLLTSp5uXNtkuOLCpaoZZZ6HZCxST22lEWZk6Nq
mbb6Xs7lTAZBnmZJS1Qp6CH0B8ThKJoc1ACd10CyWP5FIUx6Jd5RBFI6oHO9/3luSy+KPKY+Q+Ja
uylzIH8cBO1QWtBW2XlXYd6Ax73GxrBM1z7/yjMbFMXK/O6Eanm5WZDKXpsiNTgP5MfNjAFvWdMG
OkI9wNyv1g4OE1EqQKwW3wwXCfmD3dIAHhO+oiKAoKVvi3ZmblP9OqZqQXm43OLW4639ccsmM/ps
8xLdNg2Dp2cunWYoxDHpLYcXdUWnywJG21yopnfC+KtngW9TfPAVxJmte6SFCQPAuA0we/wu3qYV
eOlhLN4O/a6pGXelxlUX+9BxTvEnn0LILg1JTw9DjNPcIENGA6kLoMOH8nGXjhLkY4x22nYyVmnZ
m6XrhGVGbymMRuXXg53mP9ijT/N9BAWW+Ywcu/HQwbUwxlNgS9RLmf/EDZN+PC8ZtNLAuuIu1S/6
KRAcz8q7icowigX3hzI2ShlpzZRBrYzkJEzZhblpjRpQSX8O8nLcl1OCrAuEbLjnXwEA/RYRXBka
dHcvjxitg03yt5SpQeK+/8z6FlZ+3YPwES7O/FyNJBPgutaB6czYpp9QFTkSUDBc7O+1kAfFn09t
QDGW48BDdcuLfbU6DiXC4krQ9d9spfJu5jlS3YBpjw4XSb7mMUe4mAht5lIenl1+i41Y/LqXnxnv
gVQe4pjDccNRdi4dyuEobJyz66FjZUjOiu9c025pmhhmOxLNoIe4ZQQ+PzT9N1kVm621/4fX4P0T
ipOcVBie5I+Z7wJOSZUTmP2LIp/M40mVj8YrWnyauteqkfO4FHI1inVQIeg8NxFdMYMV7mctURJS
QZ0qyLzoz8ohpzLA9C5AK5bqNcc/6MrVcu65pv2c4yFGqcp3Tlvw+aqEwmItez3PvFMjoRtmpFfW
wUh1FY8Sc+YaF8QRh1O7/B836UId3ZunqwWfMHvgR4I5lmUbnSYyWzeB7+hKTmUTjhUS5hahbiBV
7oSWd7mYFEhRCUBK+lGqBiWSY/K2lusZVewFH6BqeZ1CDjbOE2f1oHhDP/Qva3ddfG2BV/Mwm861
BGgssYliU21xWytb8sYLqc/f97xvFAl/DKnYDUlOG5wsAcqr+dTl5MmdG+rxi6WrROKtW6PTZHYV
Bjx0qua3LQB0rFeJ8CSVo7e5u8xEg+Sda8HBC0NGPWQVTTvopwWEk5jdvoILuxKXd1hAKUw/jnE5
a72/2yAGaRycpkFe2gWbbYzenG1cXcNWY+WQx0BztFL/ny6R0UscWBFa6QFsl5YtIJIvacfKGRGG
0ZTzld74gVq939J4hZI9slANbG/b6Sq7WQtIzvu0njFOGhd4b9FxA01Pay6Ie5poV0x8dc6QfCk/
ooU186Fi/IY3LSrfNzxNbrv8MiftGaTSYhhE37CpiMfiOC3dhQBFgFilqIyashScdUihPPUrLqMZ
hQ4NmrNI2Tl7XLLImsbFjC/18uRF/2SpFYkg6FWn/iOC/q6EP3KjoS2GfSvLxDApDMn/h3iFRqVv
GvCqebYW6rzBil9kPyoMFtORc98txRH/GTHyqwHVbSxbrIG6WBDlvCzVQtrPTqICrgrxzhQZS5k1
/5KQVRXqUNTITSJ0UShYBNXsm33gbK7DXmIbqL1s2Pe675r+juI6jD8060p/r6Dk9xJCQX5LQ4Js
9dRzFLm5fGuXpQFf8WinlvnPy8nA/oxC6H4UkiNzb025x+YLi98oAZ8KmY7F/B3l7mPMdZxMdmwc
wP+wCzUX+r7ZxC628kxkUSLAfwWV5HY+Wtrn5KXb+ct5Gpi5Vu6SOMZ2etr833rnsVGDonngWA8i
QZOcJt0aX424+9/GlTkBYVAIpC90M2QrUMuc1+KmPlSIe2DxCSns7wLOLRug877PbZulHvv1FXg1
dKarH6+k6kWib25HmxEnUju8z6rBjOoAwceoYAVQXrRYi9yRi0G+4ZO6kTGkk6saXXb56Pi5f4Qw
5stxEG+91VFbnRKLAw4TP8jL+xG8RCsZ/7C1sC5ZRUHALyw8IMBBeKuovDB67URnUMqBtG+EEMk7
a4zrd8XwFeXtTVkfoxZtckXVEc2JBK4X6ATWer0VGdM5BMOQYpHwiAdxDYT8QMZjAm/YG59pwBYz
jyFXqMHORZ6qoU9xSikZzVYR59utM12LELlem9ej6iwXC8O/vXpm3LcrH4ui8mfPNVE4WFe3MMj3
1dKfZK/o7ihW/GjtfMB21lzld/Ab1gZhaOBEimiXb3otvP/JIerkjsxzxJx7+FPBFRdDYd9cwxrW
Z+Y2iBiJQoO6UG7rvMwLbF4TtmLlWBP+q3TGWse1fhMzotmv3LKPKx/a5iOwAu6JSe/ERfQttUJH
yeENej+7g/SEgBtOotfo+YAwnPXtz7kXyLpjV6jG4QChMK0YS432l9FXqHDgHMGhEEp8M4nI0NGx
Bi56e/q2TNiGcvgRDJFGgR8yjKMjhKCdszQfjXORMCWzF0+t60FqrHJ8WG3Qa+QODpAvcPMohkR4
FgJzyrIMzT1LKuZYItDpS9kMpAov0iYZnG+akiYfxJmm2ejvGx4+VhZNy81x/6oRLocrWbb9h8RR
5PIFhul3niUMoDPLdsnCG/7mZDfkP7vKZ8vmRrxM/IcnJP3q5WWvlVE1I+yjOBOfHlUDEcPOMU00
ILbRv3bhZv/L6dbijFyKWs+908K83nj2gkQfMPWXE3LfoKcYRm19XynBLR6iNkYkfmiLjdIH+S7u
RPq/jYJPmuLs1p8PHil4r/jk6vS8lRMmsrUUsDyQbGhh4dUxiYM8fMnlSWntZzj3IjPZV/R4zR6l
rGGomiEc6BbukQHvQS9kue5C0ErjGVjPvvVHvp2i//JPkT6dPlo8ycM8szliysG/JgX+rUV6N9Lf
Ho5+B/2COA5JKXfd6coQvIqqLAiEcrp6pymhh+xCKhoidqD6tIgrVIdDczXZ5zRNuXmUbJhhoUnF
SO+qZlq/eQeFheW9K+yw0xK4Adv92OT+GXRzadt4qa+xQ1KNrh1KuVqVASPLAXuZcXMtGx0ebr7D
igYv0hzfYvE8UWA+g3Yx4URlqDA22oDZVGj0l9BJyHNIFZPiEuCs7ApTV9J4abpsAl9doUG1nMlQ
ef46rMNIh5fwWilcv28dQcYF7b9oUAaBI6CqqrHOWe8IJswgvFJTIA1NDhCA8KBcTvsx/FWVozR+
LlcKPRUeM3Nj3pCPg56EaCTa2cRBY1gNQFXj2JNZKEoAhFhMrvZfjmWWVMUIA9EHGJeoW2xtEo27
oFGkH8UrFYn4Ko+k/1lJa3ddYgLAjcgWyFUbAby6AoTHnpHYT9Kb4Q0ZTaOEHzkEFq/jfJ58ZOkK
zB6HV5KcHUC5IdbbGpD+hncJsSe1TXixuSAwZEh6QPn23lw3p0XmYyr59d5GF9iS+rHxW6EgX428
djCk/LF8O4T8yXf5mBeNvoHaPxg121ldpUfwSWLFNTDjFQVUUr6LCI4ROBXXyF/VoNzZZaMqWH6w
29d43fW6MxqRZ9SPRNfaoyVXqZQNrRyihS10qUjgvr2THDSJOdmkfU48DnUr+bzvke9jMJ1nf1SR
9HywDo6VSfPZDNHDWTGhTsdoE7yEZd0GdJSSUDIIPYUW3a53Ajyblp8l2IeRBGFZzKNkOOjXobPz
RznftOaJWatDc9QQWsJPdX1kMNlviw2/eaunTpnRPSkEjK5cOSRx8FlrUG5N9uL2fSqKWT+4fW5V
QcKwc/3JRfdXaRYUIarJHO2AU5VY+t19ArnVDAk7Pe6gQ2dCI+q3Nze0B+EaSi+/Ve0DsvRUOwmw
aLZeamq/GGceNKcLwuakZj/kguEjWzUEGUztnGke6b7Eh60AfOjUnUhOMXEz2A0zC7TpRmBKeheR
EAx3nA0vYMWAlbMCJu44clWX8qGQUD2K/zm97uXlPtUMJP+XiTf+coW86+xhcpO1A2RZOOGj6wQ3
1hkqefiTw0lgmeB5NpceePouSY2wzInf5bTLzLHxOQLQ/NMzoMo3o6DQzx/frl2YyFppn4Z1AEaj
ajyh7kefSZ+Zg6yDjTBvw+rPS+3fpfl6SG1z9dejSqzHhPBNAIXG1QHazA5LfLAWAywryL6JRIKD
ckD7dHIl6/qdlA8kJE3p0e2zB6WIppYX+qmYMmjfR1wJXutQMel4PW/cvXA3AL0Cm360m05dDIHu
L1LuOEq1v90puPGiIj4ILovecw84ijXelNwPOxbKbYJL7Ht4yqsUSCbSerF6NXC6C4uy2TXuRKQ5
SdfrS8mw0dp+8W1sD6s6T7qMld6+VsqOVljcOYAqg+n5FhWqS+Cch8Ssjg9Ty4oX2/gz0vEnV8hs
AVQzhboglPE4Ue6fj0pEGbm1XrCSx0dv0gucx5xqJXMOrVAzffCWXILlMkX92E6q8IQ1flWV8x8w
E9YigBm1QdmbfUwrUN04aFi8/DVcMAlXGfs8fljQB4/DVJNwCtoVYxsKDm4iMxpS10Nwyp4H9b7d
6cZBCIRQQFh+tkq7SgAwc65BkiFC7SS4Q/gfxn/87C6Np/RMbFK65TGfYnKcLuvJXYH7PfotrOeU
uEqGk/a7lmY8+Y7jiK7GpPrhwkHdi2g+e3dROPLSan0SKkkPgHkK9UQVbiRnveKBYUH5XLMOmRwe
cmZpNz7rMeKJm2TVRvWYSBoRpfcUiJMJwjzzCcc9SJtZbSlWruwTNfGtnIqPXUQYOS9ERLJygEx1
ImvEPDQVLf/OiF9RfOFZ7JoNGg7bgQHuTbX2MUkwERGAvaUusrcC819YX10hMgmuGcHM2mhADKQv
ULYVPcA0IjEmhk9pZ9H0CuSGrMmyH8BP2mu1PW7Ovrj5VpgzDByC0BmD5JNjQAscRXke/eUg6nw0
1pSrbzpia15epju0mU6G3f3Xj+/w20Gg6YK1bdXQjezbNmPfEbQbQira1gCku7Y1okONMFyZLSJo
CVmJECbpgRcOjaQuTr2bJAn9Hxtw3OuwC9dR+1F62eAaA+gE8ClPj5uMO941jcKCfn7ukPeLw6Hm
frG51EXoRynUs/YG8OPt/4t/fFJLMq3CBRSCMsEJNqMGBdiSuZKDvPnyNb39d8Ts2LXfQY4Vs0Vu
qz8m8ZFj3QN5KvZJMifVAAbN9LjtATM9mv27PcLeiNHZRryDPDosmgOD4HST8S0Wwxw7fRWIJ6VP
rAez2cgsrDpIzRrWGBEbU6tZrImYjqBHFGlwUZuu4bACBYgSPLn0wzlv9jQTKpw8ad7/ikkuFDd1
eGCJHA8G303CWZNqxp29pCJYt4TI7D/VqIv1qhVUlcajcYRKgnqORP74qQsca7t+B/VI+OGFqj9S
CKkyt0MzNhSE4K6jMOZ7hCIm2Dt3ARVq39ioOD57K+seKOFLAdlFzRB67/fjxTvU0e9SmJOgQ5ez
zw0SbfJdMxp9VFoW5dqKacPXIkG80iReVcIsJoKlK2ZIzeTmAYb3J5H5pZCJzirCaON1a4HdswEW
YKuVyjcd6CFUjf5o08DdLw5BMUnmYcSJYN3K+TKD5ZKGKs9uC6P0QUsTEYhrPyCBWVyB+5hofsOK
6ljQGjHq7CHjogooX9bwyy/G5UL2HXWoRZ0jZvMjX144vSqrTp5PjDbjjSe33sXwINGs0+R6cevf
I1FEKnG33bsijJaHNNR1YbHa81Brt0Wj3RwGj3fkIO9G90bQ6aiQKqdqh988Py0ghsTElmAWLE+A
soB1XRTBo7Qq8xALgPHTfhS9c2xAXZoqxfZIib55ker8k562c5txudaFL8JcLn8WFgGMQCVJKGIr
TZuN9jmp/FWFCCOztko1vo+rX5S9QP/aM7tZZgcP6o0kUBB5kpjUetjXWnixmMNBR1ExMpnHs8R2
Vf77ufFZv6puydq+Elm4bzjelxft6LAe6wl5kfwZRa2L2RDTKIsJJK3+BAsSfcAOHsnMlu4SEzzx
Ex4kSRShXAqVi8/Tl7IFV8Qk4HCUVnzB20t2gxOmEZUHfpuVIu1KdnlXEzNPWG6LpYXOX4QSvF9a
ESuYVhmQo1yFnnohBHoLydGofNOoV+vbR/buxdJFfzgqbP0JUKwkuZ7DYNrBzFK/g9UI8FaxC/28
MqlvyPeJbiqDYYA5SQ5CUnTRmHLrtiVilXtfbg+2WO2mRFwU/ll1kSYOfkuJjuszcAc+/1rqTtxO
YtptIW5/rCttXquUlOeP9o57K9MBY9TMitWPGcaNlFAI1NZpZ4ZAEOlvTOdMIJN+uATawq0uOcny
CKYf0TjrgNuwcpA+i6MF99ijJWXY8ZLH/qULEt79uvx+OjsAQaJgM1u4isLfL5v/Zflnt9PhEy1z
KeDCeRpUufPDPSqaR2DuAX7jCM/aiLuy0TRkDzkKRMs8/nSjBwYgqH5PavQNpqAKzzZjKG/6BtLq
F52uUNkjytSYDAYDziVykZTJ33mWPBZfbHsXhLGSp5TaI/c1i8DoTtHW/NRns3/HXuOSDW1MffyI
miiOrZ6KHDXEwXT6NrjaP0jMaYfWwkb7b3R1AuVJOUbK8UD5gBEruq9aCbI/71R95sAX4dlobVCs
XTjL3MLhARYzc/V2V1EV6Q/x0tg1Cofl7bmH8Fn5zcuMo4QqqVrAzg4xRWXSdscVaYLhas6hcW35
SkOUfcag/SQbx/3uo5n76M/tSQGGynO6ygxr+V3KU6SFHNBk2kCLDA3lJJJbq/4aRbh3mjd8O1T4
v+of78OnIfaCf7Fiok1gChzbgW6nyv6ZorXZcGwHlTvX0tCsL6msSnyD4Rjdsf81u+sRjMvHqLRe
sbbHw3O0LEao1O9cKllLtR/9OK6O1FMpr2auqmq9TleQymBrhmPexkv98Nzl3eIXPy9KdPjDJ+xH
blY5g3cL5ASh2z0nq/G+nQ0Vqa/8gX4cwxIyCVRTDHzETr+FoxDg5iU0rrjjgTBkMhE49xJs5d92
gLnk1+NQMT3/dJ1j6Jfbp3BUm6TsSDO6F3vOLzqGzucGoKKyLsZi7vEIMQQPvj8z5wO46TfIy1Lm
mbUzIrwMZo/hHNNZLJDP3sdk/xy8QbOlCm6tNa54aP90+8cvsdDdBGCK4YVoBida2TRMVbr7fSEn
kvEh/EwBbUvKQzZE+nRuqcBVyBu9+/MBVOvSqLsyoT1RqD1eDJEEdEjy+GBY0JVbTFk8YUNCmic6
x7Wigi26N1PNb2RddZwojKGC7pnpHjkumuurS2xbPCzonlwC492hZi+egA1ml2mG3pwx5oIZ70mi
fIZKWGEwqdPu9aAhhIjLF1plvlPk7HV5Gz1soUToggw4QbHlCjCWDdwmSsqL/6iw8eHRfbMBwf5E
mh8zlaMjgMJV8n1bgK394WpmCY21G8FgXdgX9XltFEq0rV2O0nBT9VVuHMTakwumSi6wJN6iXNlj
8DcqtsBwukvejhm+CawnTNSpGYpQ8lnqbPiaElFoYsXZ3Lpvr3YzbsHultMMWGaJQacH4pJ6ClNb
7lBKsLwqgFf1wzoXESEkPw8LGHjIDda6KlYa+PaL9OwW8WRoqWaNL9VYKnMnliCBuRTtQ3IdjuDM
xAbeJv3+K941qL9l6xiq0FHL5ZjGzRcjYADsokhhfoSiruhNFsyPeCrC+BwYhv9DH2ONvB8rzNkE
DjLD83O9f8gv7GAdaqcbL4hsuER+USO9boVvw5nUytRFZtugbxyX2eLmWmx+QdtEw2aiYtLsBY1F
cxcN7YTbGDJz7qY4Pw5Gped63yFXgRo/NmOaDghV5FYVo2nxhORGCLIHvNc5y1HTVfc86yTFq+ZN
vRAK8NcFAlocqYzVBsiG6NuyUs+mj3N1yqxgecBi/vi91Cge6akFDY5qAfyyUXpCRouFb+idIFfS
rhXVWSS+0+a2zYlyLAWxP9bxmysI8a6TAOqqaYt7BH9TZtwe5floil+83zVxf7gCTknMcKeAVJPS
mPrKIsjdhcZ5+iLwcPRs8rizgSEWsFr8x9VEHUBCkoKWRDVFlCr5kRbC3Ot+0e1BI8gq4mNz31uo
Bh2ctOo7+VprlXQZn1Rrbv4gSgUNtHwmFQPJkeE9W1esVVn6zGq+zgQv2JpmmHQj+bdPfbTqWqwv
wNnf0biNPRGV2JZF/MwB3aw+nd0mZ8aB/yNKrVUumabsOLlliOnBh39SV5m5SuBI3/GTAGpTVYkS
qpgGFjK1C1HLHJzJ+2pzExsRLDjUtJ9CAkEpmFjf/DKmgPHJq87lyXSACeEHuRhkvFLsXcJXEJOL
ZujcN5MEzl+89I3WSoibBTZ7JFCnhkksBlX3O23jln5riD3CRCbPBKvZXX6wGghnWBFnTCFeKfQ4
QY1bV1DEWHCQaDoVlSpnq/m/b4BFonEZOomqrkEwJyRG/kEFq+pQQoxCZ4FIhPea2alqQAJ7zUcN
QyRZbq1+oZvqu8cyfGl52DlSgaRGQW29eb4KokgExZJlSRcQi6vsJnaIU+eorgS9KuirYC07/0SZ
YFR09l6qWs73ShVJhch5wdMnMxHnxAoVX9U7qr/joBJqbk5dEEMfnu6nD9V/4zBF3dfB+YLzCF5K
XpECwJkcge+Rq3/zJ2qYHUMjFV1e4wspwJadAncWi8njAqrciHrWX6C57pXjEwF4Il1sO/mdsa04
EjkLsl0UkdJFOoUEsyTJZfDEg55grqhntJbyMYx8mxE9syAW83+Th/rrHsccefbiqQTDFIeU/BOk
/060AE1Ft0wH/RfAqft6ohFqXUBZkdbouVN57dbZx73L+XjxLIGNRjUZN4W10+VUXE9nyDPZ+yki
QFc3b2cSz21UWtyp4TLAQbdQcFG9D6FrcgiGfYVYQAJCtUvqmqKjAmBkOX999gmedDROvMEjIT2q
+LpktHcXcmbWTXWaxLKwVoyyzMzyN7j7SaKqwIUpjTv1WCvvOV61HA11IPWTFhZQaS1CRpgC4VPd
soS2s0woTd14WjeY9GXdW/jnwJK/WTlYgGgWS00cWfNOMeKnEo0/T7jY5IMlQJ0byqIFh2HNjUvo
W7BBSD3o7la2WZ3SLjI8U/H4I1cr/JYajXNwWIkMapq6yeFXzh2dANuE2SFG6qiDyuZJl1ChiN+G
W/dUUhlVGrQBaQ9QKdrgcEXi+JYqiaa2g7G2zj1OUMwW9rXPJEy3EKBWglKy3M6XQvNe3D+uTkiM
RGC4dxC4A+nrMI3ie5DFG0en4rGv2a2a4VLQDPK4AIixNgvKvCGCKh6sbw/gLYcKrtnp7CFNsrwa
geM7fNZy92UQEFWdqP49MIlOhfq/qonB23Qdk9iGf119+V/GmLRo9jivDp0ie0/OHIiyHTxE6KGQ
K/ip+vwpG+DnOxNXkDJkV3AJ8sHNsEdD2xoUwyXub8ZWXrJfsYPjNqJ4iTpB1qQY/z4gsS2VJ8TW
L10ulWNO4lgVOWC8tEOK2ebqxe2sQDAouyLJ3+iSlaPS8D3kinypk7Rs239AsvNguQdnhFc7+Kqs
flN/zIHRTAVE8MMjZuml66CyuwmyEiPTFAODVxMOBxFBusmRuqu2XkM+w2uBcFMtxhccEMOWQzay
3/VpCi326PDtpw5QdWHmwRV4dJZBzbvT7eK8QXCrfUx1cEXeGgQQqD66ZgYhOcup/OGkE9QIDbCo
x7H2rZJpfvDJUZqEGK467QalfSRqVJ/58Dz3n2h6oVb99+pAm4QFY3HC8tQwD0x/APPxmD9d2Ctp
j2Rftfn+kUqJEm4vnfAYGyHUhruONHAaRhpixDU7l+uVYfqXKnrkTGzxu0D37iC/HABM/rIm4CZs
LVjS4p4P4hEPufdI0VEgMCU2NA+5EMX3t4tdYQRMCayOt0gDdGN/1xfaseYH1bZv+7AXcBSMGOz1
Q0s0+mjPtJzW5FrcXck7ewNUVm8Fs1tmFrCDX2IYx809nBoGUY50/eRXuT1jTRxb6fnIycvPER5Y
VllNnO1CamGWzyN1EpSeM6Jd6p9VmwPmlklxQZgonp0JsyNmQ9JRg12mI4YvPX0HqHBccIGdu93K
kwoDct7+Vvb+hBRV5AwFYLrPq5KyjaGEsYhgZPk88Tz8S9WajZavqFSpRt7Qqkx96dW+enqiCEMo
ti3g/2KKVUU8KK2DZ4YKJIdE41hbORRdBz+ntsLCo0+OF+kn2SveVOTDFQRZkZUsq4BpGttb72pe
lI2XVrFEv1q06q3psY9AZarqy0gE4wkd45aXLzRed9ACdpDcgP4RPHY+TwbTn5c/emgWknCjpGgd
qo3WOkD7P7T/dPXl1MlKbvJk9uy2aikjda0BLhGc++at0X2wyvZtPPYQZ7YZDDAaSMEuaXsV2MR1
xFm1VU6hZpYLJXj6MPxpSF1YiTQZhURDXNayyTv0UmSfM9NX7DQaUiBU/+fqEgpsM+wlG/TWTF/P
Otc5kRNRwZW01DtGOHVcJJczLSaI92K9xNolHmj0sw2dDJ0DfCdNFJFLIWOlrmuFLFV7hl6T+iuI
PCjpi1Fy9ruQQO1SPvGBA9nsSnBiJXR0CbBBYEiLxMtEUCoSPpJCRocLZjq9QzqyFZMIRlGLNFJF
iDax/oOs8PdJnrrATBKOMP+5JDE4faS53s7XD+Nw4jfbw9PR7mPhyDhQl6/KljSsMApl6knoty31
ZgL4HWWZCg+IdWImaEeEfdk+FXR/vSYWdIox4NUWcnCxzTf8Tupv5IkS4sEpS6tVqGMkUKb64eeW
9QprF+ahMf/8b1FNbwrjmW6e1QmVORq8agfYeXNhURuSP0p9jePcO9W5NES4yKKS4ltSx434UVyN
QyGo+XvFlmXXcC1/Py+quNlYYCzKHQ2biyA5w5SlyRadMDzLmPR4sO0TKlmOwBpdHEr00waZr+oV
ziAj8R4nDWMS5z93e0bAn+EizSvdmUDAA523/y06ovmcRK/HvqZFyrcGSwqoPmfuyy/vSk4EPdmo
1T7aIaNd9SYfSgARP+kPkyKWTczc56k/bVsf3cHh7bdZRh+t37ol/QysTzR8Hvauj145qYwazVzt
Ks4ikcbLYGE3ezJ4s9cSMdMPIcHeHxZccz3dFN1AraA3SkJXdPmlF4wTS3TiTcKH8QWa//oSkLK4
hxwiCVAkhWznxcGV1lwB0Wzfbbw1uLr1W3dPzQkpInvCfalI0BY/nmkRHTTJV/Grwae9uBYmLpxz
teCMrTZNZJZumPHBiVa29efaIVlTScU6SNCBTb45E40KqIhWj70QNzrX/cJ6+p+06xj4l+1cwGFY
ffFZ5mls5AWQi8H13WDGzZlp1DvzrsGovevjD9QgQM47TXS9P+73Dj5Kp+xnQcXWgxMdbOaFWGya
Dk7Vw3yoapt1nbk3CCkej87/SfUjLSL0D85RBgVRDuNEnmjaCCKbwIwgNW7ry7KtgINaZTljYMKZ
BO2HnFRljK4H84WUWy64srCCgDGfiqVueXhoYlidpF/tgF1IGpnstCdo5SzQKZJd2CHAzlKuB5un
zSZ30z7OQ1DMlnZ8VPpBsBs4qvoORIF0/yp0HPG/AFjChWghwVY/C1LoZgLduC7j7cOHw61GRrjV
7FB1O7iD/62D/AHVWSOhBTOmxteng10cg9MHlnPjRjZ2L8QNZLdt3t/nqvZIgdJm+qRSuYNWLdPp
Gp90Vo9P8KkdwX5A5e8Ul32fU5V5bR0scmn+VihKF9aKzK6YSzJZ/XlsiIE+0LgXKj/CRlVoHgvb
reuishW+uV5pvj3U/xQWBmMBKr7e06TAan/n4gtL5W6DxduNxootRS+KzVbRYCUaV8+5DxjJZdIx
cHyshxwA5l+xzVVN3irwIlY7pIPhPmKKIW9pgv95Eu9QHU3PqdK8OAJzuFFho8qWJMG+rp9xfY4e
CMC1ttvymbZYjd1L6MuwKzMX+pq2LnaVI/RZh7NiKkpn1oqLWehR32L2Mq0fiZXlcqqx/5lWOFg/
vYJ14ZzypPmti8fVOcbHt/Q3SGR8nstycmS3HG/uo9VNNsk4fxYM9ojL1VqW4X0DoolFugqS0iqb
beF2NRHX/yUo9a6zgir+Op929/b+PhDrU8DppO7aSm/9yxF46lNYIa4wbWFdxLT3GkBThJ/XmSbj
0Qu23KITCoNfm43zPhfwMKPj6m0JdXybVVajVccgOMxAfeT0b/6+MkhirBlsTSNWEC8gPzjCSk1I
IqOs3BE9sFXzP07rgSRXpdRPk8aFfg8niKwHfoOCIgWCAvWHYXlUcJOLiVxkM3gUoErFxI0xqqjA
lHEv8n93oo3TDR9/GmNRXAnfHFd5o9tEfs/GajaywegI88B48LBBZU94+/a6nVdyQB3ISi/oJY9G
fxorJdgquPCNXM916ME3rBKpEhiLuyzhZPpfigfLq39BYwhJP/Qvu2P8UQmtnCsEN6zu/LiULUsI
HpKtXAnbhWeAchSZ0f98MnX8NO/udi8WvWQJhGN0xJNXOq7m3tjmCDoo5ueOkA1Sg3h0OgH57FcA
sVG5kLX1qhD9kolDWto9DgVze6dj50/zRWLAH4TzupoLqRpBp60w99X5djRLSVJFHYc3kYyK+ZbX
Xdv9b2FTAE36L4BvYpVmUv3Vf3hXppzSqLmyuD6RvEWaIDNArNm5svtNpMsbWESVrqQUPTUWqf/l
fJBrjP57DNr3xL3ftW5zkD1XIgQpx/zpW1pXwAssB+dR6XcPuqTFUt6Xl0QtHmk5T9Me3PJeSr1M
tlZTeRJb3Awfqep+H8nEVWMIN+TmmCJFqD4bfOcgCox65g4woJwjnjQTfoErTCKgDZMwmQuaEFis
Q/+FO6kr2lOjxtsdC0OS73QmeA2sxT4cBCKlKrIZigmeggc6+IPbV7BeHMdREP8qrFOpBYhShEpI
8oYEohIY0xxpJ+vUXELc9Muz2XIu89wQ0AtUx288EeleUhQH4vZGK87+x4fpot8fZ/ytDhYms7xA
zvgvgVmaS6qSeh1ym+CI6A6g/WnDYYAJWkPxxDk3I/flYqMTiALSLj9gPyXvabJ533BgHR0gHyvH
evOnjypRsohQrQcD4etps7pjGPvIYamDbhJb6e4WT7AXTpSs/1GcR+2r4nfKeUu02Pfml1OY452f
O4RyPym6ZJlPgDUJlLHymkBy8m63f2eY9ot2IC95jUxSEZIsKv+hzsXYIQSQeT7QG/2nrKsjiLRD
Wluv4Q8SZ2jXEgYfPr5iYbqts56zxZ6F0pBYS89JmtgrGge1NEp8qRz3JamoayLUcKmB5usbTZ8B
aFisn1BnqKNP4cG9w0qiEUO6gMtJtLcB+KXoHpnNCdmiy2jFOMwE7tyJ6n8coGch3clDsDFxEeAj
Qh0jvMqqXI+2m4UOntC7+VQ3I9VKMh3B7lT77fmrCgFnXAqv0S/dNWfXtYm9BPrGWMlh1O/FcL16
jEt1kjL2IKBaTMhzsbb/6hggnVI10qviaO8TJosfuN8mtJ6Ffbn6XB/2frgqVIHtna4DpNrgqXvJ
/xkXcEAuw+2m/TnI43+dzxJOC4ZjPuA/iQKD4piKdxlzAR7FIqiiQauOroiFfgbT3qD6OJADc2W8
iGnwWI2UVcAQ5Egaq5anmoJt4f+kgzO6qjlfKrW7+NgKTi/OlWwMwVNNW4SLxVC1KHRbvDCwOeeQ
UGMTV/PhKuYQOQ72tT62Rg9c/E751iAnuxtAur9Mk8ypai29V9S1FzoP/g3iJ2oHwePJ9GqYyhIl
BVbutb6qRV60xOaM5H6FFepFUSFM7rT2Z3dTXiRyIwPclBu5DWSqwLOZUId85V4U8yBCF9yAJxNN
SUlcUz5/TkFsClabtlDGKOikl4oZOPU00P6HBaB+O37sZToEpGgKibpn22jrpWbTUMCkzPp3smbW
WzP6rsHCKDEoh+arVoi0B+SHC45RoBy88+gZFFxaoFHqLs877qrCy8diBflycDWOyWKQsP2W701D
H6HnTM08NcS7WK0ioesU4dDm4M0QIQtlPf5m07hNakpM2W4zIo4ABAQhsbR0HM1Zjp/udJOVzSDI
YaIfuv09SWUOCuAmMq9k7E4WTUBzs2lMPkJs7tgsogQqXBdKoRtEFD19xHPlBULCccg9Mpf2ZC39
uBxc5RqgBhiBroFm/yprOvr9BsDP5/yd0KJQj9Nb5xoZ14jLa7J+Kqi3gErllWCO2D66J2KkGyqo
QDLXzTdeZsjU7JIF07xG6uK/mUNGO5c4hOE/Dhv9g0WOH4AP8QcgByoVMzeN/ToRAj6K6Z98cqQh
tQnWGdPKk/aC8JvdkRHZ4Yd1ckRBFfBIj/wNFTMt9wyycHHrMmmOseZQRYcv0HpbelpmJ3sEYJCb
0qM45QYGDjeIx8P3nS56wYUafMikKWHQG3YTg1neqnqm4B0zMYLrig9MN501qAwHsnv1SqSXoaW0
HsWVaUOt9hnoNz3pb806+HZJiNrsNOZfyS2gAw1Q7JcZquXuQFMihIvT12CHebh5hJNyjvdbKNNq
mEjZlnvVUW1nXDqT0O0j1SCO+Zts5KPbzsyeYYXzdUnHLX+dfXo/RifStniyaembelgmhQL40v0p
Bs+uOrMgmveddkqhnB459XtG64HneSuuiWvo8N2eU9+Lc5/WLA3e3Kuhpn+dm4fC4tcDI5ONpst4
tJAfxOcDhhXjoR2c5TC4QFnTi61tPxccrjRhpfnjWBo9bg2XcEQKJQ37KUin338R4L7/VPO9U9OU
g8BAeoBfUACFTyHfzFT3FVy4MePGVh97Ld6hpr9R8fhg5Vzp0ReMXGY4Hr29Xzd8i9e+pcYRZ8hT
RI0nd5vq4/CKO28yN9TOEj0TO9t+8ZTEnyeqEFkJqlF29HaajKjlDFlMUcUGp9PSPldgWNJts9cn
sKiuNWZVENdMFlMte6EhS/m3mrkDtTPpy6f+ILEHV1eJBDdapeP1Vg40g/jOh/j5Rx8nDIkwiIW0
uElrdowVGI1NnXIK416E0bemgi6MKO/8KJWSBFHT9a+G0p2e8nxXr+4asFsXwZkFL/2TlKzAlDHG
V1r+gh/d61SEaiRty8nwkJV4qdh75TPXN4ns907PwoT0iq/rN6sVVFaXXmSB1NAkp1KopBWTU3VA
UUP7/8iRRymxzXcRxSLqlhCEJSYrqenwLBsxe0ANLkTXVD1cZOt4v60LSJdP74AEQ8A57bcM670m
vuiWx/FExo53byOPmt94a1UOzUVQ9ksBZjihzW/s+DfNWGAqkUmHju0UH0/yIOWvcOsWAvNL9Biv
UjJUoTl697Ml1lNurL11EWJqHmS3ANc9eniKETYGMWwAHXMR9Fanssa2kCoAPlYVKbvGnzAacEAz
DAAVPiVjQ8AoHTV9IxMWnQI8ejq9H6iBnVLn65QBMHGh+G0Mw4jlO1u09VkeNj8wYoXRHFR7Kdig
YFhjw1WNMnVBxWcvI69GfHAWR1A41J/sUmTPxcFIPGINmhg0uT2sMyI9pmCwmVzbAYzrqmbst035
drD/691M8Ogbtzr/cQvLvih3lHPbDbAojaksiDeaSQjympA/OpXddRjAd0M0cS4QTodrzd7gP0sm
B93N1cVS23ekphBjJVKNGQYj34UvY9A/MqW5Aa6ZEK9/lpolRZ4e6M+S9nfHtPitJcCTJA7dkacd
v2HXK6GP4nPnRdnfXxR9EESbfJyutzB8vQpU1OwBdZNMJFDsfB9AKHukaBYWcggJzHOHnuPrq/Mp
W18PcseBnQ2biBMtfXOvNWivbP+O0Gv75+MN/jqf690NriZzZbGDP+jtrj1Ye2e5yxC6yyfrn7kK
y/lmT11kXNKXtsll22Cby5ykH5ZeOFba5dtmEA3HoRc4JNFcpX6RVwcVUn+Tse2ncmLDUCafodiC
6lrA99ZHI5FBNzV61rPJZUZulmxlYqlr758EN56YZoPOL0ruPxJjlj5WT6A5EAsuVxLH84sGneDm
EV++Te7CeTuSg2vE6lgJq5FoQ5CPvxhPhDpGwJHhxS/XLBbo3cfttAVhEmJV2cK0BuuyjVPdxXkc
ZSdWG8QryS60X/wieb6yofTU14wIMkgsqiCIkoI2VAu7+Zam5q8CA36XuaHfvwzgNqngKIjKiKwB
LSOZhaLqkuMT7dLHje8zsqcyJeiAx27v1lel34KGxhppLUTnZLRcihG0UVRPWlih0Lj6uSTnjFXQ
9ZZxPbu5qj1an7nGQlOGCosrBNsAmkvLjjwgbO8PkwFkLiMnXzlP1axZeTyzUhGMzr7PV3X/3xDr
GIEE8zkOqCWTPuqK74wuh6rs8T51Bsxk9x6PrwBqKTVA41f/CwWV/RX30PlGxb/lED0J8CTjlEaC
jTFakzSb5Ge0Jf7AN3nJ+/cfDkkW4BqHnqG857+FTAlaytiBIsl1GXw9pvN/xteynkQsInlCG6Rz
b+xlG6a/eoCL/lQ04MqGImLoGAPpArSJIj84iAokIUpodSkZSOmimBn2kOh4kFcnZVNykdCWZeZJ
ZHx41XWAu4Dc3k0m/rXUcAynJvd2wdw2D2YOLyZKBJ/k/xCyulH3qEqk1B6dCj863BRWHX2TfvVQ
5xSaaCAWURTTE/6cLpKRAoQj3uNRKINbtxFgujzlVrZc7mEBnTRJzkt0i89Ca/9LS4qkdMMeKeKu
xYe6A4VH7FttlW25GD0jL2eUNutRRkoe4u0YGzLLWO6kTM30r+Dztwec1aR8wMDyqJ6WrkwtJv5e
lLPYKTJPuVk8rDRlSL4TYapwPPQyjTeXgu4+GfZSIz3omE1auJ3fb62xBr5QCmnm7o6KTIy+/D38
c801vM4Gh82qtqtXiBF0jKBpw/veVDcnaWhySFpZ1UrRPu55D8F9+D6aCYYFpXEECL8LgeD60FsG
owmAPEmLVgSJk0+lA8iW86XSJ00NotChS2PWsCTnZZKMy52B2ySUsonpMt7wgfx7DzH6xzDHdDgF
fLDQs4CnzeSnzFk+cadJ51J436swmTkOTybRGw0j+XgboiLD1uKpeN1UnuWvjMiMV4U8SvbjqIaW
bzTJ57Hix3vek4QJP7EqXzhbE/YrUcrPuefiCmQDWhtBAvXeMi5zX2e8MA8EaJa8z9sSskRFkFCM
prIyA7T9EvPF++W6MTsZpQUDT1f8hnS94uYr0+gPmvCD0XO2z3YYh8Aw7nBYle+YK1GcvXymXfiG
xaxM1wm8RnmWMF28m3aqugbQuXPeqihbkKfrOPhp5a9xBGSE2PrYtd9RbEYjqNgcHGgAL2XwwCWF
xsA3doyDDPoo9uA7zScvHHqZJ4J2BJ86ti8ABmMvTUFNH7Xh/RNcN4xx0kyd8mEDI2D7NwzFUmbT
6WdGM0GC4mptxImkqkLwafge1wUv6ES01J9HSUJ16T1gAC8jkL2Bgn1zsVwJo0bIfPtV6Rw65onf
u8ROp4C2BpwV/p81jkrYAqqb0ml6eZ8z82mIilG0dSsaP9jZjKwfrGMIRuzSI3FPHU/mCcy3LBHU
Af1RTMDpXfPKGv5q4xRksden4ZVNZlkoA7PCkXDJeUxNCGA2csqJQUTIqVfR7TAyKJJqG/yAey2D
CBWYM5nWZVIBY72LCaXObsjZ1xiwdtpX1g0UKKalBxAyZZooBYUF/OqSwXvvx6Bga3OUUpIyIKqo
27og7bi9VQJBNtIvRVaBM9kmwymDOp05ZtEx1UrAv7JpDAJmscCq7VOxIEZmWhvsMYaW2Q0BmTAA
x5oOBE7jABFAhcDAYcf2gL7aLGTOIag9Rgz+gDsnkSHXIAcsaS2XeRZi+hxEUVsDTkmyJDCkJKU/
ggZTbjpsF5bVjFIixINKQETiDhalO3Eqn99j36UAaRa9o5Ulj5/3dE5r8fkMy1H3tI+gAnlAEfUd
KOsAued+dYeqvfLCVDPRUYJ0ZPeRGL6gtL1b3WUmsEbaby96TRHNheBBsxugaERaAJUDzQDb5hTG
Ty83wf4byupDRevCfADP5CRpAOvxPDkIX5SyYoTBnS769Qjdnl7edCNLUsdRvhbh/8o/iwYmyfNx
mO+3cFt8n+ILnWBbBF7fDfV1QnNdIrrsrLGzwkcQx3BsnpaijU8Dw1uTSwlum/tRfUo+FLlvZPTj
TPTXxVnTeA0L9Dio4GyX05lXr/EWMDOuaIX4vE0RI5Vg5KoGwbBuRDCAKUdojXhCR5/53SPmF9Na
hZRYsyvTfFXURuvEAQ/Ir24T8rVNAZ1DUojMNWmzla43Dh+LvLK9O+ijPWrR2PBg3mv5HyJGot5E
rz1y8ILEnUmiYUCQIwoz0DQgvvvOg6OF3DsSjW+L3eKI6NCOcjn6kJ8f4LxuOld6OvjpN8g8HhRi
kfBz46b9Dp+NSzDBAEJFr1VIJSV4GMZzYI+f4d3t5dbheQuuz69anB3ZfRmiMruZMm8Ig0UwzzJz
SgRKk88GxIIS33RQtTGybB5on/XpIi3sD9nDTzRvsTV5DhsP4cmlKzbNGlg89ZHFoVFmpR0i6QpB
5xdsECv3NdSqtZ2/pZvHvn1SZ4ONt/Rk0nhK4ZTEJN0+P4/x56TQcgOIGrp3407vaRMBMTG406+w
hFMaKtoZSdiaMbPx/Ied4hn2FhYQ2OwyPaJFYXwgLrhCptBfc+zJQ3qoAJZ4y7FAg34s2HtTA47m
vxSg1QBHqhz7aGtUBCebZMDV2vEIF9QIKjfXJHqoxhH1T+m568Vam/XU8PQLkw/Qp4fFOrSYfMoX
FTi8wxZJbpmgY2GEiigpclBvSGCQcwbyUvZ66M4rAltySa8uHJcv/V0jQV7kkm0rt1qkLp8Yq8iu
3ShexNlYGMF+BmGK4bXq1ExolRZcxQzIWC7IaGfYNy8uRqZ7/NQWl1r4whbXwlzZKGZ5y63jvU/5
YO3wpu9MbCajA7uCDY8xGw0E2Z+1gUFWI3U81fVEq97IAEKGZu+4vFEuohDUAxthhHI34gXd5Uk3
jf5LWYUYj6n2xw/MHQldhNF5C0NGYCG/OjSuIavsGv1G53+x5cGkparoR6x+cjG6iY2bWatY5ARf
U8WruoYERJQaEnCOVfAACwJbE58aMaPZWzd4C+nIKUcFjbkQtuzZOVRWEjAOPImrXnXIVnNOHUx4
q8ncM9CsDwrebkM/awMDS6TLpOG0pOEnzNvWr5Lp1q/6mT/9Lsr7d8YE1l+8g0YxRYNDrdDBStSY
Nr3+3nGdt9JFH6ISG53zZgtY713ADE7SFJnXTbgb9b0gIhYd7nnvjzBG0dRbKAOzJzU1t0di3gd/
N4swK57Ro1SyhzinT+/ybOA51hH8K9OWQ3Mnsv9Ww4TlnENiYPFqhhsZXaOo2Zxpqtdu/CnqQzpN
rzjYVDOSDopJMqEzgr3HynO8ekAnXRSjwgo8ZaFNmgeUO6CbHfd4SH+Y+/wBUmwAaKJwzfCkqkcv
eUk5kp+nNPbyF7MODVIBuJrwlRXy6lU+IGZD7foAEFN8MWnK6sxNe/Jnr/s2LlBDNSFnqOV8CZC3
VL3ANPGHcbYhuyqm8f4yn9lrdH8hp5kgpi+TyBwUka/qR9xKClTXnLa9/hKLD1cADGBGDB+hYUa4
f/Wt0SpVdrwI6qAUZwobqeSOFx9rrwsGfJ5h4w+KjDluCk9MNh2Y2cfslQUqGlJCL1LJ0kWa57Ln
FuOE8YKaUKeF0q2cQjz6crB4wxBRL/WTRvCf/UML8aHEEe41/d86R5ntOJ52Lw5XtMPHgvmnNGxE
ezvLC4de2ShjnS9M1ZRDftmwbIKmcz5jAn7m+si7RmdGrycyegXXZ6tV7sBDLXOPbVllV1qWrRou
iFRdwpeN0ZCxPlX1XXcTu2jd4Hzsa3C/jDLmPLyQ+YD1NegHQHrMNRGAefpG2gbxKv8O2bjJdaPa
j2vcfFpviHBxHhagDM6XHXCwAndxspBKLODfSg8xfXDqbF3068VOJL1neXIeAJyKdnNNi2H6KjU8
2sJ5GGt/yN8bJJ8iTRx7/PQInad2sVZiFAgRyyQKa15n+cHoNruboKhz5vwmrVcg9XGl5pOZhPf0
Zuv3v5gTWJWarcUd2hTKtuVY7TLWLu6K9JcPKyXwR3U6hsXsEUICiO5XjJP4p8WImbXhjE2jjKWA
l300Nl48Cp72lDL+ln4WDi6wB9Yq2dPM7wa1cXT2cDpuR92kl9cF/s8KsqggbMBBBGDkUtaXSJW8
mTwRzrpRcV9US1QNERC9bTOl2l7qLLFFKiyf2CD1KwhKrQy0kl2ybCblIq358keJheoyQmN+Iter
xeXZnRoXA8pkr/jqTo0BAp3sOESgQ2MAgh4nWXIlL848oU0n8n5zuXCfcl50wWCHU8Ff1X/01l6r
bQbJOMMyFxcovkSNG8TGolg8y0kgGAhPmMzzT+ShlWLlVYZg4psGwkXt/TXBnIvgJSDJZP3xofTd
ngXSTHAZCdadX7Ov9UX6qzLhsh+S3hYylRMzfQfpkeF+lAk/mcx2Pl4N3sIQmTwBFtpDNZgM7+Cq
YujNYqtS6addj5mQa5OZJVVfrN1Nnv4Q2OOhUXZ4Y8jw8YHz7yoGIgy8569Gw51wQhK501f+yYYR
OGpWrKZ/QmXaqY9fb11qb3aK+uBFuMRfpWm5nHJeaUiCjgNn7KsgdEGS8r7WxKFicixtLbiMHPns
Aa9wR7YQIgqLj/rxLqH3jVNrVn46XfxCEgJHNNrpVk0CO3TRIbWlDm66LL9Mpgv0cb7bOB0c5t2l
ZKABZvn4SL0yskUCGHe9vNhXiCIcyGcJse25pL9zr5C50KdNs7uJNYY0nJoSKHYF1A2Tzx4/32lc
YMOX93mVr3Om/x0mKDwECd3R7U8Eiiq+OiJ6QPOE1zR+DAM3Mb7Ly6bVgIbfrR3cdnEUuSllkqh5
/E7sLbec/fDkQPJUVGF8ePSItGbtfsSsaHsSUvTNJ46NyR0FkcCNPcpUcSIe8fEIC4BgWK8C7wd/
VEXiOHqfxqbulPR1wgwPOWT8nvfV4RQFW1R2eJUx2ouDgsMpuo5FHR5rCGPIqfs22tTFf9B5nhVW
dLT1oI4DbyBLwngaSZ0WTDB2YGmqHXPtCSoXBPYkZhtTNc2DjWP8rp1AnMTdORpmHd117JFrfzoT
y+iyBOFK+YU6y8O8WR1cXzF3hdVV+fsJls/shYunNQcOP2yDHFjo0y/svapuVRKTt9OZWwo/Mdsd
zZ79Eo+/cHWNxiuC99kJiSW+XooWU4MbcOq870dK4JwELs71BnoMRtI+bZ+XoLzOJ+Z53lK4uPIr
VTnkoXuNJ7mKEWFjxqpck2kTivc6r1Vnys5fF4gZho2QUnyC5raA4IZA8uE2MMa7/QPUmk8tcv24
5isiexx/100S/TIjE3uNaTifdOAwbUFmk/n16L+OhyQG4N/whD+qlZL0hug49eFHpOhDlkb9mKxV
3eZjtz//sH4VmQcibY8H7ZNVhD8A42Vn4Pxk0bcZIj2yFfm4B+3+JGcb8STXMjp2YrJ6D7U/0JHQ
g/GlSvHbVJXrDxLE8uMkRYDLq3izE7wngtJPTfoXCoSXlQCuN4b7jhdrEsMwNhtKhNLz+Vd0/AOt
JTEvaO7CkBCwCec5zDkIF5ZKGV52mPFyPGoKe0n9I8tG70YSmit4bwPlbr+iNuMfGQKCVZcbpl7F
5SBNY2tZu8YPrijTmUiTAbpoUJQWpQqIPoskV7klfoLqyarUtHrlZRQUlBQqiXEhjkQriB15saau
vf+oSpJu/mZscELZ1ULGkJLdHm5WUEPBHRlCk42vGFV73qV/967tNjQuOhAJNo2jGTBnvPzPGgv6
iNeUAJ0MKyM53jDFTYf95VtINStIhM7WxboM1e/wMjDC6u+qbYqkmzonbfi9XzxJagCB89gqeX7V
mI6U0VOlFOph6cIoo/NeDwZR4YgP9TO1L24VhzLP5e8Ayf3Aij/+iZgbKIJ+wUhnASdGWHYe1sZY
qrBZJimKEHZkbsw3vdzMlWXRSmVFp6UdOeZa5fYNCGuVH0PyD+r2Y0orT71aOeXCddirSZQrw37I
7tiuFnfrz+uUKF5OMA2Cdiwz0e4rV5/L7hVrfnf8Olo3EgLi++EcnAfdlYyE4n4xyhTdcj0C96PW
8E1Lqx2TtVgviTH2roHFx1W0LWvGbE9ffZ2Z01lueVlP5atyKdX70GG9Hc+N/nMwCTeG4nuWsMMv
3Rc8jr+4tReWjE0/eeOck0UUwoEyswzcVLBQDpQhRDXskmW1SEZCIcM7/EuuY9hNAgFYto4lY3aw
M/uZUSCDEjp8GMNcR9/DV/qCgIDYJyp11QdAgoEE+pLUjX7m1ZzDnStyDDGSNppZaeo48A6xknWX
0Te8mWX3J8r4Zmf7u/0qwWeb/RcyAwpDahNvmOmxrojq7bk2lvUp6Dm/HGko82jNwITQ63R7RYMf
Cq4buZvThYBvPosmTgqk3mnNC+bBphc+bwucjjmLKxLPq+WLvbYTV5EJaAQvACCmNsaglD2V+szN
YyO4DdryQC4n3c0Qcs5cQoADah9LLWxTWyOd5rZfnLk7yZW5M+EaHKFe71r2U00r4AjZbgq+6+Vy
WCTwDL1Sn43/rqECTWxwAX/1B1PXM+7WylgrOQdQqilKX9EV2OZwJlhzimQIFpFABhmGXzlaKto/
PaTAMssT4PFANHGhM27XlwQY/1A1K+/cgIz1ukemv9MWmh7AMlzbBkeRLQj/eMplGkF+ktg7biNA
KU5hcHIDOyekRL6I6Bb3nIgljj+HWhuLhX/zswP1fpDOcPumVvrPOe553++2zI3r9qAa3JyjFuN5
tvZo7KswYveerphOcl1beYAksZAAVAJKIHeDcJ7xImSV4nj49fWr4oJhJdFg9rJB++oOqCy83FKT
maTRToHh78QQIp2Za1dCGCziSCEiQV/qpHfdh6+01yuGcjm4T7eFqHF3QtNPZyYQDFmFxR3nxjHF
SeqNLS+ERuOTGlEh36VEeaPZwVLCU80BvAKT2qLXEsXi0HU7ttoniEpMLNd6g84QB5UYAffjSTV+
SwklQDyJfpYsyUqmVRyWkWjl2Zd7TT72+yT12rejwkgmfZZE7Zn3HKUtIo6dxnxEVNcPxC96ec+W
HuqGcbKTJflgesIsJ0pY56XJS+Thy2jeBCx8REecv6atJQC4wNfwTyXyCB0yjpk3AdFqmvT9ubIX
CBFlUPXyjDDRswW0U6prUCFs9eHTiie9kxn2++zcedwW3vFhdkBGDGMWu8rKszvF9rjXaO8c9QIy
z6YZrP1XpSZbo25IFsItzd1Cspyht1olQSEgz7GMZ9z1UqM6BEm+DHCncx93cAJMEakCAjie2ogL
8YWk3LQtRH4ssHhwi9blSPIxi0rXMiBHimbWmnJHKTYkauKmST58X9tsEs10yVPBlC8mbYKSFj1P
lCG4TjBV23BEnYMEJvKl50NW1euejw9w7eyYQucyBHVn5E7UDqjXAlBKMhbA96YIwG7mEw03zQR3
2jq2vvuAvX+tFyTdyaiEB1FCaEanxOXDttQ59Kq2ltTvvxgZx++G95wpmbKBl9F/K8p6Z9qdhWUk
c1vGsCnoOSoZ37kfoiP84TMUUj3ViJW4H+p9LNK3wI+zUWZYYGmt9mls+P70LjSpS17boHtPPZp2
/cvdDTwuO3X09YG+WZ+tMuq+UuTVZymsTLwArlN/Aqo6VOsT4JQTQrDCBVXm3wEIneB4/n00SJvJ
dc/uyJzRn0i+QfU26J3qkQ4Qu2HcLMdr6y6j71NDQdJNAfx1A4QbautMp9uy56O0TG9aJ+Gs6CCS
IraveSES2slCMnueaTh6nUnXD/k5VhPKr9Un8MELZOj57am9S/u5tN4WkgX51StAiE73VkXpqVp5
7bUkGXgNSc5eK6gDoE1SYeweFGzIdIrzZ5/XDIAFSO70N6r2zmTtPmUcUjzTTe0dBiWkKpvuR+7B
H/pByst5vtV3TGnqg64Q2OLcwiN7TDo/rRfop0NI+X2sIIQkDvfJH/Dxhvl+7qzM1P+IXIk2WO+c
uVSkgqp95hPOdQQNn+ZA+9BcSQrFWGgxislLGopTbxSZgQqNRD356TMLkkHCGq9Mhp59f1nTh8rg
JDRb4Qn6f7jd3QDU/VBf2+Ep5oc+y/ATbqhvlFcndbEmXVqu5XzQoBNqkcO8eSG44ekIoyKOGBF5
Bc5tvrj/ZaXGnd4z3u9NR9HvDMDixWHFECNX6qlZKxnQZcbJkOOft9pP+ijKTg/i/KFu1nAGY4Vu
lD/NcFXT8BplWbj1IIsUqoNXlpbdihsRZGnr8vcArqoyGCw8G/vqmmsKHPoAjN/91klNUytLPCJh
PgGXZw4ah4IT1aiIB9U8SgM1Mc/3TEVzfxINmSKfDZdNxJ9IcC6bL2p3K0mBTN/vTbVLIy/CLEJ6
1EPPZDMZxM9DChumMFL4m0Jjjk3mkGZ4fnB0nihFZrAWWRsoUJx8fFblV2IgCIIV2DaLZ1TqCQWc
3nFCzudeuaiEVwBQVFCm4wzYSlRKKF8MKufm0Ryx3gZsdvJEwyQRJxoM5yPVEMUn7A6nx9nV6yFd
1S4Mgk0F3eO/ckOz8TX6CZrSgwUYb/2IHdqLMMWrfdOWfRtCv7tLRVDsA8UJ5H0LkxYRx5Fk1I4P
cQl1I72dD5222g8tbzZlS/1konF+pnyMK+wQWGiECTvBhSncpNYrZcrpDYojL1kcdMwg6zM1L/Dk
UgS8M6ArrEVg073EN/pqfnpke+/70vMbWkc35P/kQCqF8QXqJ/TgUnBWQOcX1dSYdQFTd81u6qRZ
kl80u/TT6YcTARxajupXfVpXMGY3i4/Elt3qqfLCeudqhrzyPQwLTXPzGNZ27/esRB3iydeRYvSk
3waZ1TwL1SQYhtzIlFQHyoCbf6X/Ntte8P4rFONQRIs+lWpbWnZHE3kJGBnYcTlwC8MRcFY48e58
DXQSQ6JUoVg1gjRjYjQumtzrEpKq+XwG5yHkqyLsGpuU8ig/n74wX2rCh3q/r/yY5VAmWjy22P6g
D85XP/XXiR6tCdhosyfcAJ7kCnkWeJN5rSjvlfODdn92nszxDZPwuILXf8/DIk0AOD+n5uZ1qYUw
fXnKuURl0BpdLp09PuyK4J37G0UqGhelQCXuvu9JNT/X5tX2sfH07EIcvX3k0wlh8GuYCpsp8/rD
b3LzFL+4dJDDWJyft+jm3tWFPeTSnijds49btFXf9Clvpgy2lUtx3ofdG2snmq5NavG2x4Ko45ew
sPxZedD38cHeG+I3F3T1XEObJijD2c2FWt/0zDRIFybugxxy8vFUNBU3ll1FasYGasNMQ8IhzO54
wx9lu4J8mXWcsHHvcF17ofPA+WJuJkJ8GV4fuIVAbfzf5tmaxj4TkwH90ZI2N1s54mB84ff5FyFf
tAeHOVN1BLQG7n6zSurBdWXn08BCWoKFrIVZv925hs3TA4dLnNQTtjrx16D/cOdWWqb2SCmSkgA9
oI7jdBhvKUT1dJYOGPaeJVy4EUWr68ns9YiNiNLXu9Dvbz16nIBuvCTu5j7HAYdKnVM2JJEgR1fM
pXMvZIcZXdE0nsSmiBc0mpK8zaBbmR5/b1xom1Q30C6KYXCLTjBAXSQuN3jaMvUJajQfx+m+TuQr
zC8Oz9QBruAA3xPjBPzcrTVP0f94JIC1f/Hn9/pbNxTvov7LoVsnuunVdIeiJp/hg5s4Ml5bH2E6
VOJZQtK4bpVgLXQlNjw5ZuhBpuSr/PXP+xLUJ9P7toSY7Jp0WQ4pWv3AH9EDrxrxj7RUPDs6go3X
utFfgOw8gS0o260vZgCesEzfHE0PWaJbnmxqRVHnxSb+KiE/N8nx3jvHFiyvzRbIk3OS863jO88s
AizPrKRZJTZi4dQPRtGsVdkLXjcVQNNgBqyWd+r+wUwlibwzVt26XAASBRCbNTwxIj9ysXYGTC28
L7kHVQ7h2Ps6NRkB7oAskVkYOpPO6zH7ZvPjYzpf/XtJs+a/KGGuGuQ7owtamlilIsxEYh+7n2jp
rpBysl8Mg+X/y1isCt6HIf6SPGdpY0vxzGCZNumuyGUUbwu/6YNuAEBdx7Fjqz166b0w++I6/o/u
HN35ZD9wmiHDEHAbDtMgsgHIkhHgi89mcPvbZupWZfWTMYxY1nEFRjCkXMzt0RPgy+9huV979Akz
s56KpIWOAGWle/ecLqD/aWm5J9QDMW20XzwnIS8Qjo3jpcJab58uVGTqvNSnXDSoflZCfnXgQ8Xy
OGDE5eMG4hEhgjCUf+Oc5HHNpJKatf3u0/ujjK0bha4yegBihtt9lDRC1y1BOe6YJkJMa08PYyay
lvWp9qmlfeFUfmtX2ybuoyTM/ocyxboRqIyffAt9YLN5Y7XMYqiFNa9+aTEHRGHTpHQAqoUAf1NJ
d95sZL3rA6JO1saVifuBj+e7eUzBKXbdhiicbNQd0/sE3ato992VTGwNqVNWmH5DpRbJTTFQuRTA
Ax5wA/JrEy2Qj5byuMaUwsa1a0c3iXhYs28IO/+kPsnrapmbkqzy7yUlbxLu5Kzla5vTbyuAuQXr
SQ7K1jr19wilpFTpA9/NNEoDwiIor87SeUrw8fSDxjpiKVVmoZfu4TOe3F1M9+zt3IEVrI7sl16I
a9TlrPIrX+YOj6xI4sGzmCFii7RCDqPOPST2xK9Z/GUTp4YHypFZK2CCj1S3jyRLvIi1GD+wLO/c
pdWa9vfbmw2iN58fTMmmqs+IqTlrKjuxvA6txbi7HjLfipFLkYZqChbXqv5ZuCbQ1wgoybExB9xb
oQt/YfX4HSHUuPsl6g3h8Gil393yowWhv05NIHojEmV1k7FYTxMPMQmBZu72KgXX7XaKJnQTR2iz
oSebDJz52Mhgk857bsYTUZy00NEkGvKaBbDRveES1MnSCwYXmbYiXi822dQbH2KYVD5Yqke0Nlw9
1RG/HFzcGTBrM0M1r6wUYUFzd+b/+VHrCO69YqYT77D2Pc5S89r5PRlXB5G/qDTlG7vAmpt6jN65
Fq6BTjL3z4tMM0BY0h9uB+mE2NnAXMYz7ywGjTjWN8wBxXNadrHtUVCoewQLABYnGDvqWYHlMYVZ
ac2G8dR2hVz4chGrNa7VG27UyppyqAvqP3/nDySGYW9wV29bgmqDuRx+Dz2mC9AenJg5e4XQz08j
h6T+HO4+FqrXEjBouQyOly8EO4KyV129DHuHjQ8vbW0A3jljSLPBk7mMTHSkLRqqrxZ9FH9HPA22
nHbf1mnzK9Q6K0JJflvAsG0QnnfXLRjB4E0K9Hkru6jxOQj4mbYJfiA0rVUP1MdHu03vtDScq9BZ
CtGLJCXuzCs2XtYKiYL/0NoY+eCfUE1T016zwb5o+wiVmzIuyv3D+LDh03pwZ0DDBQYkVd3ZXVSi
Xf4pbG5Fg38rDuaDyZ3QI4XmyxjxDZ8sUh1QFsq+n22wQl+pymRzvdsLRMkZwjUGV0WJulvwdwWw
vTYGZ9naIOduz3M9HVorHAR4s0jBsOVKUjAeOdADwZ9HrGFiXu8IbhVJ6/R4PB9a4ud8bXHuQkmD
WFTNsZcDTmFSmY4J3enebXlCieIFtgRP67eOFFTN0GWA15tSmsdu+IFVcfkBdOhGIURPjdyaFb9y
tvpArJcBWqHNoqtA6GO3Abxo9jFXToVAuaaW1X5m/SHcls6zvlzFangdf18mP95oPW3m7sK3T6IC
3TydmJgq1PGNwJv+BAi+cRPpgXJn7J6dwQh/SixKWRA15fCDK45N2ELobBSLRtkuocXNODrZ3zez
vJf1wKlG9Ss4g+3zyj+7oxnP75yyYlCC6viTzz2ygqd3CJkXC1LxKTtgyOshLJMYY/M6ph1GgTNk
cd8qtUrhUIsxnlcmAbifL8LjM18sPp6WeYfpANh/JOEbJQ+7b0MERnWbOBKeGM1svWFDjiaGJu90
kLrkoTBD6cZrLULRx6MyzJ9+bijnJL8BYDmhAOvcuDZDtHrQGTcsx2eExmmBNwBigr92PnW8y0PW
hzMJ+TjzNj+Sg4NJ/Qf+c4Uyx0dkZb02Y1hAZsj6muVReC1HIclgwtZMsekTSzzOaGjWjBbfA0lQ
Yw/mZIfM0cE5so1Di7dxLB8nGzBkijhlS+B2XfPf08ss31lxbEXnEWwRv74rrfkJTOaFR91PSynU
prGbDEwrv7yP8mTmAmzvWuvRseAuybJDWIXDYynjNoC0rCYeEZwwvsoKOUb7oILO8uqsJ/cdWzrA
knwWL5K7Ao5pbzf49mRG41b934gLOKDFqfqK7O/il8ezqlxAESsX1to5VN/3ifqodJnEHRAAn9ZK
lno0PnpgCM2L7k72fh0GpCcYw6CVP9HvbIoeT4q5OtrWT19WdKQTPj3e6RZUVK3CmbzNQY7nKDQA
I7l7f0+2lomkkvVuUY0B8GjliWYrcGn+ZaqlU1XBGi4aP+J3bHlrR+hbG6aTP3159YSdfkYV1R6H
UuejLxv1jbt0xZdhuIvwjm6sqmB3+uj/VH+5m0rqGoCbdbOTiXlEU2Tdt8a4FU+HGI7WPRd6MRt0
vP8Cx+tBo9n8DbAftGXzpMyYJ/KYPqsRoxlqlTASBIwoucocwn5k2iYGtNAgxSgv+dJM9UMtlVn+
KnDtF7E/Ooo46Mc4Gxy0mRLJY1JjKHncsxMLg8IMsP8nhAqhapzB8hb1lkTkOOit7yAecK5Q6q3k
F+BLWUScGRug3M6WUoBJl4Oa2clKgefOKE6kwTmGqBg1MJ63Wc76rBfAeXUC9PlpBuU6xAkRuG3X
BFNx9ixnU8umGkDK2mjgX+JBO08L1kezYm0PTzuoJTfEO5SblnuNeXqdY/4Al7zAktglBvOAPxgY
ybbkfptHEfPkbcnimVPr73VKpb7m3mjVFFUGaFb3HTXPaHzNXlNDwSTt1uXmM3RIK49HkkZVAmtP
wTglEX5zGBC0532cs26RTTZMwHPG3+SJHYlDmvtPMgFAAsqW0BamBbpx7ABZuArCdzLU71XYjY6C
hnOxypgElayF7zL7cVerOGl9RjEqzY9NLeJTQRpPSPzaDFRnK12r9WD30eToLTsz7gab772JeXfj
CM49plwKA+Vj065t6o3hymNxhv38S2gNNZFtfsQzAexA1l4cC0PfcVR3poJg+BgW1EnO1Bz518r+
2Pfd5b4np0Hbz5ZY7JNRIfF7nwuXlOUF7VeyAc2712GSbH7jupVA+ufEGKw8ir4caCPaP9m2VzqL
fpoY9jZOuqFAYTc9v0oEojyv8nfjLWE/AvcOVmM7PUzLI4HtIj3wKfpicLqF4rA4HVANWUHP9SFZ
/mbop/zsXlotkuGBMUb+iooYFDtdDolQMT1QTmeK68Ha2k5DIfNoe0nQBfc0g89RRWXUfBqx/pAG
6bIal6AFJ00E6WZKKoGpxeJeBOCRsYqrammw/tq/cYYIJkkp1CwVgllMLPJtTkdesmEn3nDow8b5
45ZFV9Q1WnO6Gn9pWVFaYw6u5FOSQMHv+DQkzlwky7pZpxDlfu7TpXxG3Qvl21o8+bg0yiSwPDHy
jbVv+4NpKveLU1to6DZzwT8ZSAWS7To0XeRfDFilRmcl189d/i/gXWmeI+LikWxS1Q2DjSlEnnyZ
d5ObK50HVG10ZVV/mCQXWoDsaxUl+V9gE7GupbckQfCZJngtBvkwsoRWQBgKak8PjJ1ogbn/hsD0
KiqRaCE/QlpX7DX7PzoiMzth9h5juY2Fq429NTX2TXhdMu35rswyTb+2YtSUMYiwraR+uHEi2+AT
SEWA/kJb3Pi9lrnENN3q9E05KftKu8fYBnt/cNK4+JRwVLe7bJV26mMx1xjWDdA+RYN4LxPMm5q/
PpCTYsC177JSbUIh5t0+D1gzktZ+qewx9pZFcM7S/a0bw1oN1t8Y8D1eEmtUluV3RPfYwr7H+zhL
UPbccUJuGcuAwu1hEWFdGJq8OS3Qhmox+9Mwasy4jgb+RaP5A6u/krZ2bUSlsjTnirMoonLRzXCn
4JCXO0uPR7I5acBrpzCQitXbJU1owotOcQg5RTid41mEvSzqIBYy31X4C3RUtJFYQL5oC6nLyYen
r6r0+7LQ9TfnxE8HmZTEFjfzkbPQTZdcN04BmzR1CUWc7RjqCH/PijsNtRg0c5PKeDZAYkHz3gUN
/mrastX3Ej2M6PxFfvXcTqTHToUf95kAz90+l/K6ApEK0cxUC04YtoT2ss3BeYBuVDEqv+GvYDZj
tHPPrgHwBaLaOL6kFihu1hea22jl5u0rKfXFG721rS9TI5EkKwS2P1w4eI5EuGcOZ/R1aGc97Wau
rMV33MWrocy7yWBUxY65EJj7NCS3J2LDU/qSOOc7dl02n4yZFgQaVK5okdgGngRfIafWRZ3LNYrL
9W8OlfJw9+5LtevsIIgkmySqpNcVZCv6qioPIk64lmtNInqf/lD2oXCx8D7oO2U82UA/RVEMQOTg
EIWOJMD3s4jhMGTqEDmHNGR2T3VUZSQYaYhgnUEYSUvZRsYyQsUBeVq3lDPkfaDjlz3T+eM8Mjh/
ZDnIon9SHKXmzlKB354dIQh6YEuRJ3R8V3YoIcO0qmW0Is7yRVKZgDbUjbIPPChjJyKJjuJO183I
ddtpFmAogiGx7rfTD/xyBFi5hEBAmLUXIsiIXicQ5fxJKZ0kR89nCYGwh1iJPRnKOR60HoMBZNxm
LhIWgIAhkRmpfQ67ozbwGJiAsejRjsW9gEHk6qZkxhRMdn8si9fc6tjslIF5cLPVF8tFYFpRu1FG
c4cR4VF/Au+dGgJV3WzWVpn4M58V0uApyHntYogHH28JWUdTgByQ1bsLds9GlKJ5CCqbr71v8mjp
TwJPKaXjIBi6ODDMNUXcA0QKJvLDenSOyFYdOu3tv+bHG0c9P3q0h20S7Gms5AAhVR0VHqnVEBHL
+BRyowW3QcaQEKlk3aiy6EIMbQK5fjsR4uROW373IzGWuktnl5VvJRSPJWhLyNeOZoulVIwgoXUx
JlSqeawOop9HytWgl/J14pNbqTwH/tEwacOeDlZSKxWxPbB8iSIR7G98+l3ZtQRu2uNy5aqvL20V
u/gpcHfu7Pnn2UvkjfEsGFP42lVe9JCMAdUsAPRwNO+AXYRYqAyK3qWiWMsEyoPhXDBVEcL2U4Ou
h4rTFiJ41QC0S5BkyhKbADo6vWA7WW8HBs9MdH/vSZbWVJO8sulHlivGEsIageVgfKtRRMbD4XKb
K8AakMxLOvOHZEPsT8rm9aM/IvPHABtcqU78NhWuhJTM2/A8z99lvkryHWyUbnWS7rhDgjhmntOn
VUCDcy49lKcA9D1w/nz8+hBrV9RH366yeyR+C74RId0sQzmwowYQhoT/U+bTtyJXfHbi2QWcyEMx
YOBCmqBSxlZZdN33LOQ3vAH3ehyJFQkj74Rj2nh7TGanbXc5Kgu82PEzY274Rf3q4j7rdExP/YM1
glwc6wBvTqdkb+5akMKZU561t3YftY62yfLa/3UzLdKGi3vSieWign9BsoNpHprBU6Mb760HOcsg
WfviDjfuV0ZMvRbiYWFCiFNbg96eI5IFFWyysMqok4D6ugalCD4pgvdnJh5G4RlTmaAzw34eE/zX
3uNix3TS3t7+GSqipg2sG0uwM7x8ysP8DkH/AkvsgYSTUjnq4W8IR4vrbhzJxmwPy+KZ9GfbBBwo
8dv7qQ3MEicBSiM3Mkz7g7YYiBmufK0vhpf/ooIsmQaHdlrfKpKAs9+KXSqZeH2tpN9MD0bt1SQL
C7dbjcDMKf8fYUp55nqRyVzyIAfmSkEZxxLlg1vZqMOQvoobRnmn/mPhoShn4h1BI6Kuqcmhrp1x
tFGxhkNSmmfGIyTPeNFMZ+cNbfgjsu85im1aaSEkAFMMgUhZlWRqWL/5zUn1rG5W5fXSkQ7IPWRK
OZHcmFvxjlPtgPJM2HbdnINDInNv+LZei/k92OB35LQxqggdK/zpYEBX3OLnfN/3VdjQ5RUVKuI+
UIfz+zWo0gyja7dMDszmZ05/6Qd+I7aop6zJ6cl+/GHk64v6hTvAjaPfhbd1D/9x6B6JcDrGCE3p
O0NgRG2wLnYdHq7DjOrRWt9oDk6owwoTx9fKN/oFvAAD0Kcrwll2v5eSOh7+cUB3bMz6o2GhW5AY
XV1mPCHYjT3TgOm0UgQzkmMYx9fVl25peIze/HfwILJQfl9npAU7xYKHJ2wW/FOrvOJachF7qfHV
cJo9WIFof8vlH4a016sdltN87p83sGK/haor7a9/9OW3OQjub/BlCdFxdTCK2PwE+WlATeSdX64g
YnesAricOpVLfpwT9XmTmu/jtaXHJ1ynS5t6K8iQ7REvB9DBT1CNLEQc2JPJiFVNKUiqg2Vjd2Bv
cYFCcvXBA/BTbyZgPNTxIb0rqidcWrNNilSgiVgle5C6+vZTBK+4ErPl/KsSrcMgwdZaDDgj94pP
TuraRJpKU9FDNRQA43T0z1deHzGLD+K/vaJ5nudQ8yHcxGuEOi1hd9uLiDdbcBFAaJMxQFbfqTI6
j6gTKrAvZFgrTo211ytpk76Mpbu+LHNDCzKGCLbqWux4qRkL09NtW5OStyurB9JU4vP24JwI4hoD
1OLSuuXnIrbDb2cIaA7T76/Ps/TkxwmNaAoxvWlEMrO+tzPr3Z22bmSaQMi8cPKDw5eLNx7wmdj2
qk114ydFHACCG4FZLPPcukLgx7hDMsZyLfpmF8SeyFiwy+fnEgKodkQY5btP2gOK4A9eRwrmAipn
sHbMNb/FX0NIS7/kks0wImJMr0brWG3AunvX9wOgU43bSgMUF3hT6munWQq1eG/YdoDiNk4nbAL8
BXjNWlpGnaSkh1VjGNmHKYbRC1aGfaBuaq0HLkrA7uei5r76n1FA1WL5rohSWV0hrtrKZGHNaEiS
Qon6/bE2JlqeD++5qnhZAfUtDwdfnqOR+Doo3QtsJrLxXgUCkiLt+lhqbgVJ+oP2H1syJXa3Wbpz
S2GSg3v3lU2lun614WgXm1jrIpvExC4DLDutJfcu6kA4Jf/IAY9T/z0sFU0DWCIRq22A59DnhRYx
SuVYIax2e+kNAvnA0eQpB1GrWXtLyt2RRDX0yC/hX/76vGSm0h2Ps6rSzoP+b3b9EpqPrmbVWmF6
8lFbTMAjOWHNPClI2zKV9DDvzI5/uK7KrbLOP6YfQ8pKF44CUq+fytcdSuEzSyir+B7lW/OnerkO
BA1w0JHi10I/B88v4jh60ajJUFxaX+B2Dz/mfZ8wO7VYhRKKmumb+pUkr2gx2rAF/U4lHsDrjEWR
n+VDeRBqajwGwHQUzn3B7mQK+4Pix3x/DD0tSx5UOZYXV7UXPrrrjn+o1zHibEhqMCR7g+mNgAfR
GeIo0oS77a+Q91+8PWv35PPJp1WlUIvBukKpvUbDp5ms3CLO5pgu9rGr47QdJEBuHFEGBVPDUfRG
E/uoQ9QcgW3gQ9zldA7o/YRmWo1R+KnfEvYYOyqDjmPTPXxeK24Z/UlWXSaqnXfPPBm/n/Prm9pk
jSU3nE0lpOWaQTqhyEqXlrhIbjgFzlEzv2HVuzBfhorur+9+bweV5oVktRnvmQ+xfpaP/pexh4Bq
6pFA6cFtqD+Nkpf3DnHgXOIrolnr7T0KLKXNK2KeWacYVYFSCbOEAmTwAsbdM0OgbE2S4vToHbhv
MjEtSHTbSTU8JOYYyo1fDI+gdgEXEAn4UhR5DiD6cPq9PqiBr2HSyIR7MDmqJ7/w68HytkDHBfsV
AAV3fhcUoFN+uLK/Sl/v725wzgw2Se+OOkJAYtJK3XoevxV75GjnLEm4b3mZZyK6i1tzqKsxeEH7
eafKE9CWrEa4MsDyq3+855FfdY9It0jiKTAhrZYM26bqijwj6oOybcitOUycx24GKRBYIdA+HI3H
r8569KUPa0eUdN9AqgCMyOv+vyRCdgoCoPffFOLJGjpW2Q8hQdN4+F8WkKR/4H88lu8SX83/VzZg
pUgT7OTCyvzcDZO+YoP75+eZ0VFbH7GVTHwSojfs7iDoPmk8pZ0oB1IoqTCFUCwbtyatk9btbF7o
i76GHzByFuyxRqnITmitrWBM8HIVSZMFCbpLeYOI62hlxCBgBEiip0zDghMH+H0tmVDwRmLcNiK7
krImkLtYUtY/2iHUht3rfjTWaHxaGPpd3gCp/OgAmmm19k28LAgjutWl03xynEN87LBI8XpzaPAS
yOq2usF57WHXgQDlGXh2uXSIP/0vvqBbOxPyRehbmnF1HFd2Swdlcr+gN4MIa95KkGtNJYi2xVaG
dU4ctb22ikGGm451X5ohMtTCakUEUjeNrmIjuD0dYf923ZCv7X/vP3FuXNZTtG0kWZarJAUw4Leq
O9zvpGyqLU+rtRexx7di/LW6/4uzaUleH5p0iP847RDYlxe6I99qm9Mxy9LkWbawn1TKq8Bjx9rX
9YpPjP9PZHAbGbe/724qpu+m6oNteYZaM1DQH+xCH0qX8KL6V+OIZuiThHeDsIakPycw7yHKvZ/1
6Fb0LU0STeR6skR843SPx/VxM/wuW9w5evpqUYXBhaj4q1umH9F1MgmPosUlyHIU2IQYuwz8gGvP
Yzz/UZqk53A9k5Jm3yDJ2QjNyn+0dNX5u5kIwVrQZd4xMgH1R+nJh5ygbLORmxiQxKr6s13Ejg9E
HNP4RHdWzl63OB3wrrdeHrMgp4njRltbE8YfVCt53BNqmtsJA0i5Z85oRQPtMqrKhg1Lihve8y31
ZTEM+OqxtzM/Kc0TNMwQrkVwRNJ2K1nQiBh0XJOlrPA8p8tZ/dPBUGI1IwRUhAwykdnaF07ApJPk
UctfxB/8chzLU0ktHJe98OIVM4LSfWcD6NT4lLRj9yLuklxD12S+Uj0nbOEicr5ZZ7g67D8ABfZ6
xjKGvpA0oyUZnNXSV9faIb2Bft6RFpP9/x1TC+6z1r2LQISAbIeLnZyadUWqSmgulIooIvLsPoOI
GXow6U0f0QJ9QT39X3TOWYO/Skmew6s/1BxaaRwXMObxolpsTHoXpcla7nIdJrjNEZn/eiKIsSxN
Rqi5hv3rEBXwiaD191nXTG7+rv4YXH2L6ZABzdZVesvKiHXY1y6l0j3RSjkjTym3Wnxq6LUXgRSE
TUUQCREiOu87KExd7V2ojuTbDw+keRI8UJcurc1gW/khJvJ+FE7Jqx5maRBrKoNgZlt9ggvMCk32
oldiBBHUzrGXIiWFH/tiA+AjjAh0WYqwpEAoKcaqUf5IAgL/hGEjx4hbD59C9aOGTSP3o2Hm3f2S
j2cE/2eeJFkyg/2+XlsT6PjmG9KqL0pp/5+cPMeMTiN8oZEQcUJgb1NUZEHAakMy0JM70hXCWY9f
qQmMr2LvN2GwBCEF1qjpSEwwA+PxOPJ79wNkFUlB06A9ahVLTsLWY3lxyfkAXHxhYF0MjCBUliBk
F7wtJah2nJ6VIwK9rHq4rRsA3MzBKTMcSItMYGooJjWfMFJtY1odPcbzhSmOlzIDBCle+yI4A0Nv
0tEF/WcL44Lz8BKNkLHq/y/v6cBYH5rYMmcUitip4+hoPr7D+XEA/z94phzfxFJC6Ox7bQbuLCMk
qcva/pCwBbfe43ifO/nngQbvuSAlikbAPH7Zaeaj/uzmrH8GoNG7AGrOPIAVyXOUolJU9/RLe+1l
r02W7JDOBPi7RH604BwyT6PBhRFbh+b+4bupz5kRf0wzTDJwyhhyx2mXWzHz5bFVpCRC0zz+ar/g
pgVmde6ik9ua+3fHeH8FRh4HNzgp74d7EfWQe0DC/KEDsxXCVDL0qZGUDYSnqaKqCpu/pqdtezKZ
1KnYAI2tu9qP4IZYrSBUSpA3sLu8Q1CFe6srtz6GNrWUSwFSOgVcAI/4CW5nlBHmNasrXObfzx6l
MR12ResbMUVdkrz3k+deLvOLrqAycQYvQlKuwNQ0JK2VTQQ4qhkC1uKBLLuvB69FDY5c/9ZB5wqV
gAJ2bH1e4ytsJVXrHD6UPeVBat5eBJ9WvnEVxOHISU3QC47aig/vnxYfmkUj2q/aZREBtyylzUFj
1mrgzpLnJYp8UQqb18XXHiSaJ03idvFsdCVaUvuJ7cRc0PqT4eLl76xIm0TMNl3wi2rrKapyN/fw
OQ0ivhJaOJILKfH/K5FFDcJo82spi4weqS0o/8SpBY2SG4j5VHy7RsJHwPnYKKzBECttKiX3DGAW
etg9uYzP8Ltb8+lpnJtmXVkPDLEv4Ni8wa6b8idGSTQVuCDTUYt9UFktejncQLJGQAk7njSZl7eN
fAWirjnEr2ZJqEBwxKObqLlxj41Veg4kGE2gdxtMiGgWZVS5yTKZjycR5QSGiHWMvOGOuEU5HGxa
OblWZ8M1uUHJiqU+z8mQL7p0oQrubC93K1IyaK347BCg9YEa/6/c12zht5ab99VGnE+hKLt4pkHz
yo0bFFTEZ60loVAxMBsvzG51alFqVyWRUj4RJqv5xhHPVaVYDqMAswYiyZA33sIoqcry3tpCfcoT
Nf9gu3QiyP7n/PQ4n1KEWBGQUnozW4bQRDLRWK3+rAveg++gkppWVj0DBWNZ4BORrGySHvAbeJdQ
xqP/6Cx/YihY7BdyCbHp64g74Cg2EzPwzYKzMrUYUozCXevn7mOi9WJUVn2Hj9uUgkbHq4TDqyOS
sXSO6egTtU+N3VViiWgBfhnFrhF4in83RXBfO0JaCnmSSdqGOJSHEzdhmSsaCFQ0ivjh9N//7xwY
XrLXaUTR3vy6tmPvxO92ttZficZViR+T/wmBHRNUkKpSFZx1EHTMs3zDjeFsyxDoDoCT1QW7rsFC
KCJYY2hx2UK6TryWAA/19791mEiV43iUZGIsd2s6jVEQlc0ilrIbJIQLNzpy6WNabtbUWlfZGN7c
qTz6sg8CMwcnzNvrkTQH5/+8D2B8BIJ3CRQGXEX6eDpMrvAvdorbeeBaYTpzqctZPle7eL3e2XdH
7KJTtkIfOZd87hx0owVJ1vZ4toSEwIgeI3N8/OR1JYgEllIVJYR7baMXS7G5/DzkAC30Jt/RZfZT
0fAwX7Vf/pnwRKIojzYfidXDwU8D1fBzdmAmlB6JxKHcnoI5VQoX8wIC7KbXb2CvisfUkOFbScJk
48tN/Q71Pjqcw+PIU7cHOaqQ3Ez/b+YBbdx/Z4VEojg34IimFVnQyb3ljBJr5lU2eftOTifeS7jr
ewa9fVSwenRkw2L2iwaZuJPF/YxlRdYJt1Jn/V3cxvWxuv3zRZl/JQ7B6PAFOx3DAPtj3ih/Yr5s
0gNzbzLqElo0sAYHEBfyR9Hej+QLIfaOX391cz7Nh36LfembzxA4e+b24EVq9WUSht8WWc4KvtQD
z7WaIKBjbvlaegUZWSW7mwSH0hvy2G8QSYVslQUmKH6upNyF7o00YXSoQiJlf+9dGyZ63CPk1Kdh
KkBOlJK3w2NmVP+dZwoNsHDq/i88f3JVKkpn0KP/59bS7CC7LUPvlAgpnZvXaZQcPkJtOaYmooJ7
QkEBXfMVtRlhGzaKozZ0s7gCnoH64s4bMIO2S7IoqBJn9HveQwt17R9XyWDhG7zXXfPt372M5ytR
PhX/19hMDwVt3bkn0MT/3W9VPDtqE0Ns3XiCv8xCMPeoyyucVbo6l0r1guPBQKRLnuXSzhnReC81
4nzQPF8yS0i9lk3RJjEYs3iWxhKF+YQk4UmhouFuRe/ggqCGVPWmXYeaq5fhSrH7CVsHDcII9TOG
84DCESHwwyHvpB1ryXDtRVqvsIjGaKXZTKbJdKq3JG+ZEfVxGDuv26XCSF3P7Vl0mtf4pv9n+Xbc
yTUjeKHEcsgbc/DHNIN8o0u2HX6JQksgvCRtmpslb2+VBkkoSZ1vx3PRrBq/JrU53yZTtDLV/LyM
dIbowOHI3Vf/DvpOVtToYojrgiMKe6+VOUlkORa0jUM1mbdp0ZikZsp6gH35K53SDM7YG45wOAH3
MwJu9HE8wKNnLbEOUDq+pHbY88IVWHyrdWzpYaX7LWeiP7M5e2yK48SZKMpRVsWjn9Zqr8S5RD4Y
Yy1JMCyEzHWhR20F7XfNvlIcVPUpfuf2yJj8WuFuVSmEzKc87k4h1UrNaXzSBFRAAqLnKcfSbcpb
D3g1Vfk2Uar2tEOOve5HEsaGFJJkZSY69Z18dGSJDD+iXRwTmKbI9/JAcH7t9DjHAj7mfHBcUcbV
7gSZp2fNy3DEGc/DnlX4fQrWGXmebWrhErT5YTHDVfuCkWD5tDBcSyXQ9VwX9WNJo27VszE/RblO
lN0Y4A/kkJkdHN3BQUIpLfshqasgT4B9u+Mu3TX1xr/MtvZ8peG08oGCnZSiC5Zb7RdPjqJiCZSs
yVNeC8Mgr+Vj1rwh8WDyyqZYETkDuatLxwLxVlooM5DmYD0DqxvgxwkqARq6xjdRMRZptlMWM33A
GnX+PaDSHNXWHTFpgM4wUxRd7BKQe57LX5TawhWg9bXBF38nVRw95G/9Ed/cSMO6jZuyAnaZghgC
XO/Y2IsLVOrtqe+avJlAN3XUrAFgPXQN58Wt5ya/MdB/wQV96MQFsC+5c6Y8EsvGVrCS6a4n6COk
I7+5KwlYtqdv1EYgZoKa1l2wBWTtqyHbu20b7Sc7y01W6R7g2+JkdBnVuXBnnNM3WmVvga0ifuWF
8D4Hxn0tYOajoPD0HFTTrMsHm/GwUI9bpv9EGLZc+tV2B3hVyMRt8QwPbW/ZymmgOMn4RNUxGQM9
OvYLtmN8i5cEng/EBKhRxgk73U8HDdiUMN7yUdPe1Y+zwkf67GjyHtc/dARIgv2x9EKiTqj0z/dH
B9S89hOObAHeW8twNn8IbxhbwHCAJcp4EbZ3G/w2Jv7ZrNVV0ujlenPxApuS9tvZTAXmUMxwED+6
YCLh2mCOH7J9MRDB9YdSzH81SYXtI57BtChyRM1ZHZnltmE/LCl+yS4QCM05+uSf6RNFnffRNx2b
LE/qlyCboG73Wbe0OZRwpcvk6xncgcov8ZlBCh6M3A28xLvFuXRwVnwtrZsc5tF0utcb4iE8YVO9
P2BwmrdnrDaNOgy7ZG2TERqTdQffjN8cPBlq9Lw4PpB6Q76dXTGZJoUUCcC8YTjxUDu7D+64dbfc
/qEi6MLaDm8WWfaaSIOMJTSOfe482M0nDHDJcwj/a2niuQvru6+bDcmxuLJqJVdEKot8esfrsdmL
gwCqHZEfolp30406Vi/169jjwyS52uterdH6Uevjxc49QOmYrusCUCxFe3EIpoJGhDTU03ixmAra
TOQqCtZtpiVGCkN7arVRs7DHhDq9amn8dguT3LlvVK6e0KRaGArbrbwog5vCSvVFhgG53k9AD4P5
rGTFYw357j/cUI1HCRsgYlHFyKTxGLGTNZbykg0eJ0X7L+yE4OzIZC70BX7duKYIEvbPsE0GK+Va
gzcH/R4VrToSmJvGK+DWFQw52byz5ft0oFUFaCs8cKtV0qNZjXKUZnjpu8hAPuQ0fyw30vKCwxCO
YTwfULfURzfl3pWS6KmOmlv4C2xmIFzIUgRKqTVGOmfmYvDua2OF8t6gCQVPxQEEv2pqHT5hMLkV
9YZkedeEhscap6Iz6mNgb0W1g7aRbZaB9IM1ciVEOkgpDQOmoZzGWQ7PIc8mXPASxuSEsgs77kmu
/qmUTkQR75xZisZMi+AhzciwIW2bO4yMhCWanDqqnAn1SsDi2vltjVNhQsQnzt3OWGNnBBm+HpmI
YZPh4/82mdvENk9c6IHeZl/GBWE1TV57WMwaL4HUbjIL07+kzlQ6CywnyhTPtj8oRxJbyaEKLPu3
+jUdGQZP1qOcbN2XbCmd3ZMTwXun+LwCW7bWD+IFjfUaTMIT0P7vmf7/dQcpfdIyF7Jwf0e65iMQ
f/vWWW+ONk+SBfVnGdSdI/XqYbRitt8rz3B8lHJhA8VPauUToktN6ExvHstNAmzzasPVOBU32eOo
lBG3RljDYRxDdjHcukUyrbcT+clgJR4gvzQASHZaRPypXCkhMMWy7WeocWBWwDCBC8gaLyeZm95o
KqnDv5vfp77RWjDcOTMm6RI/jTgnWzjgKomrmWR9nTAVc3i8urYCJ6bHYVZFiLM1mOhSnliG97fW
jcxnGB1OmR0926F8IwWnibWDTXX33mhlfgpmm6CzBos9GZ78LxzhHTtskaO0p/6Kq4zUTGQRmEa9
lDo84TKKKB07YiwcfBfE93VPeLJaCpZAii65P2dDPmCCVKMgZokKKIZDIBAvFFOD9pFE0HaNiuUF
HRwFiPhHfLsL361tYwzwhq6MTkFl5/ibAcI3Q8qVSR5sM44TdL9bxPsRalJjITMpwfk2+HZ/TkXl
gnTh9Z9n8rvNjztKuzNXW1bzrS02jaRPcJnkk8EZ5kKV1ieBmcaLXFrn6km919XXoYoPjw5y7CWu
yQWzXX6IkFV7XVdXoQRD57guVdQCtCSR/B38BZGfJovbNLCi4vH9WVxUAaAgTgXfhY3FyfZgoRnz
OVQCzPAamdWycALQg0SWeetOagA1/UAA+D32WZHapNdG9WdFZ9GfOrDGtcVVwa2oRFGtxTqX7ToC
XieCw8uDKEoU5VQpwkIBvuJHlqMVfKxo2i2SwaEQtvo/67OmVgf6bJbD0nprFJakjySbGlHJ2zjs
qwI8ZBqb89VhEKyUI1XeuTzYIffslrs73uErjeWJT3LkPHVfjnBHJQf4OBLfh1vQfyHX/FKJ8Rr6
pZULJ8A5t/QVKuNRBXn0ykO149CRxJ2cnNaedmxhf+v6+daLMjL6IwuHkZKx2MMl8LmFcZEHDBul
PZ99Orc62E+DU5EL+ObUzOQd6oQZQsOAJ4RVGdwMxM9o96DvvW1JiJDQ6i2R9pgbOcdNP5uEyIR4
hBU9Hen40/uNDuZjblZfkBNxMPbnCNljvjO6GzsruOCXKni7qGB+gKZKNtlqJRbzkeGOWCBKW92O
fuBzpp3XyBht2xvRLBfZN6u0uh4T3DHDvWYqFpvl8PQsysCoX5qRdcQuYl7tmS0UUMLJSrsTJoG6
lqkcb3pRmfJHvi5QRVr771FVGda+8LmvljR2zSqCDKwSXQcD9WWqfpV4s8/9hgvxPLK45JP4PlML
ECxHOTNHtLIDPvcwN4ZJgj0/9Rt8r5YtC+1VV2JHAsos4+MoL+mc7GD6uvUE9bPgM502YqcGU+cm
2j7K2kUqgz2mdEO16hh51eBLPGfs6UmH3aQOiPRS3QcjfSAZllROdoMpa29IXFGk8usncjJUm5eQ
kNee0o5IVYvAzDdqJhvb+MXMJ9oMYbDd3JrNK6NB4bG2pZCcX2WF64Q0fOT6VoReo8TOpgzY2E1p
odRcILR2LNBUGzQOXWSpt4m0DEqA08m6t77r/FXzWVgvuGwU3RjcZPhnqXIUCzG5Md+mFWTgwN10
29jM+2kqWTerN6jBsSTGThBPR0YnbxOUOXnTiJdbhtY07aazy1+56B93iJCDzHB4WIkRehvA7XH7
gg+vk9xigq95NEPl2fIPTig/En1NFT2+bLrJOAzG63NeFkMs0FA1T6OGggPdXWYVWYhKwTG3TVes
rRnp8QnYgoysYTi5v547x/wkGZT+hG3c5n+hrYLKXWynftKvTfPO/oTK8Rltl+ZJ/UogWFVmgoYZ
ybss3kVYTyuw6QgCj0+5Ek0w9Qu5HsI0KAIBb9/chNEmBueI/EHUQvA44FrHcM7G2Gl5mtUrNXxQ
WCu2EsvbUk/Gl6CPnQ0Zt0IYj/uqErZeARVVYME+54CRFkrspYwJDpMqtKRxPE9hn20/CQT2UplD
Smhiv3FXiD+a/11lRzgizVZJj/x/dtnUhsBaapKiekvONIN1mr/NJyi+LLyESIaQWFbFtIDiH0by
8ltg/mAvOEF2NOr3/p8BT8lewMQFbrhms/anR6X/FMmI1B3+gBRuPJ9C4zVDEByvT2uVBh97HGKo
hm1ZaVzK1X9JXXZcKVbeBz9my/BL2+6GkC2srw3fUuN28WeaVElR8FPj1/WV7UySDSBFvxQzidWl
U/Na88R8wXMS/WyRTzV8NN60sybybIIkEJbQlBgO+B1CeAUTvRBOSlIgNZvk2285iyl9YgdeccL7
No0MWsjAu1IKE6c2/9jRzGkl8om6Vwsp/YDrkKBaX5bTw5bsWayNxOEU0ihbDE7jH2BPYoKBQowG
XMSEx0xN9gquKWvZAOF8uPTYvhRMu4eSwPUoHh+zA2K46vRIu3mN8jadoDyksS3GgVj0Rb9kFXv6
3nSSx8klouTG7hT8f3JjMyWq3ar1k/6pFCRd4HydZiDsMtAsYIeJ1At97cNAy/BFb0Wm8Nq49voh
o3kinwfMi7+X/IpdHNb0skqkBFElsCRJvbYqDEnRjag1ejYj9mLgjlLFFF0iF499wRuED+0w6Qpd
VVEzzOJcwmBZ2FF/8MWduw0ffP/Y+7k4GCgb0Dax2RYcFqSewopaXZVefWNKbwnKy0LCMlHcZGA1
B/Z9U+2vB00AaN+fzkPnYTlaoSzKPArS/aHBb8sE74PHNzmPBFdaDv9BLpTOvWNZDZ2YnsO7i5f8
2cxL9K+KYwDdBAYA7s3r23VLPsJiF350TbTdyni1yLsUufX+9efeGyIdxpSuMrW8ArVN+ADhnY3r
RRT++s4Q5Qkb9NKKfYKfgVZ66FV5QvxBJ3zmYb4Z5i6xXdCAw6E7T+jjEHZwxPAluVRFct5FJaqq
Lxd4G5yhbZvYKLZ6lRUkp+w1luor7eOv/fmHyqNgFr1ZFanQNRhmndTXzB/Nq5Lvg/CIKH7G/RpY
PInYNydp+GEIrWSYe+lHsK4i7U4/yYAIwWCBS0CzzR0oZfJnIKMsE7IjxS2bEBmoSIOCGISUESjz
eXw//KDcipb6Z27JJyjauu0klWsCcGOPoh3X9JQlrXcpfY2GE2BKAJfF0RGpEsjsV+4eVzh2Tb+s
lv1ZuLoyB6ifFdCckGyIeXevNNCdt1I8kI+AKnom989+ceTqyCP3msu/gjd4idg0DA5P+5pRWfgG
2dwcAcwSeRHUtgkI5iYgWqUNW7i/OY0nRoCYS8oPkLx8IcHHSkCLT8XPnOGTMkJqXPDyOHEOJAL5
2y3Z34+oqHXj5UNXtebI4g97Xr+8tuoWqNtNR48UU7mbv2W7KpHtGz1VVvNCYcIrGKuJEmzkAt8L
HW4g9nx/gQuM988I4TOuC7q6NMmQ9XlVlLVmivfpAICrKcI4NO+uLsyt9fgTVpAbDULXFPVauxVE
bPgbmMMdMPUMZ38YDFG5vI8Vl/3JfvzCE9Rz3qVErZ9cd3kBL/yccuc7XASbSJ60wFQi22aEJSH/
67K1hilZ084B0yCjjvxnwLKR3H4vVBnxi4nm8jg/3PQNDRnk+S8MYn72IOERkVLsAClpysJMQlmq
J51OJNsKNZ/eBqiYRoveMz4zWGMxCZBAnvG1CbAY8Xg1Abq+FkPJXv4/R29ECgpZTTtvlicpyFhp
Qq/h4ee2YV3vXasunxqoTfcWXdL5bg8C8+fjuDKHGJH1n9KiJ7GqafYYhFypbhmCwbxDsFt0p4DB
VdGzJSCfn8P0ZlJsFC74MdW5CQRstXVnNnSzJ6MkvGxHjsIqpku02TeSebG34OVetNOzj5aLLWgs
6Ka7J95QPD/xC4xwIcFOmVVT02iyyT+6hpT/t7guj78aApPDURYydX0FnnfwJAvnbYfHDWyqj8tP
S1d/HOJ9v5SVFF2NRonDCcsx8iI5xylyOImYtVWkd+FjHo+QZ5GKK77r0vOIe8dManfmylH8OX/B
n5IUuU7laWtH3/q+4EaetBPgbxKa2s0RJGIZhzHiYe8HfrD6eZ3b1nc8Me5AJ1NJtJOUC3KcyYSA
tK76/+5Q/7nBAS1anjayESxjvk1u3RppuLGg5FtAgd8uRn+sptLL9YC1j7NMOMIPNBM7QORTo7nv
ms2igophc9NIAtdHK4jzpR3QQZwxfJZPlykKInYgXX2vpi27pTHCl1K3cie/zk8UG/U+0oJzUqUs
erN0VGAttNrw8pWyN01ZspuBFSUsIKvcXjp4GOlFLtLSgdJIsPeFWeoQjSd+DmcaGVhNXjO3g487
msf2DhnADr8aZJN4LPFDgVl/NuVMnm7F2hOhAIGFGTcmruBdhemiHjQaSWZu6A2f/QfQp+BtVkFk
9PvDm/sj4PG9Iakb9CiHnJnwEB/FCofotIVLwn1xVfKxFvq7l9qKSPB/cSF+vCDB/xy2l4FOGvLm
Xd20V0ZqFelRAbKRZE+10KHvG4dtwcxn3QyHCbsejLp2eitpppTZm4kc9GME9BscXVgm5aKXYjht
K3Ojlik7p1/JVkKqfQy4VeWwvfLJ4KxAGXBk5uxAOmYANaeR5ayA4y5Apz4XpBfcdqLIX59bSVXS
dGhjiwJbKvnwQDK5X1umNhzbgzbHV+FsZJQQGwqsw3nyzdJFT0kZfWvCtxAqaTyOuaE0MKa2cngP
e4Tc43+GEVKEamToHDCbDHsSoTNRhgnRaR5wwaIx6tt1L3E8KiJiH798FDzv+QnfznnIHwhPl0qs
iBiKMNwZRNCVNf502TGal4jOWfU7TKDmDtyQrTB42gVXVa/jYkBVaQJv+vBagUrOTqgfVUzzs9fS
tJdnA6GK6l16SZGfZD6CXUnz5x3bNsUz7sIc12598P3BV8/9mgn/vcURH232v9ZPiUU3lFrqmWv/
ALvGeeWeoRZlnhy/y+qEBTeFYH66MoGXl+A5t/QH6x6MwFeCzAfhR2/rHJP3lwaIDimInpowMGYt
HFaAGRL6LqvuWggzwee6R8A2h0yGrYQgTaohKsxatPbX1bRdDVUQNR2aHqGP/HPepDRolN+9dW5F
eYgOin9sKbSxtgqOYa4Eu8hfrhU8loUP4agBw8+ScHzHwAw54ntWZKnSrnO/0hPbED3OXiVZ0i7V
yEBX8Ae896TqchJUCF0XoDA70eP4yIoSgWn3Brm81C7kUrE4Dhk3+m539RzFLM40w4L95Zl0DoK6
LJHMGpFykWeZdnX/lAodSAx4RdCsnP9IM8hYyD4oC0dfzSG2d7AsmWejy8y0EwJ8yA5cVWc5TEWA
p0Pkqvk2h7+8rGH5ALSu7O8gkOljpq6YXuHxKpJQsM+a57SskBxFegPlyKSxL6ARfFCuM1XFavp8
Yzloc7DKTIF5NUD9TL/ZpSlZ4Jnn9St7lNX9rSTlXwIhcAY6+uL8MkGEjLlCBeWhnQ5vJHHjzKrS
sWLEzSjTVOIB9PaPwB0LCF9ZcZue4LRKGxfXaFwIduLuF8P3MtB+5/4RgOTjLhjExjRokhCQGXi8
N8Dnz9reTbeGgUxkdi/JKS33cGMq5Y3KaqG3rHfOBrPI7QKVTvupSVxrm2AxBmr/6Bf3lQIyVgFY
MUGMePJotglQnw4njFcq2NJAgmyuQrYJeVADv3SarU5GnvMGmp1aFTp8o1oA/gcoWPPHiEgjIsdk
9SXU12iHiErRpylC428CAf4TAwIoTt81+VX1SO2v8OURxzVLKdUfBhUmJZ2e73dievirXUEmuh6v
+2kCA2DNmFgkJhrd5LM0o/9ndqm3smV/pM9e+CaUYURFbtXdZme3bdP2KwygMueb0OLqAB4d9H9j
7AJ9iwRU3zitDFwlHAlf4TxrxiPQMV0/4z+fNPVMhOhDw7eW9Dc7elhU1tVAwUIaE1L2PqcG6X0o
MPazIgz3fa5HOWqI/KMsnC+3sp3+rmzpxYmjdEu2iKyWolPwb9vQzxqalytmAGp5ngDZr9C1/hO7
dHSyLDv76+eTTz6BZncjUgdujnGzl4PlCOCGpoLoi8r5wt6rkS2jInDZxQfFYWNRbBIA13Lih7O0
rmrwAXFTiiaywo43b3vz8pDoCh8LPaM2ORcKQen1C0gPHsu6g03mgsA9q2/2c7RBo5h1D5FmOs+a
ybMMlkD+w62h+tZ/PnEyvh7P+7zuNmN+lQldgSsgSDV2GCSgEJX0kRPiMa6UxiqYShXrnC+b1c03
vjSZvuEggaGMOG7AZp+mJ99mKdkJm4MJ3O/UdALrJPVaR5S8t96FOJSgPQTC4b8YCj/Lr3m4iQRe
E6VbS3ihyuYbp8DgYJP9MZaVCBh+2F1gzWTNGUgpUy0O7co230i186JQBXdpgah+WPG+G3broONk
4jdZdq5IcSFGzQtWdo9tRDGfMcwk0pmSlj+Hg7S95+nruoBzxp6rI8pLh90Z1Gzl16U1lB2g0l2z
7ty1JEhEqDCgthsr45Zt3u0jpuFCe7copgiFQ62FAkElNyoV/P6RoSKP8OdgcT/xMVXg7c2rzT30
AHzhW3RQwix5mV03vrVj59Jr2SZIP+acYzw0SpwI+H9A1w57gKx0+/MkDTC4/bMMuR93AtbkvoB2
j1JCDGZduXuM86+YWC7Z0p1I6o9LG0JTGBxJtoIQ0ujwZy+2iPPcI4TLr3NhxffVJnBLRMXCkM8S
T7/IXInsrD08ARUA9WphVqDWHWv6kcJufJ5Cdj/2ZXD6E7VWbeHuC7ZwXAOQpKCtHFn0oGROO7tx
FYgZx2rQi1dSNmhaWwn+Ws4tpJ9dBoFtY8g3l74plMkzjckkIQPNPRerxIVAWa2QZrZtt2YKLpwN
jyxokJrlgix0aLenY/M5tq+8IL+rYzboUCTAD6YluaaciLzxg/LTfJbyuuKowCxO4NOaJb+7SZih
ECqEEXafpT54VVwq2Mjgm9jdlXzZxtFkGlLcIFzCKLJt+61qrnnXEdgwncfJfP4i+3/wnh7acTUs
C2NcUBDOfTV6sw2H+4Uc8RjmToZIh8ocvdJZvqdhEeY9IzL4b/AcinaY9tBG3jT2TCI+NDrfb26M
f55YPmV1VI27dH7P9+bzEi/+bf7W1ZWASAUSg1WDaRHPe1vfRm8kSSNgn4pefgGitONWNfEFg7EA
tU5gtlupnfaML4c7eMbLP7hzroOgF/CAiHdl8tnsi3+zzqZ0zRhT7V2cTnxsgSqkT4IvOmP5kgZz
5CzkaIq1CpTnG5ALF3FonaxvLefyT43p8PGXNCH6f7oGJnhUsjl2q5Goi/J0508IDFSpOC5IqLmT
+84kSza0gmuvjAAfXHiTigw1BSLdrDEkz/SKgnoSg2ms91CsmxKfa3zoq+nijnnog8GAAU13LerQ
DsWuedOyBXi2fl6gNTkIZzGEFTMVKhzPzlqTrzeKC0G0iOwXHde8BHle4c64qBNCv6VDs7g0JSYJ
kWoEzbk0EnoE0eY0QukLxU46sgKXFLFUan5vmD4HsqFoc/cLM8dH4c3dTE/dW8OMccW1c0Rz4IxI
mF156YZPrB3s27xlQUkvbmFqSNRhGrI7mAvp5V34gJN/M/jKB99ij2LV7bNB7usONJuW5+ezSyPG
3qAto6GpxmaPjQJYyjTvCXLB7GC8eOXlaI8a/0KW67C7ioEoeqjpUasUoJoih1LYh87y1319n6hn
sL2+IWgLKaz4d3Inq8QTuJ4fCPOuxh28YppBv2vo0WC9SdISyZKJH7zeDdFAQFPc7Q8sCAO1aNv/
iaCmu4Bzr3aNz82hGs5v3LjXTCFjK2flGJzKpW83Xpya478cwXJBrdZAckFJMiRndlNSdw4j9uE/
dwH5O/+Dx/PgkNK+rpRdppDBOWbsOOn1T4g/qccy4Epb4kFZp3UF1AQm2it3fOY0iQkgC29aHnn5
G2/zeLAvRRjg6VDoxsOra+3IUfkRWvsMPxiUQfcTUFtM3eJgl43TToW2X3aLGQm0FJv0YdHw13Mu
FKvoxbZN+u4wXSgIg4+Pzn5zS89tNrX3vRelf1xLOLJml2RBKM7nE33BRSKS3D4QnTIFMNGASm2d
mQp4fu6adJpYWxnjYLEhNBJlCaHtELGyRWpFpVdjBalx60Frbehn8vrjsnr4EeqAWbf4ZnHRBXMI
tPjlHeJwMdK+ktwTW0P4G6HgtvA9yxL2RlOZD5uzER7M3vlLu+QlUhA5wuU70WZsYIrrcTsC030P
86t4PAgIxQsLOPZMgtH5gyEaW7Fe+ZizJyeIM1+BSQjc1/3+W8dFNtxX/d0ai3saMVUh+FhfMz1r
e6NBJEkbILozXOka5fmCa9tw9RIvj0wTHnK4cOXveLlPGMzg5yjd0dTERA5hwyDZY6Dv4z3jRGQM
7jlYPJXKVJ9AM9n64nMZM/MV42wHlo2PdPhBIpsQ//K5Pvkm9/F+0du1EIJdN+9FeCooIMNLXIF9
368AfklSbfR6UJT0G35izM6x1TMINoqiuqySd52zSjO3JomoRKpv227RZG2BO4Je5tPqm5fXP8zS
mwt33jsQ7Rr1k/gKWp0MRgfiDkQ789tYDRZiS66SIXQbl+E3bd20fNJL28f/hsU1BNbIBcuOrpsk
2qaRA68qRGpEUpokI30onoYsZkoIjy3zQ8fq6mV9cM8C3wg2O39ty4bIitaPaiPsQg1UT5o2iZKH
UP+5ONeYo05+fbvjCJULuyXXN8oRIqA7VoWgwImYcHnGDv6OvjZzpj1+Ho0VI/85ADwMuUe69P73
2qmx9a6mx12lernhttsopvj0bsjvsClSCAUSY5e3+m43aGz4gbI530QfA//wBuKWjRZzifRquYg6
YEVnRavGypzBO5MtkX2kEpG4DDI4tTfTqj/lki8rlGgNc1A6lNTUEuSo8mOj3tWgTs2jKepGzKsx
YxT9ZpAYNMSWhDh8I3hqKdXze4EBzpWQKI9iKq5t6HdkRgLepBGR8DyIkWUOqYiC087P5LE2r352
bFqURdN3BU6dGY3Z2bmwkw3SiH9p+zSMiCxX2QEYpOMaYnoK4+bAaGtb7+v4exFnNvdi50TUb9W4
cF9mOQ9or/c6fmER3HHeJvtjMXCcAAWTq0JpDa/NWx1nMi8H/fVz+C0tsIeWuAzlRl+AE5FRvpaE
wyxY4rJBN2uoDFsdk+LJC1ilKjNvDSMHgYOIMAW5GV5jV2VIndwACJIC0pSA2F93OrGpm53cUaLd
EADN+VY6aNCZQUz7z2sC3AV14kk1vuBD4Iz3xRtgcFBeIUvUQxIFPuI/6dRVHg9U/XkTaEQw/URW
+HnfBw7EUFnWpLktfCMZ00XYtSJq0Qa4r0OdL2B6ZGS1UY9hLU+HqbPVh/Z0NKioIfe3OUIUbxoy
VEuv61fF3CYTEAy/Av4BINo6TshkRanK221hljNpN1LIQmN0Wv2NrnLinrV6CMzdZm6MsdVPlZNx
yLUfCelAmpcWQI7NThMlI6kc6u8HcEIYmbUYKVtw9+woij6b9/G0hxBLTC9kF1GmEGwr7ITP88Lj
F0hRyvM+0lUsj2V9Zl5Kn9b9tpe5V2z0bcSW86hh+pv0whFaxzhx9qzWvtFz0z8cub+Gjw9qcmJq
O1nwL0097WyRjZtl9dkU4T4J5vXbSYb/4aYaOi9ImpvKjRITLlZjGgwhNT65HZNsxxlrLHXIxyla
pMf3/s8LslLb2mHNTdPUKL3EeD/4kgakw+LUArRWlmKvFRWPbo5TmqhNBLEItPv5jQ6Lc6dgQCOg
jRiSCzWrOTRylb0e97TOog9fwREqxLBVqzB8cAnOr7UUuGtjO9xYUaQDzr0aqFRBBRbmIJGpTADf
PXRGy1hmk+XOd73IWQL7kRG+Jb2w0/SLbYTy179xnFQJCrbu8hZZJ1lVLMBKu+uZ3uEAP27WECuB
x7q8N3E1A2bOfDbDiQNemtVDtoqlKolKcYujTIxGtJNxCnfUtaGG9mo7N4Psb4CpFetkj/v3sxgd
BuBgCHR40whxu8YwjkJ9mIK1kyJnrbU/oSZLAdSB27khdymmalVxM+NMtpR/X8Fz3jv6UO0PWIkC
JurucAWf4htlpECBmyndY+szg3HUNnWI33YfR+QC8xYsR3yDFBBhxpj1FmkiBlMCLT8Iozj6/1B3
X3IShUByBJX3XbKY3eJqe0yqCSdqcjN3/FQZ8PvYV9N4NX43GSF3o7THl0Or7q4TbP1ErVcONE0t
4eDiXHdyRp1z1eMTvSLa18L1ZmAoZ+Z2MfhnsHsauvcEAbtNZY4WEfaoYeKUmlbMwKgeL1W2DF/x
Omgh61bu9VNhrcOySXILzJlDcqs8qAO3aup+NbTIDl1cDSPfMvvF5Ls72JBulPkl376nHR1FuDZL
TZR/qzYasP8D4m7wEotfKljf6mXM8sWPTfWCcQzhrOrSgv3JBKFzuBu/d5zlYZCr9JP0GBAobqbg
pyv6far1TGWTdRIwh3RJa0tvYDClk93EoUMewDtQKGuDVb59KjewzpykY/eIurSuBB7dU12ASIhU
i8lR+Ol/OaP7B8xzG3NMl7oa9FQCjwkqg07KOk7o64B/UA//4a/iYzOz0Jbvbxsa1MM61J2j+Pxp
AYrberyzwxyE7jMeg8EGB7fmWsgnc907IJl8H/DJP5xjqZhixrM3iFmrRkrlONMQ20CsSi6z6RDG
bRWmHc3qe1x2XYM5YsLsiB+a7lEHvK9Vv4co0CblEZUZhOoPOT7DzvGaEBW6p3clIrEi8ZPVbxGQ
rOcjPo7Bk+nZhDQyj6IndacY6FDikE/jMIZS9FVdsQxPwTH/qTNyorsPNN2tCzb5DTN9Aug/h5Oo
ehTFJkagNFqzF9zR4qiOYVuj4swsiyZSi45RNapngIAJ8o/hUgWohAyCWmgxZNCpgOkocf0zTfNx
3hl/AvbHK5Fk/QDwHtXR8haO0uIDeBad+sjElhbNXrOfkwxQEKuyPzbWp3dPlrLRxQOt/9dURAaF
Am2zghEYR5mhArj1OKBrZVcWcPzb/A8QOXawV2lSJjXAWZka1oEqgISUYD9Y5ey9aEVCYecjtVr+
OtLVjFIDmVFjy63bIBE/u4I7gZrZeP7xd4muUJnpAcrFu6A+Feu2lOrH3Rgm8L+KWqPgySa9wLqm
YHcFrqNU1ZFucoVoThlc4jfJx0iVBD5BhoEGFr2/4/XnlMyso9uY2hfEidOPf89dj4tWO04DdHgO
DkIlEK6NTf3T96gK7Gb6+6kJGpm2nPO4SqCLKPtAcpLwtyUMfbDDfbLHMU4MaSfzbayPNXE26gXP
y+tKwpJq0U7xBSQK31NagQ+kkqaayPtmgomsjrgv2ekanlzp51BvndyUjMiXQqiDx7mqdx/ZtGmj
I/u5lWT2tSYjCW4jqfcNAho62NUC668wI8fXeAv/kxeKzTeSnymVroF7UzlA+H4JlOfUK1vta9c8
Yo3jbepm8rrWLqLd9Xco56RFxaqH1oNItaXlzJYWpixpmNUzrH5EYDo+4sRZVeRJDqLy70p03Gt4
lRoxdjGjYwF4q+quF22aVESue2S6TQ6fLLmrUNL7dnRjhAalxaA8GgXv9uQhYCihzZwp071KgJZN
57+4+wyfoVJohC8+Ct6BrA3oFhKnrx9xLBPwJ4k6utJSQvEjxm3stkzxum3RucEVsV+LeZ9R1z6B
My5v4mSLRYUHAQ7MArkaWaum/gPGKpaagO2tVHYg9LKV//vPRi9nuHhr72L0bj/oHOR08+IF8nf6
D4Mf98kHA1bWZC2O0kaaSynkUr8u1qEHZaRUNwTjYQHwFYB0WQSGdzAq6WWl8du0Gphjj8Rt/Vl4
GPS3LpgtA4z5AvpYVgrBT4fpr3NQm+kgttAT6BQJf1tQfDorb0HcVpbie9q8E+tcwaipTuYHFdqd
zBl9UrAMFW+AFOMLuYsJ+KtYJgyHsga3ThKsTN8P8Ml7xTTgzMTi01ldkRHXamInjg9qW0uLzYXm
wv66Ukz5IQ7jxqAhqyx4PVwv6ajIYNVSs0VzDz+EZP99ivXE70/qnbQDArB5lu/UqxU+ni9udMsh
BbjbNLHWLjwelMKEOACfZOHkbi6mBAGAnA/XVkAyctfiOhe5SJbUsIm+9bH2wn2YVhMLvVPtiq05
5T8ywUEUrbKfl7kUcUF7yCfDru+6wrawtJDfpzqdvk9LC/eqhb1glzKG02rHE6MZD1ENR7u6Y8Po
g1vZSv31mDrhE7BGctaBIp/E9tZ0eNmC/HFoNwudMaAKnWhnNfYFwFfGuTOBSqnt2cs6K/NLsXFf
G5F59pekyCP0+aFjrtQuow83pihQrvVfl7hnA6eFZpxE5sMmWr6sp2Wp/LVk9T5XIs1UdY/0VfTT
uOLBbTrjC9/GiSHC0AKGq6JoY0sRNzc6yjXiCLoB/+d0eWFuv1PuH92EkdMpoBHEQiv/VZLd/v4B
vWJyX6Ld+21EQcfSO4WwwYDPXKBuQJZFnHgYewCU6av3V347YGCx7bBhS68Eb/gr46kGdFEbSmPk
bW4BmvZdtfdNG1Bno3svx1cKlAtcmlYU4+yFJqwv66Yfx48Jd3nKUD1yvb8G/4b3Fxy5/QSx6dWH
TV4NRNmf/TYnnm9mAQyiqyBxrhR29URUnUuWU6Ok4HZtlgYYjwQNXHnwD8drPH9O6T2rrC53Vi+H
FbEK9ElkBrCI1NiOvaJm7QSarOMHXKHyMXSQ/do1i2Ego6SARMF6bKqeEJ1ZYcB4CmyOXStWsiKx
sC5RAiwV8cjYUzDsCCDAH7J4+SmxNP5ttfF56V32hJAMEUvOVgpXkmcreIcm/UTlRMOlAh5DkkVj
J6aqRwYKNg8S4B4v2p57rkolP9Ha4JT9IQ0RSbXqYMIHxNsaxilKzfiuciB3epCKZWMB8z9CIBxz
0AVdojzcN0Qa0kcpHIJ7l/5Aq5PHmC33Q74HUs3a4ZFwCV5oGv0Ok8iAeWmYsQYQepx5BWWOciHn
35mk9xL7AUBLn36RHFltMYYzUKegsXJ9GpWEgJqJ5irHKLYs+Ps+gJ/lrxoQXKiLGLZTq7qAFAYW
mGZWzzNifyqv7adIG++I/2sgkCA2bAd6LkvLSsAZEh8sbGKgngPO/LC5mkPotmDm2UwOJ3O9FIz9
D9nASP5r69LypcJWBsCP/KzFRXs3CqHHycSq3jQk1Bh5pClYKxaRtwmpV0sxQaA1dbBVLPUGKJOh
gxpEQcmyF1m7MpzuPOXtG5hYn49rKCcB6iDmuv+iGv458k5kTMUWWuRLbvNso5gtYuYIyZvEZB7U
byxbZdPOlij36FPSYwxUwCK7brraataHLc6UzGiX77TgbjyfLG57Flh6YULzvTWHSLMVx0FFrRMj
ASOJ+jzGFPlejdEoCWMvuxh+U9U6Tox3hQWvgKvfzl7iBKs8LzNTJqTsFTz3hgs8dreg1P4O8ir2
Ea6G3frsH2DDnz2M6WimWiUD5yHyS525RWW+9dvAlJAJNVlnCOrdRNocNwfp7LIRyxDMyLBUl37C
1MMZ7yWmS6sBv0qb49rSXRO8Ic/C55MfJZ3B8o+H3hMV68XKM6rRGb+QmlAgZ+wOjaaUVcUAVA1N
GSEl06vLZXtjxisX5FppPFSc6ytASMgwwWvWxFb0+oB3bNct4tP8tjL+WfF557fq1CHza3LDzrZJ
AelDy/Y5X4zImPnmnwvNFZwCv+ke4frz2TuJZ0S3qGVyS9kpFR+oBgDbTiPLVFW+iDAEnmXNFKD5
TwgpJLe1PMAv+9UocZyzX1e2UiGxgllje84+5esej/Nq9c8vdZ9YXkDeK8fjO/p+XHQAUI0XILAO
LAPB/v6t3HdexRHLvPxZEhEr1HJDNHptkj+OUmdxRwjFWcWne1zGYM82iLBjGF4lzd3qDv4nQbiH
Q7mifziJzVAt3DV1d2tC/1yH//UuDy1HqXqDCJpHEOArWYDPFEIIttw2wQui1lJtVD5wkVSf3i9I
aa24mkqpFbK9+M/uHbeAC9eDrtnWjgSYcszSwmwvHwi4DSDNf6zFblBR2Am58dh/u7G2AdMyI4VL
arVi/qQYW9/t2vq7a4qhIQ6BzVX8REJMZBlI4tw/KLqwhQq/1w78ZCsiacjEvbBHT2SIw5c3VkHQ
S+j4DC3vSgHjQNjcZ1qKBvhUOKj6uKDKZ+3HqtBDrAg+HgGQu/hxO6FvilO3j3wU7GaevuYimWpM
9zG1EFr+oJO8CHnKvRBG8B/n1N13i9Xct3FUYMoOhzcml28MgGBfeZgPBlqJuq44YmdY5aR4L5X9
tWiMxePstbHQt+7gixD0DOlWTshanSZSjRHaS1PQFCHbdan7ZrvhzdesRDm+LWg7LRfcnVybZr2m
3eWEyqWA0itfI9VARQtIDy32LYK32o04co5GW/WkNKulr4x41osxkOA4/CWs3vQJwg9lRk2hRVfx
1CVTHHDRlnldMeBK2hsyGD2RRX54AqtM7wsheF37CFygo6a4CaGTPW1bq9BX9qkg8PNIzBHyOG4D
bNf1tOD9xu7Z6T4+4nzop6uV0XvUwJfH/pirrCO2nDu/YwgXQk2Yy9B92fspiFWV1Ot+ShpzkbJt
2ziP6hZHM1O3BWgga7QI3G0gCboYkuqNaRsMtoopzVTlIuiPmTBC7b7mn9hzI/96Ifg/C97yh/9s
2OefMKddA9pZo4WV+n8RDMdNi0itl2JC2t+y3XYcIUa2fF0bNU/BiTak3y2j8XkVu8VOt8haWo0J
/wLNh529KQh34h18OOs6C2KONteT5eY5It9zzdQ4noHvDNUNSA4ICXMg1zu7pd2JQlnED17SklxS
v0t9/6qC8KiPz8dz6XS3ZsZKTjKbrxTrTZDIPg2+qm+kUyrLxh7Ekyg3Pk7YbY7W1zSBC2axGqqV
onZh+eL0i8yLMzzY3E4DzbHnACr4IJsgkp5m6VRy8mkIz1qISj94XM7QvsozMuNz/xZ+9AGaJt6c
t4nBnJ1HOxyP6sPZQNtbM4eRxmipzm/uhJ9cMdANCN9ZVddgJSSc7oVFr2vGL/77cUa8s4OuWUZ1
HxIvFhCJ2Gquxucy2Hk2eN8fe9q0lD8VaWeQ5JWEhelJhuZSjK1lrRo5YW8M9U93ya3ZHJ/kZvbH
m9dxlnwZ02/AbbmutKlKk3Fqns1QHL/LGJwY36KBjLPC4jKJpOz83ausu48jJ/IkuQYLE4Xn3ELX
srL4Rg7N0xIo0Qo60f7efQXI3bOfC6OwZGB3F8XxtkvCg5iL5IOC4cE8Pmfe6uBTnF8wVxCJFAfI
tLTOLWntPi4kWX5lD2DgszD3FxjgSaI6D6XpnusLsCzboP6V+trst1rftin4Z9feu9Ot2dwdu+yw
l34u+kTwVLCmTgUnhVSKIBE33dmFvqJbF7hsyZmT0QTdAtkc4Gddh9SoqjGvNodlK5g4p8cINnfO
sdQvVQWzeuBoqx+84hqS8Sem3fm/GYwT6ed8M7AEyG32E+AGtthW8WEO6b6I54qu9hfEtOEVh7BK
8xhHty2plOOnsSMmq7tNMexR4J3Tr/e+SVV49BKIMbtUp//n+FECfdzN0Z56eMKm+Lh7G+FCPASk
e3go0/UsNL3PL6WC63/fB8WD76f8Yh+wWRP/5z0WKsIWttqeasi6q7OVHgkhuNW6nd4XbW2tegPd
srJ6v0XyfTBd3qvnQZcMSmSJnoLeCkt99EJFFy6CVaRQ0pZlSDW7tjNVyC3OfBm0ptdcyPd2dc6z
F6xwSELMEcu7a2LU+h8p+Ar5M/isagk8K64g4JhPNZdSD6QDGrbIwJgcnzy1qcbw/T/Ae20+fvFF
ElwsYWiOirnek2docjce8rxtzcVRqk2iSJcz2ZI+yC8Zd3g1I5KoJNhedwf2AkXYOc0rIovxZ3ly
lgMSPAB65ReH2QzfnwKgOUKTWfaPmduocR0zf/KGODphgvzByFiZqLudx/lYk+DT/FzP46qRcakX
/jTOhjMYtGw+xPzIKDa21TqGuBz0vh8Rp+9q5f624a3hW+HXJt1tqRHXFhnv7/fAbx6q9AOtBtHQ
LViF2+qmQRtGtn5X7bBAVqzdxlj0I03e2vnPcpIHDi6v5cZ2JdzVnbmsIw8LJiraBRygR3b4K6lj
G1fPeo8yrt3fNgb0MjiJ7t9JWQyHDfpfcIhA/3GhortS0NvkN5lqLlqY3txm7Tb9qDg3fyM0AqEy
1p78JQZzyeyPCbUlDRyC42YPWY/eUp2tVdG4K+1N0xzM/OK+eEjvw2MRVdzigZZV2U3meIo/5UEm
/WoHOJkmZP/4H70H5Xk4l4P4CsA1C/UuPC9s4uZHgNQaggE7/64Qx/Eg8Iun/yJoh4v6BdAp03AX
+faKQO0GVTCapB76VYL62Zp4fN07GqEJxo5K22gJxwgn+GR5BVTgVn+wMaM7P2KC+skzVCP2syve
yr174WHJU36gWx30/7eX2y0rGyCmKMnALE8WwoY/NARyOjMGnxkAuiStTIeNR8Ucz8nXFIEVeRpc
6kYbBXSyfw70sQCmkEIMIsHcWeAOJPOHdhWXp1KUzdoNw1WYWTit1PPP+AA71IN8z0dSyJIMbAAp
369NGjLS25uy6PALU98t8xxe1xgdXEZlFY0Y683FRe+Jp2BPWNuK/KURwpSFnVYl+W0wogqLUB5r
HqEWCC+TMgMfQLijvv06abmpTnFa1VkPuOjGxN5eE6z+R/rcVt2z7aim4EQI68TlpoKu8SvXDLwR
KDL6xcQ+eqESS2gGLBtTYjADiySrKMuo3ZKe2TszVUTiQWSON/kn7Uso+8hHdiG5dxiOM2MIoZzI
Sb1ruuP2leW6VxJkmUIXoITkhoTOv9ZQCTyAUHwKWYyCiRjceuHpBzBZxfrteYs7hh1Did3pZ+WK
QJD9YqvpKoiNs1hzlwn/j4fi2FWOaANzBiWi9jwRCZn/c+8heRkukkl7+5wm5JtHXfcnjlIhbmSK
RX+rYDM81RoY1y0baC8kQlxb7IQb4hCrQXrRoclKEEw74WP+UzeYIqroNUDbfW57LwFaL0Y2wV8Z
wormmSjtBgKhJiW0f9NxRsNul8tBimOkb2DFbeVqCC5WHFXv8bCvA/l2kPw2DvsYa2mP9cfDwsgF
5Q3BKcH9qdRZ4Ri0qj+uB+wcwb/zbhr+5c5TJv6m4Dzjn1jiJqWbHSzY9Kj+TvxYQNvlEX1Yv7DF
4JThxhDgaZ/gMNzfvdPfvR2gfrzkpdFJD+6dN7GXfY271aW87HIcuL+MzOgpGduIiUQwFNcN1HBC
87LtPC8slTgJYNnIgI/5g3UL94Cc4z4I30MYFriwgiDUTcw4XzYchJHfgPS7maZ6Cc5/WVY3eAYu
BCJD6OM/svEw7NVcW4NfcwAIZXHHZs0XsPwV3Ue1kzzScKEGpTWzsxzFE1OE0v/klvBAjSGtOMPk
lLniGrWF7u9/xCGMXy8HyL0bQUZe4F8JmmXrdRGGZW4efjOc4iYLEhSx3TvYZSS2Kqgd5ODainM0
oSmYJk8YgQzatMf2QSUCa1X+SplFr8eEYcyd9MNzEv1OL3gEjdTWcP0nb9bnnWWSEjZ/ifMXhASM
Qs56Wu94KSe0y1qtuM905QeuKORqJs6/mZxKKVmAouUiyMyj1F03E0fJe3ol2yYklJ02kRh9hjmD
pQdGCxEtuBTRX5uRJmXtjlbGNTyDhSQJ2fUa87QGMCpY+Xl9I9BOrqWkYlTzVegK3A5uontb+UdG
FlgzbYZvOtuOauwVDXu1EFe7mVSHCDE5LYimk3HUSsKw6Av+9KLmnrFryiuvyhRpdDLkqBbgfCuW
ZE11mP6/AwcjLvB0kMuMwV0dM2EkpiznDh3Jg5eVU9XAXO+3N76Cr1BNcvrEBqKzZn7IaMbqjOcU
HjOIyeJ0VDuQEW7PY1DZYCFTmrQM9LfArmYGBPRY7lK9k5pslbx/EcQaYW7xL23i9DOTi/mYVEIr
Q/1Pvfqjuj2a7v2t/ddJaxkHRq9qbASiK9p83INq1HRpsoNQTvWG86sPvCi+Vti3tO1nL0vwSdeh
le/jghKIYSFuWe/Bxwsi0QCURgLzhHeNCtgvmlcQi1FEIOkJYZaIfqKImImkJh32BhoIPPugAGAy
m7Yg3jAElHrm5mhdDuQJIHdYhYX4PoIodyEKUgfMoj+Ng2v6uPDBI9IA6MgiLfOLdLeB/kDWJfGp
1QG2cf48NXfvdbnP/Njn4uuReKh22L9qwDMmeoiBXu7ihND6rGn9t+JpcJ8I4B1jmJ1PMXw/AyH3
Z6B05uJ4vWASAmC5VuJipAI3lTjv/mDl89sLfy9VEJfj/4yWvTDgTHX9gAzKOLvJdxiSc00i5UZp
wWw2gx3PNwCQEtfBZLEQ28S45qFg4fMACECr49OcDx9k8JErANzf1UZeyxzdciUOza20Bi9OD7R9
1HTDAsboYuuv2YKkERzakEVBjJ1BAskH8xG36uygedFB3SWOB2pmnEq8EGjm0VenErgJqzbVNlm9
5fBySvIWxNepZCBcKjpBbmjxGvuXXA6VesoKTNSLYRusbU9UnDbP75JJaFRy9rQzj3zpV48jFfLP
Yt15+VtNDzGL36HvEJ6qXSrKW0XD8xl8BHfyIMN60oR9OqNtFUatV+SJdeKgzrVpv7n++wWgg99w
7AUq/Tn9zTdLZWJYPc4ITZmoYC14xDjIXWbYpsjALJZIol7GyHygWJuVhtCMu3LKFnDJHtxVknRI
/UvC1AnV0qBrh1ZSsHZJcDUN9xDcxsfr+KvQ8JIXAu0T909DA6bxq9DJN0ycPoXJ/qhUMStwTfl2
P+sZr2+JF0AatwMFQZ6Yk/YBUyZFNyK0Uaide2k30hWmp0Qo8v4ULqfhXIoJVpMnhGOT+WrBgXeC
4GtWy5rsRdm1asTdwKE9optO2XMlBHoDiY6U3M+wY12FkAueXQjzDIFa3mKPG7I9ir0WcRjSZC7M
KKnbDK4lk3xuAjJ3hfwdjdONKKjdGM0RGuFMQsf912AOHwc5bTlXDpCi6ZwWy5PSpmBdkHPi7D0N
WnX/Ql1FHBhKjAoFgzi6NNOjQ1l0Eucqj5G9VH/8CLIdhtlckIHgx62eg991cTnOkJoNtnHIDBes
V1GhJFD9xZ89EkF29zzB/RcU51hltTTVfhFonYBNT0vo2Xh6jug6SqSzq8W4sBBcUZk9GVlldxTy
CAoZSuWuUd7Lxip9aOkr0JSnbny4yIjjr6pfNojashhg4eDh2rCwLAOwER258auAWcw7al+7yjww
kaVG7Zue1jNZCJZZpJEa++IJ4mBj2qLeT+EwqqQ190+p+NSloap7wB1Q0U/6Y8/suvnCX51lx1Pt
oiteZlwIWhD6bTw8KRyhPFgHVZtx+/vytaWEPWDt5eEZVuexVrPFzx5055dnGqvsmaEql/15cljM
+Zyr4RUblVJl4JcB45x0qo3DeIfUFhixmEqi7ZRg3Z6T/Ayj0v+wxabZVDuT9i4v1YprfYVmInDT
U9sfS9N2lONWmerAVxpMcoLPokWVIOPt9e6Rvu4BUBQUqXZ5eds038CoIuUlEcp9RyWSxqf/8l7R
UpVztqv7neRY0nsFLG/ZdE11UixTjMIPdPBFJ1td6I9Vz6ZC3SvebqywDRg5M4hJ0G6AHYCgke+3
Y5TTMigt4eyJqZiJcz1cDnUJ/MHTwVirk+cImAlac7za9z8iPVBPp/Iofn1oMWPIFHiBRI+haOfT
IsDmuMwGG18NyT/WnRQsyi7HuLn8nSUdAXAtHGetOKKjCQI9IrRjH2XpzquYwLuzIaFs9ztvgRWe
ihXXalQ/p6CK82hUQV5i3vxkvTXP7EVDc5vwf/9lvkEr1VdYpxg35ANNqgBbgA0EgNCegTRlKiT2
66nGFuksqex2Tv3N71VhduDrwwQcujnqL8YQd/2WACyj4AZnAWuHBEiy2T90kziAvOrTnFzrL+JJ
U2q2HKhQusZYvNYfg2Nml7HrtqHiCLAikSayCkdELGI0mM4UMhKspnIl79HkHgjLcIc060p1yXLv
w4wdMBMD7e66JL4s3cXoZ0EtsMGYhc1K9Veu/EJMBtf3PKVT/sPLF5TfMR7rtn38AU4XwjHwZYAu
GUZr97b/ftBg90C1bhKtrCKwvAYVO70KioFzCXpq9Pp1Hsh/MabwJU7tJaIve2F8sk+xjzinI+O0
iYRpj3plBdHwm443jNLnzcPlvmWVCRPOxNqh3YdNqR6RFJk+lFsD9ozFpJAmGlKGEmow5wuN5U3e
giD3bRBkNMKuwCpjEWKNipHWnY0zTAQuIht++73f9tFkr71XXpScYEuzjNTcxeKYniCrG3O+ZWNL
CWPCbcmkElMwoGumbs3smfRmT4qYegkAAWopTQx7G87JWaPlM0OUaP2MCl6Uv1gT0H8uKzTi9sdR
4rHefGrFuaR/Y9bWfRsMkbvGFeFFgHQLRmUGUiU8FLjcLEqH/AKtdnmhVlq9NUHQozVsKJAFcc9u
YviNiZYte7Zo7366fAleqmNkTEEnRSC9AtbqvedqYBL3BMnnC+4y6o+EHMhfEst0bVWnRGAGfxNQ
mMpgv/7H0hMc+uFmaVH1B1+C3W24AaZFRgWoalW+BgVqx/9PjRPtejb9oprzeGm3rKdgE40/PB+a
BTC1fwHn8LV+Eygzm9E1L9smMULZh0LFS2VrtLN4OgQDos+gbkQi9+4VCfDfHao7VsgcIGdQ+qr+
ljkpFi4mOAqoC2e4lyL/jD9DRd5aIyvUrWkJ+jObOyLsE3r4HVaumtCTRH3SWwlRKuezOvHteV22
+XnFwtnAXQOFkfa+d5544Cutm7nrOexWkiSNBdFEczLtxDlEyQQIfxsRrDIiQ13rCe3FqliwQUf4
PG4SvABdb/QmJXB8DK8QLRLSGSp1DBlTI+fFWLySLefqYe8xvudRuSPyFSw3N5mJ/KGOxWjONs6c
L4AgDNPAnU6pj7MFX6s3B2MmA2Fo54yvPdiqwXnOKLc3tz6BVSGgTfD4ZEauiZxRmeqWREzmbIW4
MhvM+CG9lOIxO2VSSRVq+RFQijxBYMI5ojNjwoRKjRG09aSU+GANDPW2mIHK2VoSyEQlJ9m0UTLO
2YmK3BrY33IwOqIjsdrMoTt1JpJCzsf3sJpzUTft+TXys+VVCJR6Xdz6AckT9plQtKlBwTTK63YV
/MZJstlZTARnO+tgoYEZpRJDPDjzNGQ74Sp3sN80zF2vDKXvSHaAR/vw2vhdH3hGTF1JBpj2wkbu
QB658nWY+trE8nTQwE+mDUVwSuhFcKD199kzTdGYPSKFTiPAhWsXyk6NCWKfSFz4SDeOycgGnPZ6
DQ7FR38QunBs0wP8AG+tQyn/tT1aRK/rWCOtlKvKmM7t8FmdO1RnB4zZ1i2pjSuRMMkfGtExpIXW
jRfijjy04aO/i3OJPYzlyPvw/5EbULynkBgjqsGEvBCnl9n4N3rODqzxKWwKvixrvxZ8UMhf9G6Y
omjH/o1anKihdNhyF5vzimk/LqpQP0Ktx3AxpWbrv8O+hfHpr1oknEp8X9Xo4dyXby7UBksheyQJ
fWm6qAl27aR5YbFYWY4i1wh0QxNkPH/VKPSQ7nichUR0JV+NM6jjH9NX2weB2LChogA8wABpdhQH
78+SyTeEAIcezXAOtAxFCWaMkqnb+NiASlYStmyU+u5YsZFHLRU+TJGNtBPoDCxFGa+oC9yfDzdx
ZYz53Dq4ub1DyB3q2jopMk3eT6RKSt8bftAaS7RpeweGgV8tGzgYvI+jUjLeuEALgmwHqh3G79Tt
2g4/UdqADV+tiNmcWCaa/Q1UXQGgq86S438GY0dL2bWhiFL/tHLLzXQjeDrbzSt2tBQDYK0+Yp+N
pgALXGV3j0BSMWsm49yMXZKsGSWyBD560LQ/AEkTTJWx83wItapZ/vE+131AQlN7y2+5m4nKwwik
TGHbmCYhYsSlEYHJQBykCeoswHCbEHXiktSc1aOTozHi6/DGUxk4R0QGTapYC1g/a3fhrwNNL+Fc
rIALqoR7lqAqS26MlkIk/nPdTPRw6qnPDiZPUEJMjsSND8d5cWyWVXtPiCovVCZBielb+mFZWJkb
gP6OSo+ZUm73wsyiHPVZkb9fHLjp4xY4kiOVOJ6O7GnVWUG6BZQjCObNnA5065lkZOEfe9Ki0eGj
GOz+ukLqI/SPR/r8vpOjefRXehKXdpklTKWZMjjjpz/Kisaq64yzoSe1cdom7rGFyKktu7s59faQ
CuwINwjECB9SL4Ni2bNFdfzeP+5vTaSfdjiqIAh016MCXi4kh8mhSKlePTLwBW0uf18SiudEvQZ5
K3t1+Lut5SGq5USZ74McSrsDD83oS3fmDfhTD6ubC3juV2dzI51wOb6qRetSTcpIRUrOOkmJ1j4B
zgqQNpxnBt3aYYUOjLRfGaIx//7jDwX234urxdVAqQ67Ry5T9fyOYRKxbICmclF/QTF5wxFmgxg5
BZd8djB++wGLOw32VVhDTqUAz6pECX5z8V9+/R6yfBfYvJPgnY8aVYBNGNnffXPHs6z6bON3hVv1
To2NbOY3xzvrRbIUp/eObjhafYxseFcLls6WvuvVSABFDFkSWQs1se1v15SFVRmVveJxkhPweFiy
uWrHs9UbKPj0xlE+U+wU80/cOcdlOhJ36OLQwj0T2JMQ//YKEGS+jJcnJKnvqE/nU7VGwr23+C2j
E+m0RQFNRZ3veJNj3VqpazS8ZdEou5IlgiHFgIhqh6iBiPAI3z2ECOgy/aWJ0c/FEuFwAsUIkleL
lF7udJKMf3ujHWvRW4kDmh8HvWyHBFxmzQXxr8juvQTelSgEPPRy4INjd4PErdNFD1sJPsRWUtpA
Gj/zWfI6bdw6j1M7B6A3/g6Mf27gPgpBUqS0FRQiW7f+l+QMkQKlhfATpzyI10PsIaqxbq6+fGdI
HDgiZ9yIri8ka764/We2D7aBq1FkiMwEV0KaTQRYwWGI2UfepjSHF6gR5k1e+5zPsuPhLmBt/uUS
tAmcM4d1GJLfkPmSXd62PPrm/nrubxHS4ntyXHox5hO9PwLix/WZmU/yxnQJ06jr9e0SZvzV4Vvx
98BRre8W2AJOZRh9iTzbm6kOU+dh4f78A3u29hvt2N7K4qea8LrHLLV7kZQiDlK+I7JGtyFHRoJC
xWXjhObaISbf728FnuoIW4VeGEvtzTSREhGGrNgSJgwHheCJTJmu5qpv1T6a7Rss+zrjKWnzQg/q
vx+96hy4seezSP+svuMRGnCwE6iwk0eETsTRzayo+uz1AXs4fYTh+aQ7gX6dB3t7fUNUN7FabTbQ
BmduGedZA8yXc0kKdneOJoKhnkvGOHI9Ki9l/NzzRxbEcoRQWN9EFpyAyLLq+4XqloXYRx3gFGIM
dXeJtjY+xvcYYwx9krUoGLEdKFtXVKwQg97NQt9DNo/f6BjMhr8H86E3l5Ntews0Kq0SAsCyjAMK
LO5Vk2glBFjByZ75sBKYzvDoZHxYXCMbNCcSYBxVqEkQeLP4aj0YEIhHCFBZw6XOH05xNrwqGUDj
SpUzBqB8ECv2wOif38YtFnd29HA7iKHwB78qQIUFFoalEQRu7OMcGl6+TqE9M3sl6/rkzJEVxlog
zVSMfRh64mdWv6WEZGCu4xV9AnNSRPQD9A6VxxTRgQuIQvUJdjcZ/cCgwHyMfzga1WeHmX7Oj+yN
XtRx5kdrjQDvCSPL3dm6ECdyG+2B/ZeVzey0lPj0CSF1kTHAwI5nqIeWedTEOhJEQM5FDGOvXqLb
xVcNp52tLh7VEnKHGuKC66L3VcEs3T2mHy8UDIg29+R3VcMWvf0mi7P/GTecrl7aDiuss30+YKWM
m5lSQ4FnIMEaAbbLtlBvJB9uRt9j4Qub3DikbQXtaaIdxBs9MWfsmcZGnIjfMGBGaFzlbb62bW4B
p8WmQ9Fsu3gtHnP0r46AcUE9qgqu9VQCAzUZx/5JiCYFNBFU4fVC7gpXCaY95CkyAXSfvRswDwVV
tXl3bfwWn/eD4cY5Ua9TumXGERZ9Pb9EmPbwLEFG7NeRV5wMWbmSexZtoaZZPXJyitHYc6qD7Eo5
Bpy1TwrI141zCrqTPWqv5GD/ntbrN05WOgPTB/eO0rmUhXB93SINFVDKO3ZrEtu7aoE/h+rp0ZKc
XcGb5eeJfSzvDB9iHE11t9Bi1BDPmLrqaNEFFCLdSNxfJtCONYj93tK/mff5OLCarhqRTavS9Cas
oX4uF0EbyOVHzkENaQGtrerAhGSm35bw2+DAKCy26jxba48LIrBJCdUlIhj5DR9BP+HoP98QkTOL
c+ruTFgRxckx7oeImzQjwuw3Dk4h6AxuI5P0AxX3RqluQzKVrblYoZDrmKcYK74sMDdks0W5ctp4
CFvi/fvTw9yHT/2IdNnWXMdEyDeFbHEnRx9pULb7w27gvXFAhaqA0NOfY0AiCB/FK8AqjfZn2tyv
3vK9bY/6utJ3BzciJ6S5lURtVnfLuNAKvOG/N3XddBOSBQgRtvTU5xtPNOnPUrTHt5cz92NGUU4V
qNrYd6Bh+MSmvKlGlxqW9oGdDxk7W5LjgSg3FeatP5qUfX3EwUfRRtUe+1vQfbUbaQm6iWlc/TFD
kuU3jQMd9hfA7ubUVmTWLSbQn/qZW+Ro9vW60og0Fpr4uMoOsrArDe0DtjmuLvIav9TPOhCVPN5S
CDo/tYOG7hLM1c+34ZP7mNit5GcQmfeGKQ6deMHeSNh73a35WXSEfQCtq586M65Ithq71IIc3H8u
GZqt2rpVRyy4tW/xhT3EsMVHEglq6zWyKYd9v0pzPVJBWKRTeNIfqIP/8Nh4iqfNZIW00foOLjx4
Gut6qcU6ZM9TRJu4eoZ6eJcSH3D1O2epWLP5K3T1+IzPhmn+/wqi0NFZYYE9GvBhwmfotT1l3iBR
b7ibUrI/yJ4FbN8wQqWzPiSoDe7l/rmFivMgCXlFwdisP0/HU+mcXqmiOKzQUcE3ono2+iriQQTx
kPQx17UjPjQNrz7v9RgsieoL0iqXzo1W+6B334nCW4snDmpHKzSNdqbTRYKJKskEgxAFm3GOvaok
NrTiYLwg5UdSDEMoAw8gwJa5GCaCKC9KC2/DHJa4fqv/I/64oa8T/HvnBzDi+8sTpGnEaSfYS+DW
k8KaOocnuY6RI1srze2mef3T4f4HK3xU9TcpwY7I7gjrv7dWdvA0Vgy0gSBP34YjouzMVDlatffW
6UL0pHM76SU/9PDQOYf9Ytn+ZPUUi0W5lc+PDh2LGwNSdunNpkTaDL/NUpzNMPPPzGlLs9tWyE76
1gsToXus1ddvIVvoUWg0vHKbo/u1d0X/yzIjwQ/zRLxmOMkRVUWDp5xrZGE9pvAx5WEk48Ktqo0L
X0aQswhef9JkVpucKXM1nR5pRO18a4woKE6MXObkQBkDA1GA47KJenn+slugAX4kJ+PgKBbTHU8a
UaP6rHSE8u/RN/D0COi9ShhJpWiPYNeDmKLf9ch/+FWvtUVLOohw4ei0ebwb63UKyjNn+Pjnx++A
xeVRgJmW9t3hbn03fqieQi716Y/49uCsTfcyM1FZBpRUIQjturGdstTDdPm9+H6jFsdKfvo/N4cG
U1xDgWXrlwN5gWSDhTzuvnvtDSukb4+TYPwUYldVpdxCFN+UcS0GW407KtXxOVbRRLBj2827p2NI
Tcy/lg3F88AY2/y4Ge0kw8s2eL3QXWBtFuGapfRVjuquyDZ1r5cuBzsN/tVnm6fo/ieKGF7A3gWx
R9BNGEYJOWHeGJttGGATVtyBC8hFH56jHFFpNrhl3ufSUjn9LBNQUV36HaqfL7p/2jKb0jn+Lzyy
jDVJlgWshKy2H82l9C6hXirF4juM6gN6ylJO68N/L8DfMAsx7HVboQt9o4PHTajYRjogQYqfaJso
zX4K8ZhmiE9Qw0/KHv58S/1yyEy8xM7z4FhgK5gTR+MH77PSos4iI4UaJHCnuZdiVElZ96acByPj
Lv0ptQ6fjiqWFJJXoNBvroXHoGkwKzIMreLO36fBhePExi1Dqw2AQ6jFBoQzCJOuttqarf10S7Wv
E0CaK06jUzZirJlFyDeFrGr+SXpoQJRmm7NqZBeHwvH4rpKb4F4qYTyL1OYywS4ylvUcOw4C9H/3
ifwXMAhy3kh9YNdileEoeZSlRWPeSma5XqjVKxV5IQuNe6CqVRg8KCmTYq4e2hLI7u8840s/ESr6
6w4MH5qzXHqsOS3PHOkgO/QVhNFdwloxY7hPKJWPVKO9uG8LTPwv1E517rhKlq6HpkmU35fosYiQ
J2+iz5VLrCXm9Vt/dqqdrWIm1Hdwv7O3qBwkpoNTbYkUvE/rsR57UMmu9Aa1Ko3aX4sqloqXF4g+
Nx+wFSRTZFJ7Wvl/QVtINmNce92ebyj1Blibqk7oKUzwy1CndzRx8vYHvutwFlcyX/+88F5PJWgA
8kFLhibxKBi5u+axkeE5ulF41NTip55x7BQjuVlEKVZJH3UUzpuCbE36LJk+ki148d5IggapQdjU
pVe7zXxvm5/3xPWoNQE8HcL2sm285uRfePhwkH69zTzroeaGIOltQZMn+KzXiAFMUPaWJLHKoixG
IgZHJtyrhcRtNJ+1v9nM/Y203yHhkSxEqTNqT+NAwvYgX/O1xYxqKdTgdrEqpmRD3052+xLSmVXw
c0YLRIxOV1wG8egCL7WFEnf42mKGoU3PPpZ0IVX8ItkN/xATeh7ZYTJ1FwaGyuyQB4m76L57+Yh0
bMV87PpLVLnZxs+VhsDT2b3ADFjvtf0eMJ4JWjjXoGilfRm607ZvRp8GA1cPAUUwDK10zlhFtlCK
A4Pl0i5BgxUjco7f3JhsHf+OZFTajFZsPgbjalohuHaYE1W35Dl0zkN7iJBgsD1mSRKZMMRtViAa
6lXj/anfwVj6rHdXKl3VkuVaGY8dTUQePBseg5eKNy8BCdpEMfdCLlyikBUPPGoxPHP2TBb/lYPH
OORBEAIeI+Ti/3z0HZ5/2qgIQLnXxGoV3TMUKT3iOZYiuCWowzOX3fF0+iWOl96YpT5pV9bjr1yL
n97pikYBvhPS1PIiiZ4f1a4QV+p/jjlV+kfMZKvNi2CPqjGi/pRkjdcKpduGRQc6f6/lms3ggQWM
HGRddMZ0MGc2Xy9cVNO8XOtEEkBynTir091reDHst1oHUjVK2Fq+M73BjWb4rU/P7s3d5Okc5Yae
nFCjuZwVEwqHmXb3MNaF5tRGLZwc5TkkaoSRwZKZfYel+3dIkqEhrJ+DXa7N2Nyc+pbFJJYgM1sI
05/twNrPnRqIKX+JPpOLgyTm5xfe6oofGJYElf9nYqDUDLoXgA2GaDVswuk4HWnyYmQA5pyHpO6Y
NiAxLjOzrJ7h6Yek40IRlxZswNwVN50L/chXv4WKBvxuDLZ81GTzE9ArPt84Ut7TyJM8g58ba9H5
QlOt3+R8SXkRGPREHTrEBw0y1uv6eY+V1JIXBBReucmVE8QEZCpnZtBMvtKWjVHtfUEagqxUeXWP
Fffg75hdnudZl7H6h9TCmyXuIRJrbuYKAMXkpgUwljquRm0mWJSc3/vuaccjIYe+86r14ofRvzJV
6SKvyUDFqPLV7hN/YfbduK+LZF4P3o7PUGCIZWHpgSVP4OgHyt0P+xKuluh94cJWv/yE//i5S0LQ
C40VFdt2bf1uTgF+Pjb3JKfATg6gr12SS+1TvwinWrgjg0WzCMjC4KnQw+Fm/w0Wcd02TaKkvRfV
yfXvRl2AfKm7njAe5rxbXrsjDskcHtOktEuRMSKjcC4GhzhXfe6yGL6PlvAGUHo6iUTi+36s6hv0
FvyGJcaWgiAJvC7sBPBAG8L+VuODbzA5cups8lwUztaJv9V73JKxiRX69X3AVrugfwz3hu5lSzt/
eowbYW+r6Fy9kjb/VUqJtgFE9OUOM9o7uhvHhczwfUzmsejVP9UZbXO7vx/NQjubKtiNgCb5EkVf
dk9JE0NpAfTRfcCrmWBZWdTgqQT0g3putMYzfrsKF/oGC73tX4e6MsH+Hg1pzFc7PdngpJEbfNcg
O+AlpBoqZlay8yCqWPEzxEe3ZbmyI+L39lcosCeevQH9877uId7Z7NFGiQ6uHdU1mWFuky6T4tlM
QKffT0t29WFJurnqJcJCyYmML7Et0T36kbLxELEFj7GMgqFGhg9if8UJq+h8jOn/abpthxqvtZSX
AyLYIatg0SimP/6Ve6k6mRdUaU4UnJnsiKUvF4woEcAdPzKdRalLbIzjk2N7L7RVDWPXAcUE4DyT
Bh5Kci7L7fIo5twcRy7m4LkRZk+pXRg/wTCPTiO/dXH7+XiJgsjFivO8CAOnpgtm9qM2fe7e99W9
5lbP30mYZ4Tn24I02M2i97kmzUccM1DvH77OCSnqQsP5esIK6xpvxpPptcx9NwpCRq+lokad9xni
rgs7ZwjA62CfwJXKB88TC2UIhbJK8Z8LOH+1DxM7/PN9vvzT6lqJzCo9ulZttdO9XvfY9gSi/mW/
SqOhLLTz2+FJk+hBzXqDaRKsX8EPutTJjsEQfb+h0fL1/Y0WJBkuL/Bm8e1TdzxDIDdBjI7xzpJ0
UMW9uFM5R7HmpN+ZFTv5OEtuH5jIi4nGql6EAVUlIkEllMWh6JXX+2H78K4dWXK2CtNIFaDuMSmy
Yyhw/0lbsjt/gAiF3r88Buly0y6HWUoPDay8NXrt6VOvoFg5hvIgcna5gamgsc3YjSedZhrgKzNB
jkXDp4ptCeziBmCHD03VtFynSORGVPJE98e67QoLZYx3EUKpSwA3lU0YrNK5H/MFxpPSH9N3nva4
XH6uD/4pIsQidjnVVzEWyD8Ok1L+OKz+I9QY/vsI0p9NuM6qvYBbuPEBETCspnWWoaAREV373oWn
dLws/eZORY6GjxftPHvAnJgPojVNUCNxUDhCwBmUSPMlw7RofdEA/VdvCB/4ZA4pAkKZF0El4W+E
7AL3QH2T0NwT2cgBbfx2XCY2y4Nwz+cEJHqNce95/56V2TMNd9EHtyB67BBiJYXEocVp/ROWveHa
ZwiYQysnxoccfKQso6QBLqSybgacuIaz0ocShbm7UghsjnuF0+bOlU2okw43nujRhOCVlYOSiXwP
xKaKWcKclpJkt1RISBnGp7XXeb+vL5q3/FzBpil9Z4Kpi9C/F5lBtv0sWNlKAcnLwtItvVdop5rr
rtvnR71a25ccdZgbk7/n2gE9zELqGfXs0rmEERL/HZuIiO0VSO9tiu4xs475y+WrhBN7gnnJwu0B
LYzZ1I1yGv6+uj4CdA1SQwQMnYZEwYKKIDi8ddOaYw6StC5SCkvO2iuxXPWTR0p5aPrkLrZU/eSo
lm01z4xl3/2UV7Y8dZFyo62eqyebZ7j6s9UiwD/Y4A6PQ9sgDPiZSoygwdLrycPuOEIiJ/16Uw06
hNVi+yln4qlkwr72P3wJtyaMUMwuWfchjhvM7GRzUuq3NrDUzBUTGLWnN3xDIWXbny2vi2wOB4Js
Iqy/jL1j+AHV6hteN43/ZqSAIddkIZxWVo3B9d7OYRtGnimAE99jk+rXyCvtk4tz/ml3lS9QVcxU
o679IJGEbUNntEaE8mlWuX/RFilV6NvXvQ/nNEMM8EupuC5c1dDnLHu2kGxHtSgb2BSyw0L0znQc
gZuVuSCBZMKyYwfxW2tKYKt7KT7ffWbRNXGN91HobgqqWGjWR/3WCa0aJQnQOT/waM8vkHBl9o7Q
lN6CRpPN/hiXINXW2qdVTYV1qvXnUD6hBdM4WKkKiEBzXkS0J4G4a3VnUlYdCivnwZR2QpxCJepv
9+xgc6Sn0I/Sz9LWrQ5vVEglMjoEW9qLVIz5iDNVlZGH1mY63F4aOXkuokwbaJtHF1pw0JVqWzD8
ObLLSHBjGzhN3bbv5nqcy9bfK36cyhERf/ZjGRbAdTvwIV301GGNMp5Q7cHugWHoOMZMu/zNfj8p
yJvtPDY7yNwdxhVR9tA47BuGIo/Nc5+wvlAtJt2TZCaWU4bq9093IuDKuF8MxB+l2hLif5mL+qMM
RbXWSUt2EseF+vQnwpM8gqO3xoqakax1JaHjdGGJjTNf9EV07+z3OiK5VgObglIfq47u70llKdt0
NRHHrxETfvBM9NyXQJ4ghG2Lw6MjEi/p9D5BjFOlXhEHM3eJTB8EFynQaFXeln0XII6teKPFr1KH
xHZSnqIRL9KPU9JHhyr5yc+hbel+1IRDNrLt6BhMK5n8TA8EnSuJv+dLJvfeLbPS1/lagk4CG+jm
rjdPTngnhHbur/P1mIv2MVRKDg871+n+HIpRoNHOUjOYoodDN3fD64cwJC8AoKnAOGkY0Bg+xTPf
YFyfEtf9byNIlGVYMcQI9uofJbH9skjXMOrfg7bvPixPqQIGHxb8ZeQ5nshC+jPR+H+9KwfO5363
BaHn7qky13914YLfDdITT/TTs4aUw2uG8T8nqveo8KrPB+DDwjJXPnZbBWnHTQ7SrdSQfR2BTPxP
vczibyiotignB/eiqJbVabH+HpK8kBPktwUPIos7JyX0Pu2RQgfvPhJxiDeRXg0HzPYzc8Z8bHh2
dxM5kvvrFTjNft/kz8/8k3phj+RCuosJGL+6H1HsMRwF5I8NAcb/si/ypjzv6KKHD8QKQ4K9tRvr
7vhFJt2TgElxE6t2fPqZmvS02a9xdMDjQ5NB2ugegNgSsSXmdhUYdxcTV1X2m/v1Qxt0Qh9thbNx
N4WM9Uol+xA1/5EDdjrSMc8HupfZEtabG01hR05pv0XZ2EgQ7BPaoB33PscfXZmMBmKPNzPmqDIY
rqu21YC8YrfqImpbqgVXsAgOomLkiXAZ1vizWW66vkcoLwLjmROFDeTgFshCIXcxmm+k8jlyUlUv
AoICbUSuGvypQ/AzYTxSmbpCYxZAMyPlEUDJbl0MVuEXfFzgPxPMZqLBgbclgSbGwGaCnvd8JDut
JbuPAiVZMZWbS5L0r7WyajLUeBp6CHRZRbx8sCdro/bx7427yDF0hofwgAdYn1S9VVjXgmBIRCKD
HlUv1sOWtcTDYXWMxheHZFTEtT0ezOSOBQThbGjJRUMPONxavycfzQqc+N5sYrPXm/Nhs4zFcaN8
ylvqx3TwZcZ6c2o2SyJUSpbAkZLYEnKwjJSnBQahI3yagotxZLhfCjUExUXVHKhHfU2OXs8ZKgB0
Ivs3Ot7IPYSvRsI8uMm2eO4IdUbJLgZFSwNY+TjTPKms+JXDr0rfCI1p4QQN77Jk2VrotQO92UtN
GFYvfgUUYxxli6pvMwbh7E7j1aFeVR88IH3V1I9Qda+rTU6xjvtmzQK5hdX1DIQSl9M3G+5yw4il
7EUeQYVXt8vOXCh1/dCHaDzSiqkjDDNd7DrueEI/q+GxUCCPxgwierUy78a/9TpoL5ZgzXhCxVtC
i1ZykDJtRr3MOKgOAKTz8jtmcAABUH2Mk3S5ayy4wgNX6bksBXFoMiOXHb3DiZDRR8hvRNdNMaIX
fHqlXbEc9ooEaZS3kktpJ/9GAxem6uHq+194Rk1cpYHzEGZ6BYGatz8+RKql/FcQhZer4VZtpq/+
z3FOzJUGMKAk0um8pADdDWEJGKNRFlO0WBWFOMRvuaAxkRbhjo4HL7GH5hsMoB2IzEH0DLCTTLg5
ipz5QYJMfz4SMIJN7qGDbkJkBHrl8hdv2IMOs0lfQxKZQmMnOrFwnkTdNR4ZOXJao+s7uMe913jW
OhD7VYXJm6U1fdRsCAEG6ble60iHHZUv5c+smV3I/qfAYatKVSNib9u63yNmzxFIoMwXivLbZN/q
0WOPEMdYyl39p1RcwwOnpWkzLLM2wQ7Vp3VNHWTzUY1GG2NlJUbIQsccwgl9XyOsc6MpwNqDnue6
7UUZJvgmPoCE1P+EZQ9Gg0DWfPnj5/vg/TV5rnkw6pPVIEM3kwiItFfU00xoBHS14TzbJz5F1jej
i4Vq9G35XuNLTBgCP8nf7yXoDnzmR74xYn3TmOtFP/xuu7jVCt9CAejDlzjB0T8WxYCwPibSINVW
kEL1kjMgu3HKb9BnhQsvmTWFLcy5civ12pdb2mGv62KpIpdEs6QD1ZZlSrVxqNMN+0cz0vnTbT9D
oUy8olSilhylR0uzXzWw0cgdC3w0/otQH8qFNg5a2jxtam3ogj/oglojhiq12ZCXWqmaMwxdWocQ
PU5EW5QWQyaQpxssXxy855QOPuCpzqOiUh85Er88XK36PS724+/Q5qKeja9Myges+XrXTwMV7j6K
3W0nDndFD7j3nJ+Rc2gJC3HvU/Wv6bttttPu/RF47QzjcoBDmnzvbIkp3f9r8Lm6546AtISPFcEc
eS2W8Fo7zlUn4FQ/b/2O/eE+BOxwqZaU/qgtDuE6eqc3jQ/FilnAklz7/5Hxp8ojcai8p8qi+nWv
GSDhKU1cJkFGh30z56D8eQ0iTToORrqHNGiZfC6/eQDjZ8IGi2YkkSuGvqjjBRMf//8oMU1pkbjb
o19qPAu8pFLky4wIXzfFoffGS09JHHcdYLl8/U2FYO9TByWPRKSBNxPXnHo5FcLnvGlxzzxScTUn
/Notx6B2GV7yoAuffKM+IJkxNxlbzR+mz6Pm6csWzFxf/o3ydx1MmWwS9XIUs0vMnsh7tQMkwTe5
+0Jz/OG1LPlOeWoTsSxYeUv+UqqZTQ5JADxN/2J+x6h/Cm08JxfTZFYK/eQQK9D5devNVopOBYLs
JLXi4LgNiL1TBKcBGAOojeje0D7aLdkCsW0Wdmfg3P/PFZs9fbr+k16tluFVLsQdGnn6cgndOaek
Fvccqi8sbh7knfeuFvQpcI/iGOJi3gxmQArCe9DV5V/ylM/OnmnGKC1y1g5tePeQ9kJxrz8ye/fN
si1tU+OjvqEJ+ld3c8nFWBI/qPll5lL6q3hm7vMcAJG21fCPfbFoo7jIcy6ysivAM6GqIerKuaJb
bgfdWD3Tw6mbJzxwdJJx3Rwrbjfp77YKHIVBsAKZIpdUc0PNZerDhOh9K72o0Fp0vbAnycmmoSKx
s1SWZuzJSG7x0uSdb3JOkEbNsr3rUWeI5eSz6VPfMNP/2mEawhWL1KqfGTZDKiB+UNMDwN5K7zIi
uKcihOcjsn5AxvurhG35uhCQEM9AcN/LmyVVZ5bd3lC9Rz7iYk9gbXhljNEFFJnquR/NsO5BthB+
pCc/BBCjRpAwTA/qOnDcxY6Tv/o49Bv4ANvuIWcVwXIZny+RqJLV8RYsK2mB75lRQOxpfXZxEnyh
G25Cc1jWEQDldaMDv3JwvD0FH0ea4QwAVms7zK2lDqhrF8czcq1GzFtwwb9VpRN0K+4y5d+Eqkm5
FOmkWavZA0MfvWgdMffCS8DOT7TcJdi39pZAwGCpXaTWofVa+43GjJh+wgpUy9A4vK0Wn5dXXMvE
PJANsQMErt08tVmMY65SVb+0WQxmpZFx0A0D6EL9cc3MEocTbvY6kULMGuH6lne0Tl0mGUsMaKdF
c5GBMjPWFdWOZ0UoWc0oU5TjxXNZzGzWbF9V+YvyJ9PRM2cOxQC4F+oiDTxmBLGGK/EfcdqrJHMt
InMhTDFLwIQrMRE+cNIvweViNhAkXT8Bc2VoaPUt/WG8EF/T0XuIQZPfhEy04SOmR5N1CAAiv7ph
+mg+YYCPNFkzmuVgyUSdpYrVTyWmK/IM2LOevF4xvnZ2AA9qXyyktSt5TBeDidRuXo2ddnkNj9tF
gDcJ0mN2gz5SDsvb3uBEhzIBw/DO/LGFt8Kq1WKwPYDT7u2E5ygyK/HT/ypdLOTsJO5odC4nw4KN
EWmAzwYyE4m/DeqXJVXTLRNoelmDzkPsR5S+FzSzzO+0GwqCMS5uN1HpkBgniXzwCMVtjCD9eVkj
L58uMjQvxMpduiYRhG6rHFsq92qiwoGGuIrZwRw5197RqEHObZOupzIvFOPKIM5nNNeJKP/h2HLB
9AQAHjYk+ebf/FWM4K89AfVmm/AYFBLGCKxq8LVeVQGhNRjx7oMeY+wf4szUx0t1t78EWFs3VzZm
jDBAzfwKb+IXmYt60q75d8sivB/oUXc2ebIP57wXYg8noy6zQBeQR5GZxDHNklAXBpQiVejLZoQO
4j+3Sd3WwqWZHAquGkraRA5RL0sg2W2WEr45TuEV7jTKv/6m490AZgwr1/inanfnXunoK+PHBseA
x9a0j/8mCyrOZgW8XqeZYIvNfoVs9vddkOa78CzFvHvdgvBKmiSNIsw2yXzw6DTVLWDzTc1551MB
HHRDTLs0GD1MU+QsRL6kQz/BZza2ez6N/AivMoB+EVrgthe8gOms0UtxkXstgqQCmnj4mMeKniVb
rQI3jL0SmU4Xy8DoDSVJ83sQbhkJCR5wvuQr4dW75e7T8lo/cdRsv8extcqXQNnbaprdyEYggJ8b
F7SiJSBR4wcYYCZVPiQl4Wpt13B5z3Q5f6IM4MmoIz3zXemBU1Fz0KfROlW37+8IYgjQgrnKs3gL
9QCsH2ZclU3AMG+Yxug64TgkoPPurfoIfkBdfp5jorAnkImMZ6vNDKYXr5CNhP7UZp2FOhuIsAMm
+lNS2hEkuQAWe9tWf/bhNrYfteXZDi2AltBXw1jOT5KtMPcEBFiPscFokqP9pA8lEOnELpcMDMGm
ANOR4OpQx1GZxafqHPgQwvVK+H2Ku65zz1Sehub3OtjW80xzmIcO/XvUT0nKCnHNjwko85N+bNOd
oczc/3/jf63VTMEnq8ZkfFC9MS4QW2DyZtHJ1rCTqD6PTI4bNQHQw5bDPvxTnHWwpk/CnG1kKjzu
VcloeaCcuuBTZhRiXitv+gxYVnNADezZ3s3lJLYJMh2lzbKoWjDpmj0WgYO0cwHex078m5Ttu4+l
BruVDTOZfsp1a6jRY7KN+VhbD+DLGgD8Sjm9pF2s8ljcEauzlLDoATGrazeAN32srHs6dEbum5N+
MwVsYbmYAcX00kyefBKaFv7fKNDx0YSsgnKqldQMVjt3W+FxCH9mrGmdhiYOZPGTP121a9IwH8jh
OEsGt3191HRoyLlXqhcMbrmKVlWp4o9Z7yRtKnft+N/UhgJz7HacgGtz9yjHOY+FNX23J73K3/4X
0Gwg6PLf1A//QQzfHJsFbIZJR07YjP/bBe6/ioYgrxh9NPp/v1BLM0eCpYnSEUTw2SuWVVaZhpzX
C157vnKFVlxcmYWYXxzLQo/Lx/vE5v5mg3/fpS3duTHJNPC1rk5uVBbS4KmfyX0G/78jH1SThwET
SYfiqxjtW9uCIgf93qj99RBTyRpBeLz5+4Haa00pdBW+3WDIBTYmx37uQxuGLHXjRjJUzfPCvccM
KlxlhO5VOUHkBMq153dwOR1MA0S6EO3BBtyz9jMgmaDETqWgK59feoaAk7xXzHBJ1f7MAI/7/aFL
CysQMbV2Q28h/dhCARZxGwvjCaHs+EvaW/qEp2GWKUJAMZGF7NBAzolZULLh3xNXq/wAiG4oVsAr
+ptsk1IAMTtz7W9wEZvciGEUTk6xyt1RbuwPDUPhAOI1AvM463ucIO8q5qK9gCDGH5Q5jW1ORfqn
o0V//wbDeA6xufWbAPjHZqXyMVRDfjCtemDWeTshrA1BStdHteJTaQFAuCgoP+zhxcnHvQLnVkV7
Aarzmo2cplgs+Aeonuh+4rCYJJQhROujOl9fWvxB3U+QXZdcYJkKpDD0ObaosAQMnYCg7ThF1/7U
qzcicsrv1CrYKyfLuHvtt282jaCn5C3bsYWOW+qGxVAUHzrp14lhqDCI2/WSnuYjkealQqfMZUvx
Crd9cKHufcVWb3yB8u+u6K3KOUUQGIu2bqhiMuylhF74WBaPyRsxa+s8WXMJHSj5P8DZW0mY1XSh
BoSuNGX0HAe0bw9zZR5Ex/xutZzUa+vduIZVOECCQKf5bW9ci0ea9GAvMRbVfONh5uAP8yzFOA6B
ZribNIloCRG4p1OYFBv9ix1pxknqkgd+jFHAjumfdDbEoffj3j+lpuc5ER+q1gvwsAczzZhBbzsr
bWVfFYAjACKpedmjla6z8ojlU3f+LefQtXIEANoG1/TQBAYzlF7JU/OSJwfQQAiDi69ycuNyZBcJ
miTnUffdNtC6eruJt0fN+iCowCwk0LjlAirdoniOPMOSInZHTQMzvlq6uDjJTV4SUGfVjtFDWwws
s+nvpqfZz1ruiBeWzNyQkGs3O69vQXbsznDuLUJyzkrdN2A9yPaQtMpEdLdToA9brsmST2vbRKAr
TCcsDu2VBjP8Oa24tDSEXtBnX0aTeqqvZAHsOKSv2T4fEsLuut8Nh1XVp4B2iWfYzq1p8JQcBElM
pDP/diNWnQQe+Ao0kKTtH0mzCYVfVdXcwV+e67X7d0BdiX4Zt36vTQMOMULNdub1J6lpd+s420am
6qHgAvGp0reulBO3HUbGOYyasmkLakDdxAnn1RmsjJ4kxojbNhUUPb0N0xEdbxy4vWTgR5hcrtzL
dqM6QNsRkndVNz0pooSXqTaLq66WN+IXcJVvwBKW/agtkaw15vGy8+oGac7YT3QB3hrKniErqIq5
Q0tMEh7omheb0LPi6umCPc+ccgVw0G8fEh9xm1qmi10GRmGOGmB5zdBFznBpZ8ODwWzsFpbXeazM
imB3mNfWt+wIfz1P5pnTL7wq7By5rSCGED6l8urs1BbJM/DjwVlzjW4Tvgry9w7TQ9L6S+jkhw2L
NsTucKwYDj8rgAh+NvcSe6VnPSF4IlY8J8PZQy+2Un02mTkOPQn171KgxksamEZYD21Kzi4nGd5N
3os+yWrW/M1DDJSyJokXu5xZe3Esispv7eBTgCDk0M9gtiHD6w0ypL6OSXVrVu51iZ7XRuCdffmu
Tjw19HLPWPjEZavff7Cq4w4hOlLbpCVk0+U+41uI8Q9GXPD4gyquoRp7nvs+XIhnhiq+miJfRj1o
4JReZQ5eLoyyIYkqRKVLhMSrU9uzzwpq2Lf+ZLlxUv4s4Jd2KMT0RO1pyGnzvHaWJ4V9f6befxH7
LK/w5t+HnqAQ4EM84F71AMXp1boHrCGue2z/sbt4LNzR6f5hQVE5aCULnBZKMBCqXMh13eQlNaL/
6ytsUBku31TzAKY/MjLCwjtDcSX6G0VNOSrBphXEBk5+kaGsr4KgsocudBggl1V+z17PTY33N7kt
62jwKoyraYuOsxVN6fiCr7mDhd50Xg1mZ6DvvM0x0EMhCTEqo4L62E97yL/qJLCHcO+0U6aHrrpL
DTY3XSPruBXFfS7dYAlTu/Lyorkx2YIhdbL1cB06YkI6XUscLrT7gjXGOapJ6v8d4o68YejhJDHv
fywyBLa8S5J4bQLyJjOm4zurZHI8K5WdVzYPzV8786DI9mzpTnyCSjFZA/AFVAYjVMMef+po6REk
IY+glHYtaRzThLkdRnG5tZA5Z2RpXz2NvPgaVMqSiWPRQIYrqVCfsGJRKr1YE+S6IH4v9S/AmrC0
n03mk+nkTtUsW9rIMjr9rigrtCFWjLjAdb7glwryqmr0luWgakMMbmql0G6WbJIBqqYABkUh8MWe
f0U3/vsSpwMq4cpFKYjeJLUunrQWhLlffc7Yu9aD6hKitUWKJukv775OJHqGj30IU4RzEUTlCnTU
m7Crg8zJyrpCkjV4O8j7yUW6GLMyX91beARIzqc5a73FBrGMZWfnQ910H0WUNn77nc12olp/Z4L/
bUu3CzKmwH4NHeFok2HchwfwAtVCmYzxVGl5IJf/1VVq4loVV2o7YRCO66kE29s0qvGGhXDJA0gJ
0znpXhUMpK2ZRgK2XW2n63cB7oya1NGhsao9xvfLS4gFtoM8meR9J3iuzbNZMuH10IierSQ53Fnr
sspVJpJkVfso3DTbLM/6qj+I8hD7ev/ctfksjMeysNiTG+FzM5B+0KPf0zSvysQ/OcRFtWVhWzYp
G0WWoppX0ECTbhi2iKTgUX9n+tJVdKZH7K44fcy+EVQaPgIdZdPyfOsdzG7E8IJdgfnsztnj/NKp
mZi4sxmaqP6lBcOhKUB1Cf1YtAjO+TkfAr0YNDdx2HGLjYhn+oVk+/yyarhoDWB8lyFAe05pQKja
wvs5+ukXn+tNKaURSWlBO03gDdp+7m3frUh7N2qXiBwumWH1zgGlTMcSG0wQBsPySBWx9acKn9pz
JxtwkEIwBz/ZDq4cbVS3POcCUf61ftMgvPJEru4guuXiPTrn/4rnB3KWSI7OhuNghzWgSOR/t6CT
vaXXqtr7ULSgRFrphF0K6IsxhyR7R5C8m/dNX2MTUVebQ12A1z43KK5xlQQIOaoWzPu59u5kvn2s
MjpjfYbdQdgSecpDBZjfrMLVzYVvzNwoOO+LExuu45lSrOPOJVX/zj5z0jdOeMJYIceR8rymHr6G
CYPYw6Bij9kobNzsBxPnm3Z5gj4Vhg1NmxU2k5fu6wAejXrGB0ScqGoWxs4P6jZHM/kpgGPF9iBx
ts1dCV5MSaMG21kPfI4hurNzL/+pagKIHDry2gqtn0J8oLhulswO4+yodroeWoZQ94PCKhijSOoG
B6YjGqvaJtTnYrklJMyB3/POtrrozDI1J1R70ppR/De4TRDJRIzE0wcBTtsNpRTwcvz/WWNc9b5O
ucki1RxJOtSsJYHPlqmH6Z+XYNePJHBDQdYV+yTamtG58nFzzOV0FNANDv2iHK2ufCRdow53CmcG
890y2dh0+x2yt7rerPFAXuJ1/NsENKFRHKN1RTL2FAcYX8w3HJmGl8IE5Ue2a6MJiwHyBFSCm3ON
CddVq9IDnvCG9UPsg8JIqJMbumgKnRCI/R6YrkmPDz477ZhS5YN06LxOhta/udF/JMgt4kvpgO1v
IxngMuV1Wv7dAjhY2oQMFylrDo1EBxX1CNHd8ljG7wYuMMFs+s5Wm9/LM9u0k+0RP4OqpzrQy/1+
3yNrfUipGxJERBExs5naqJNLzUJdQaCiMYXCppjNQjkCaTwnzQfrXbK+AajEoqoU9VUtttBZS1Fb
x/oddFnNxmVWTFb0Zvmex70Q0IkIo5M/79IWTBwVyWz6A5LERMu4NXam69v81pM4zSlmD10Mboqb
itJyR9ZPEWAIkSaCKnQyNy1bv4WVQyaWA5gBCYMjFEkvLqyYHy39DEzj/z6bcJuaiOR90dgUlZUd
B/CQkqkurLGWjV9DbRnU+3TiYtrBj6o6loTSIdqzmVvaH9EuCrZxtdlwaGVjmdtFYTvrKOLR28LT
F3cIcOYE5ypj92Sj5bJVmNN/8UCwug4wduQRmtTGXQAyttLKR3pdRUHXBBHLs+OQg17o445KInmn
iC4EJhZeSZsCKqelVuIYv5JtMHxAw7/k9HrSbdl5KMlGIzZ2k2gQudXabjD0nO5IDikQm2rQnoST
o99+5qNOgNtOSB3IBtUuYiB1ypQYUFbyv/oS98AFVf/Nl8yJSFCHv8Ssgl/QjfMrfKIDyY3v9Bbc
DgAVr7XlzrRynmMDXz2tDGqSdTDmA0GkyseVx4bOmAUJUWTgRQrcOQoi4iIhYpOedpqsluH66pg7
FGn0YRfayI6a6hXvVph/nj8nuR7lTznJM1ai1FEyBMvn2CPbSrLOgeIUH9XiS2fc7GL+47fBAVRk
jYSTNbk/2OCQK/DeybtZQySkrh9leJ9mxYjfcyF6f3KgLTa1nVOEwEPyya7VVdpnzOafKCI+0g+g
F+VBU+4eA4KakBkXo8+ox8j5tDvu/UwofUGqiLMHa/4bSXJ+eZIvO6h9CAk4XbohMm/QGILKCbBn
hz9z+aeZfTM6UAUOsM+K/zf6htNfDSNbDXVhN/w2Yh2AhO3HCg+BVWjIKnkry+KxXz+DBQOCx5Qf
mBMMLCQZwRX+NEYre6Om8DrPfuU0asodKbEiNW3otcx82WEQ51GeZOZ3rkMSHOYv+1N0Nc2VZHTv
sb8taiDVtOLPys9EOIjbc3rBfVxefPSqge1teS6PkpELqNPuT8CChTPkV7WQj4C4CocGfTgrKnvp
tmiQzMkep3j0nNWBDBIHsFE2H4bQn/9RF0q4iuAN5LBGdzB1CLUZjiHa2rvohNDTs0lIKKujlj7u
LO1fsYR4tDLnG+xP6rzdflB3Es+pl1Hm8MbUvj0Q/Ve16fkj+Hd2/kWMV7tSQlClWcUz0VM3KNeJ
NCzdegi1DAm8/c96jbNNxZjwH16UzZOmA8pccdu+ZTZLKJfQKzINNPfhsZtTvXN2C08dQk4e+1c9
y/cM6Gm0HLgwlUeCUC2c54ESZiAIL+SFZh8t6jD77LZ/TvbMPvyhjl9ddh6aUSJxnSHU9pZP45bO
D+GA1MB10YDTE1S/vbq9OikXQq5eo6xi3HYofrwBVxl+tNXIq8a7XmCZY8gYC1PB+4+BnKi6QzGS
Vj7dpWYM96E2QWBj1abumyn3ZaR4pjSNJDDEHJJcaM88rHP16DLkO0lwLg7Wex/vh8S5bX5vZmPE
7weAkA9Vv1+sgUbmf1nd/aMB67M5YrAEq0FaWdyX+nwoP1adbLufSaAa2kWLfr0+XLGWoltePkgT
BjHQyWb/p9wC83/nD80u5EOGYzf0Pbx5SAOeE+y+WuuU+Kwzd4pXYPirDaYnWwwJ9XzxUnKtMM3v
BeCZxX0WBu1UFulD5RTds4Nrf6l/Ayx1IagIon9ECRiDTT0U0i8lsZJJKB1wGRrQbkF+I4mb2jG+
v/okBuVoafbim2se74MGLYMIVc02IqXRZYvHNZa8blcHhf2XJA28xqIP3Vh4yN7O3PJuBRYJU4BY
RuCnwt1butG93gb1pf2yhQO5IDIQqMdw+0qappJjsAufs22dvsHuSD+NCLQeDTWh31ZnNvrQVpTQ
Wcb4ol+km/smt8Vmyu4oWNPI9KnXfVPjnOnqZWOHf/RZ7J/PgddxdEspnDYJokPK/DLqf4Q+mejD
RHNaaELF62yjeL/YjQ8lkgR9mHtuZjMSr8FGZntDprtOHe6K3apXK8Jt/i0WqnXfwePgZK8H+4QW
7f0Uh21wAPVXF9PMDqIBTq3QKMNzKOfH2aZGoggc2lrODCYrn5aK2je6w8vmFgDgE2evBN/DwBrY
F7rA9PLS7I8HUv+8/wl2yhqTcyXawDvAfxMz11i9FsfVyCQv5D5DVEuHp6zxr2x/p4JdNmBrDK8G
wMRT/DzIzryvi7+zpI6w98JqqNN81fYckqkGdnsjc4fYCeFHfq/Q0aIKH29yKfW89Mjm/L99yleL
JHwanQmFX3cYPqYUwXCyCTEOTj01b69U7+3uEymK4RGkUSHzKOtj0IXepZ+QfbbhAOJfvP/dNufI
9xFxrJxDybhLP0B18EvjLLZik9F87SRRA3r6bYfeJaflcDk4pyv50+K0ToJ6TbTvlNMu72B6RF0l
CehK88twW2pma0yiW1iFBYcprf50y4twQbVPYvRMOYd0GB2dJuCmswIL2b/P1TgP8TNnvUAJxhRX
Kb0kWRYOQ8F/DBeXHmVxQiAxNE/Uq1kCNrtiRICY73+6IsA9WDB/K+2x0Ojgx74aEm+ULJBcIsl/
lwXibLMreYgA51H93SihXQ+OJB7PvIjQ6vx2w4/DFBR67yrduVAMUBApSurO5c72nN1FjUMzSkNl
8dYyfWzy75B/UoDRkyIB7SrozxJk8FsAjMmE9MUCd1CVXPD2b4WuQ42rLGy3VZlHlj2k6nU/ul5a
EwiAVpJR9AbnJISRzZJMECxXtK/FgZ3PBLEqrSC5uO44Rh+oU5IFRMEaGvmKoUn0HoUEIuetMTOW
mkVwi0Vc+53rmFkYcA6RYIl0uXZunTHPTEvbMIfy655Ps46KweK0i+K6ZEP3xMxSQlNOUpoYbCvJ
5aXLwgzogw3BhgdD2MLDoWCsEePvCJAxX885yZWUJ9OBA6FQPcpQ+JdCcKKSunlSrxYphB3hT8yo
zA0Lllwl4houCF0SMyceQw5Qr2r1jCY4SlLV42vAXWBkSSfpE9EthE/OtWwTUJd8E1SqeNtcW2CV
0j+5vvYRyc448pZxdlctlySrg3hBTVV5ThoXk0t5APaEvnBocjDhDrZcVu+96k78t9eGfkawrxWa
Csv59mnQhKzs0y2lFm3krRoNVwpzbVBM4RwYbbZPA4wiQCQkPhlXDdD5rl30rBClQFKijFhrXvLZ
Y4uJQNYgZoEWJXDTRM9NYXMdPo+buLU9a99De1snozCQDAzoT623/8rp8fqYISCb95T5zgILxN13
V4HwXp1/gmkQ0quV/sN6Xn0qgc1QQ0kmderiuzcx97JB+RwiYF8U0mHvGQfoXPcE3Qi2mVEY2yqx
oqfIKDGrE6nI+TI5ohgKK40tSc3rizElUpObpHwmuUnBlbJ6Fl95c6l4Hr4F8pgVZndP4+Vdk857
MAfOA2x6wDUYKUOREknRn5W8ZQj3Liw7sCoolzV+Ny+S4MzsuvGYQ4hRg5XRBd05UL8YEOcUujik
yB080+27KLipnDZP00SSqQM+97WtIouKtkTJgiOtuWdg+Og9YfxgurahnFW0F+u+s95hhx4Os2F2
XsCG4Vu+siiuPDBEPRAyrD79rvZMPnj+AHOcD2sGj3/PWGfWBRwXS1nvwUxLh+X4m2ny1tqrGpu7
V0jrpjxllsqwKGZTzw0oOqUyp5cfmwkZTDgAH/MergPKTPTOSx/fJLC1PF1K+nuIl7BJtePiISL6
n1m8g1BYP9JI3FwUmNs1Ts424Uip2oOxdhTgDFxOd9vCPhNDrhYO5BiqYy3hUHdYbGwCeCiHbOQC
SgTI/G9X0l1PwKHxJMrdZsUz2YtohCsDOb+ugPUdJVjrlG53iF3gqdqVjXLZnsBkCoUcIBJiXxEW
2YKeaJ6mnyFlxVV3ey2DQzapQDAXYKGiw1r/z8EUZvlNhi0JM581CGL6BPetwJQ/JtncXD6s/YED
otdbgD8V3DA6vXc0p/+TnUiRFs4aevTMtLlumbJyfi5map/eybNGgpTNyXIx5P63EUQk3n3JaZv+
HY+2kQygk4bwT8BaHW1nz/hDnndRG0/PenxH2BzHmWV/TDZQ2rxNg60crB0MWv6bWWhjt+smo3M5
lmR3Ys3ZbwwUHgaGh+9xaWjkKvGKpyUkEe9NcnsNs0v2gNWSz7wjzPZHsa+08caU/Zt5gOgcv4wi
BnMGkKYUrXmUSlJ/v2y8hHwnUviVjR/q3pbbj5IUG4X7y5VWPY7oaSbY3+BtGXEliRvGW884xxHD
VTiGFq2t//DRJO+UBpsziNVOX7wv9fUwLSQCL43n6MxG/7mqUry5+Na2CGjYf00zYl4PFGFaPKyp
tNi+UFYd8yoD2K5smE3vk65bkd8Vd3KMbVlqVUvkXd5mpEqkdisu375p7VmXaLHWY45NXanFmRhk
3jAAAt+/GCD1KkQT4uQRG+eiVclwXZPXlb0iA74b6sDylt0okxYrNXP7M/RF6ffelSEmEOhbeo1U
e1kUbiG6QYve/gZc9eR7Xt/AkLQx3sHdJ9TyundFhsLvW9puHbuvll1ksyTWc1mK7O3BD+kNz+64
4lrVs3culrSpmm/bP1cSwBvoYzcNb/dcQsp5rNyFwDCnJ+DHxUHZ40Z+eUo6AhRydIldzcsxbtgg
qN0U1jkbEFQeXVUsmRRlzSCRXGztfm9dZMIR7jHQ6fHhfSs2cZVf5C18sSRFjKaScsKmK1rewOoX
z5FjCQLJrP1sijz9bs7wwMhMGO3pFeC5a+X8f81XPz70yWKfuM4ttNSK/dy0+ZfQ0AQmARkwnMG2
gq7kC1DnEDMiTbfuC9dmUdmB+mgduubiDL1eLzJPwut9y/SnEUecesggEAymS788tAEhjfPme8B8
eCHKSS9pA3SlVQYcv2OZa7lpIpDQzjngXrXcVYUwtOMK2xIA/ipPkCDgey2gUP1k0nNxb32yVyLV
NjWpRKjc9UlDUDXzwAtuwkgs1UPI7/xvVZBP1fyepIonDXgpgihyoCSp5v4aA8t6nn1GKZwQVDIl
rsx6dC1SCBi+Jmj4U5IaxCx189l5Cy8MPA9re8NbQmHrb4IMpmjfSQlag+4LCHzD2wscgpoSC+c0
PlWH2CoGlJU2vWJ4jFy8ZwgdQh8PAZA77u0aI1/Gw3/e0jMhOzslEqsHg6AWty4PY/9aV6w7FmlJ
7U0xY+Tm6tqyd3YkIBkvOcXmGENy/X6eKbih8dPpaq3mYqebeX9USF1qpFSixEicaY+cNw/9Lcb5
Ni/7UfsQ0nMT29SYUuDbXB5tSoU8deIHTbk4zIt498oUlH5DqNKJJxKZbeCeAOTwYXVKRI3n4Nc/
tJgpUCedfsarPouIPbUtijwUEnOK8QCptmJg0i3+lKVpyZ5LNGub0OumdWFRkyu/EojNDYl4LrRO
FQllcvzJW6gyo6ZxMqM5UQwQhgjSdLHCXcipoyQYhT4GRDqmJYTKCZMD1igH4hbzB3t2vItq/UnV
5Zidfh/KjO86hr/z/bkQAlAWlVLT/V0YM/Vt2FldH+uKzUsgydXaDZ3qvDcjaf0NZu81oz7I1OCS
+Po23c4I3IUSnFuDpGy5oHO9gNsCWjFfWOdqh0ltX1DsMjhO/G0WdDuRcQu2bEO6oTVOOVU5AmML
+IVLLGZyMAPCQt7XglYvUj5Xo84ODZnsgWC+06+1WH2StKuNToR2B3fpGe7orl7/SCD6pm/v4y0Z
ZcVCjBWoKLSlogtaDSeE2d192j/C/EU7MXyByeIkHQvTBAMDBIOrEM6vgRn4XHekq/J3a5aYf6uI
WV/vNCM519430jS7i4POHejciQxsHSot3b2BYeb+G51zRnwfYrOVNIYJZBymlP3Jc+pSpF+/CTp6
ctIMwpCqpiKPLSOzpG/kjrJ40habNjObQruiuN+X+04vfSlBWOL4HO8s2utIM9BLURTHSHBWPQfS
KUi95b8EuXOaF8oOAgmKveDkF5TBuw/svbNOny9gfVjqL12aE+BRZpt/A1Rbdx/GNYFvThASJCDo
QiMakTV2k1wCsEtejPJ+l/37eZ1jmb9/4tEo/2h8kxHgWd3etyuV0maFOTpg7lYVpmgGqEV8vmn2
giCvvpg+r0t4pKGSTALiDLuHVYULMRLaunqnhv8y9JdJntdm2qUCJfoXexXS/oPJaiOc9zC04ary
g1gAizvX1Cgca9B7+KhzczkAqk8RHsJhj+ftP8RNfbKdXVZfH9ppPl+r43ePgtj/kBXec6WHQ2hV
RD/jBgQ3oHhoCjo9e3lFIBDHwEc4QitJwBFo8s21A8jdVsM0M/LCZjCAEB/rJucOZpQmAWiRuYR8
IjRGbZ1PZX1bioIcCJwZ2GfyD7M1hd8uuXMMXJdMhnotyum6p8KZDQRyMMmYmtd9EBMGuRpHLdz7
mlnhX1GEIzTlB+9/98nQE+nii0FLPAXN/H5NawEbSEmHam91vPTCd4rOLezt8Ou/Gtg0L2L1zjsO
CYfFV60qz24VZEjvswrHQHdeB9v4G0Q7czGD4oUjnZKaxloV8oZCVWH5amYX1Gz8dDsbDGruRr50
NVDWM5KVFT/zy19Jck3wHog1/5u3x6OXfkr7NA07lOkT7vvvkLvbkEy2cRiq2CJ89eBe2wgxsQpb
0YHBaBEKD2P2/i2sXVsZDbvtbKve1cpNPNSyr84hp0pz6DluCWUfJSp37wQbW+UUxqhA4WkOO7QZ
U4f5+Q4CvJkxdQfasE7hxIsQPzXSbWOipsrwJewIGVoyeDpeaWsjxUzf4jubTg4r+ldD8n29maBO
6mRS2yUJo4NCeeZgpcLZ7cdY7e0PSXpHM+xKofiJgWcZbuWHGQcSKjtOiKoPmbCK4Y9VhbdXdwZJ
KQRPcgebcBQKGM9jSERXa3N9YOaZCN2R+ActjQkvFLNczswP9l8jp5GyJvXALW4q2MMhbEDL+4TO
EUmMdSRzc2ACykHLOaNLtUj/wL+qI8N5N9ZAdpbcLzXTgs3rhs7FeWCBmQZIaThrWTl5KDzwvlDR
3smA7NQAGfps4HA2VNqdT9YN0sy/IaVBfblHI5jhrO8AdcHL42m5gRWtt1rZW755DKoZxKgCwd6c
vlH9ObsJoRfAU8VUSWW9XwnALxvEpZuqByQUizAsbJiOhbzHWbK2MG0jJpxZKh7/gq2FWgt69wir
R6dEPeBTg+B+orcsSaID8p9eg1vGgSdzO9Tt+h+TSLXVKHAEhJkC/UXL1B+Ap4+xsktwZnWd7IN2
5Zn76cOMxcH0cNn3Q94GWxf1UQgOtDbirsRvb6T84toGwunwIMypT19nEtvZ8U6iruBLrLSN4Mmx
mTtbxErd/ixsuSuC9Cf+0r/owdMhbVrJ7VRaHnljKH5DfIRaXso9SQR/TNLBJ66uAEBqh4lPQVM7
zONSWXoL/r8dLcRcwPWIprUQQITGudTH/rUqS7uIYkzmo4DBDSKUApbWQoaiFYr1S6U31/YLx0A4
wiQlUbYk4qRREMg23iQMaG0aDJ95QdOhPw1ymTl/hay4HcQX6KGk4yAW/BZ9nki3/6MzWOvLcaeP
u8Ao9Fh4g3sw6do6yQgqMnpvJEnIaIc/36vN24k/gTFdLklUcQC1vl7EgBJLNPFNH+fFrXkWpcAT
ySV9tAjLvSC/CZJiNb9G9mhN75TKXCCPk0oEZArZlErbixmPyZJfZmBGL/odei2Bu2hNYWxv/tyv
jh1FAq3//LHPTY/jIG5dFj3geq8lTvIv2cpfQASB4DA7mfunXeXS4j8ZOByeSQkeBB76pRMgLFyF
qQ2qoxx4xFXfW7D4JF5Dhp3GDF/9HsA5ZoOISbTtzrEzdqIAj9lrDPuEDYvk+nMruU+9LXo8uVbG
dd4POCnYEjZ4zsRLoR5ZCLJV/q224qsVEKoEtTzEjjOwCIxV1Tg9eVQ8Fv2jr1vPx+E4T5pC/qbf
KqutGaorNAUDfz1DfM43k9ZoZx6KpVwmAlBO98kT/k3nVB0/B07Xariv2X8hgOplWe27OaXs/3V+
FGQ8kk1t39MZA4h/UyE18f/hy/+ZC5OJGTmXjrX2H1fbNcDYcVRxZUIgFDcY3mRrsWj6FDDzi/My
bhkFhYv79IlXwB0N4dqim92YfMhfUWip2nxizFeTpVkHK8pFtHTU3S8LLTvNiGXreY11OMLiTJBL
ihPNCFfL2auzoE6YapVX4hlZ+N3taJFgzYlP9nL2c+ungE625wWezVHXX2YSf0aMeFnWgdsw5GUs
SUXENCNCT+tsUeV/42hHMNY073lxikal8ZWMzVt/0H+rpb6zex7mAqYwerWiHzobLh4xPdpVC8lO
Yx4nhFElWm/POcwHUxNaZaxsJSL+WSU2H+MdSG4QjQug/5TW/4gMhj4hELTCjqSgZEGuzyxrkxaC
e9ajkPI9qpwFv5hb21/f+ohFaGzhroea0DgvmHwLf+CS/wyELon8N2x9m65tL2K40QFEAeOcsenw
fYrdA9rLwdrLNIuH2kfg6J5khNgeSX0VagfP164Bk/O441lxd9HfunG9QsEVjom1yVCgf56rGbP8
AxgYmltLayLPp2JXWW2DkdZRhNLcJ6FUFnmuQtku0Ol7W0y4VUGrDBt06FyIwiBxmzjQ6aF+wd9u
mDjCAB8Uzwk9uOVeE7Fi/0wjTlIXR1cApVUIdn6sh8Y4F9Id14drkJV3oRuxK4gKrmpfaA/Nws/z
YM37d5vOB9e9uayiJwpyRibAR2B94Rw1IEfUAjL79ZCURFb1Qos9vDUf0h/kcNk32zRUdjF1/GGx
jwKc/udqc/AagUZECu/yBwis0dBUW0W9XKO/RZUWN8v5l5tm9GHQTSRkboyu2F7E8JD7bThFtEiH
5NUHQnBKf2KDs0ZNve+/wSU411Jlqi9e4fqem1CA4821bP3O/KS6kPWHylkfL5YCyPy3/rxkRvxr
BN2tTtxlt2NwsLIaGukcaQlG6u1vO5h7ryA0J/feC1I3ITcBrTLTlKJLE/qTpYH+acaIy44bDnHj
58Iv24K7jSP9xaHcdfZZTueYGiIgwIyHXcERfxU9xhTyuUtVz2QHzIRCzcj43Mgn7c0c0qWeup77
BskeLIm3vnx5hqlTqpw58zq98G96HcboFwhw/oCHvX56o/vQP3kdnFMpWZ4MWABNyAlW6hdxOebD
gAvM95aRCLYZYoNPdtalQV5XlW5GdlDcVXkS+4jUqZDL/aBYHFfk9VINjLvYkn8FViPgV2G3iUkb
wxt08qC3JW0Xuz9rz0Oj2hM9oNHxG5WKbeFe939xlCJBf32Y64Y5lVk32lIOy2+J4MSZsDUIkd9f
wEELovvFgU3etjQvHA7MDLW7sUNin29L9aGgP4vjPPHDXPMqQZfuxixKQxk70hH0jbD7Ljk8vZEr
JUkE4D3cFv11c9Nk97meS8xuNJPWeInF4hoZZ0V1tkQh8AaVTzv0GyupCY42uHb9HnlKTAlOCcwv
rU9ivkPUv4bCYda73TENB47lKXsigtvyuPkuXBQgQ6KDBcC7lnuH9/c7AneRPXfChbTKwMSqd6KR
1I9J3VXPYvkPGMAwxmiKOx8HfDzajUUNgAEEUNObKuManTqynVm+BCxQwegP41blhjIaL5bt0aoq
s1MdvNuzOBOsWhh/yfOvZBShbn0vYD5IkfHqq2Oz0Muvd6Vl+EtRla5qSk5x+HlorOjnSHiWZSFS
shA0QuBtny3LkJd7MYQhPMBwc3c8B3tvZO4DAw1td9oCv+c2NZ3SspIvsaGSlLUmw5/dSKQAFAK+
I5p9dAhOGmSpk6lskiBkx08oTlZQNZ9luGm5wP5Ys8lyGzPupAAz0yDrGnXeEEnudXhJjx2Z9zOo
YDtCc0BHafg3N/H2tDVrYYK8klBKL0c/2zX7jAYlFXfkJ4FumfKgwE58a3LdEaFnBNF+8ntwRs1v
XSaBceQy/cAX2UKUxRDMqtlsrufOVs9g0LOPsmASG17VSBmQox+Zy5GjokVtmK0+p4Jo88sXiSh/
khS7M5pU0SE+auST9iYBdt4JRBTbhuA6sIg/GBIyQvA9JX/F8Yb9O07robVj7mwuo96euYYhrFRa
qBbIrUkdK5FQdDc04t8OHMbOCBJOA+aFQWI9tPeIxae74WPX0EuQutvxyRTCUN6nrlGf4x6Gqzmk
kpVpQBqWZwgACYI69KBFLjLK3r1BkYkFap0V2OOAZsi+ippYMs26HIPPBF1MvCriFZTdK2B/beKy
qyyQHpGxkTghRShzmkoWS4mBg+QKNXUMM1ujhTySpyE8rHBE8qHZwKF2Hky+WfrJajj1OIY0kNoX
EoYHbc+W8kufY/isAOzybBZrSHp39H9fy/OmUk76RlxSD3oOqa1MIhmeC1Re7qwDHud/0lNlWraI
266gis4FG4mPl7EXQAJdysqekr4dI0z1c8L8KRUn5MSIgf7u3qnFAyroCYDOrrXlTLvmDYUQE4oB
G+KR74i+r/Qe8BILx3MC4pRSm4nCoCmZZJ0Yd3ez/LOsJ+EuLkGlzQJBaUWTFle68PriqWCFFvO8
yNZ17LtMfKF1j+WPFeXuooSI6+sKQPvwOaUOsjuHYrnHdwfOXlqltHO3mU9WCTOMz0rSlofbheiG
zIg3qa4JyODgSw4m0j208EvO67LD1IqLkqsF94Np8UoJ9k97+MCTfT128XJ6co1LT6Edlsof/5lZ
0BfH4K0BgOXEUEzZDMzhgg0XLmXwAGWTx1FLkhvQp9L6XEecmFuL7Noki6WmAPhCocs0appfrrzu
X6Qk/7becIUbXuTvdpTcRu/PHugHB/8zav+eSTYjhfXKLvS/szT/3BZgbek7qXG7yAdbLrammiJi
9kmdLTBwQweQBHHZhRh3Pcfd+OFc5Q9TqZulHWWAD1M+vL4Hj4B2jcGO/3LGsUfF7tcvp9QnI2hF
AI9/wSExGayKKDw2fq+rQgmpUd/Ky1/XUcGWRbL2EAqrQYvjZXnkarqAx1mU+5LHfEiCZ/AyzZuS
J6NUeBCdld8Ud+sr6F5JxT7V+kizmrcmDJ3a/+QPe02WFV6Vte2ezr+Ss27buGUEjMCTfYl2Q6B5
HArmxiA0Za85FT9BhwB3lHG5lA1NxBpJKqZ02DwMk+oNoQBiQ77fz/ZJTFU0vL0c62LFPNgcMhle
SGQlsyXNzkCebYDH8LY7tSP4IpTdUYRS4f8Vo4cuYv47/q4oumid1fvtj4uxbWs2mqBPj3MPv4IO
H5V7DuHwA8LEwHvM4NsYUF6QMNUKQhSTodoPaNQwWfT5ioSboldYC8k5qJgm1og+gPKjrti0mOSX
Xb6awrc3iVwfUl+WHDF4H/RUlrYkbu6ZxRGQjG3fT2xvzIHwn4pRueyCN4eujqxYA9mh8v/r+z2j
IsFZHVtTmLrcpv0poV7TyLYu5mE3/hkTJtkuKs3/LdmCvc5oA4lGgEhHv5itTZ3XwdVCd1LTFbMH
GfcB4YxGohDOaArljaFchxBR1VXueSKOFq/CBc2j2MRRYMpWyNPdwIOWJqwb6foV1U3HWrX+FyuY
RffHj1LaH45ZlanC15Dk9tCx+f8ZeDmINw3nNXZlBCDWcM5A6lWeQTEsvZ+9VE+PRlQretCCLb44
PVR8YtaAik357B7AvlRTm2ZO9z22c5/l0DH5SN/zkgQ6qRWBPVwXF5x3p+dp/rcnSED//x6PhBZs
Kf/xtQAbCedbjFYN0Upsnlvw9zoqhj8m2Zng0fB/XDQ299HXWzpIkWO+7HnnfGnPdh4dUkQ/umCT
xbmrl+nhvUt19/j/kJxRsmhvc5Ob7rJeLEVyfqVJLMwJ1VU6FcBVh38prjSVY+rmcADQ0XPkO0cZ
EPB1rKoendvdsbh19BjBy9JusLbrQsGtzYq9yGprCQCHBd+/moyDshHr4CbLXQiskJpurkkG648z
qIP5e/K29+faagfjQTwsnzITiljC6uDKkcA7y13JdIotu61Aa+C75narMKpcaYZqlyOw6h8Hqryw
rK5g1iRjg4IAhG9uOnvfZRxmWrtAJTbXODr6k7ZlTakjrYJhHf1g0glqg6L65hjB0zv3YM9rpvD3
lTpTuKbMERvheKhuPWcMTacfBw9fG1pZN1R1z8AHspvqmd1xPvtHFdCw2aa+c5OZ0i+CHEOWEnLj
ZzmSY+Q28462YJ9WXDNGfIG2QQPixnneMin8EX3iDuHhXz8qW3u+mOxZf1v5ylWNuSBds9B5mLpd
ZhqIROZCBvEXzKj3un94w2Q/DjuE9v1+FeGF8wIY9BzdLFR2kGp6TzgZpRbY1Omd/aY3pk8ShbfL
zUcsKHEPVcwMPoYhQIK7AolmD+ziXg0npghTq7AyXYXgmPK/BumPMVi3TcE03wmbifIQV+PZ7n1G
QKRVWGSBaoYE8NZTqpmQPmFOJLj0InWFUbbJ9p2d6Z0dGs2tZXgaMTGK7DThVdCl2a6rAlYRomke
nNvB4ristDLOIqqEawLDZk/FcfHOph97GQXgPnW7sxKeY7mArxYMSOVHLyB7KMoTNgU9JZk60iXR
D7+VCyV09eu8SFAlJbOoZQOdR72djcGcnbB3DMn+KVaJg4ffv4DpXyLu3d9/dEasfLHtgdesCgIr
KjJLe2r+iVUzzhrb48EoQwlAqnDs8N7Q60DLDgnKUl0fx9h9MjBb3d1Ft1CQakdJdXcm/ZtjiOKR
dzMWGW+pz2MbxgZAlAg/nOGV0P/U8cYjQJlUY85wxx56RL1ky93daWT6/g9d2zbMW1b6CROnhzFn
46+QcRsDFbJELlBL4xW+oTtozfQI3+bZq7NjUup7J2paxLFoEk9vrw4kZKpHymZMbtGH/lUdPbqd
jtckDLz5ZyLUcWp3UVT2Fy1xGwSrXaOsLE1Gy4X4nieMteAwy87xcrWjMOHdbjmtiCf8QFQG56y2
Kpj7aOdJaTFT+++RIk1kSoBBfD3hQjUduK00effotTwSeKWzNJexqR1LHSJLT0CxdMsda55UH0kc
K0fs2fz2g4Z97/pQqa5PKe7c7oWY0H9nyRaTrluWNXSAe+WacgDrafiOFzlGoxKFgdZAGRLwe15B
zsIUTQ6XFXSawFRxG59INQwEkINRON7tVdS85GFVGjzYqb+mm4CTmgfy1jF7I8OciAJQW3t3aVXM
kBXg0/076XYiVSkxjLqqzrBVgxQYYAuP4k2sXkzIPisDQC0lujlUB5eNFPIjb0e+fbIbcB5IWCQz
NaxkNRmchY0TG1zRskuMG6FUz71ZIuaTinz291jblwPDxIL4p1AAzZFrB4AxdGH2SOPSgvnH1jjm
6jKXCu90uwVb3c7KDWPozvS7nl14usHstYaZMBBf0f0r/o6WGqgnq1TGE3pkMkykEZdkq4Y0C4lr
0keoZpiJtc0+J2AjMXvM2lk7kkiz+/gPpNYuwJBaBeYAJ6DYKlEs6L7J9FYlWZs/D1tFjRn+YL1m
M1QWFOV1RIO07wL94XZAmmspbMXuhZS665qE4qFRRKB78NtSIL+pzp3IpZvSrIKLs9GsSctHmqtg
CylbCIglVunM39EwIuKPLWiVE4ixtmSf43MEImHqi/QJaxusK8owAFIjNJY1nE/WzmC7s/+VU2Nv
LVOavfoZ2HB3pXhHoF0D5utqwRZzOgzPMI4Rb8e/M/v1vVlhe2ssRGL11aEWTrh6S+J5rNDROFLn
msy1x/VedD2Lc+NZlL9C79P1J3+i9ePQVR43ytKQS/um6JI3y+mHj+5vO8AMVTWhE9AhnhFSUYuf
v68xSCgriH/ykdCrwBWywzMUOWOnh6D4g/ptmV/V6VJimCqakt9EoLPlU39w/UQHJ4OvvP1WjmNX
dX12g3tYSui70ttCXjM/UK1jt0lgk9ch+bqtlrZXD0d7LhL9qV6totdV0DGxH4eySPo2U2Ly33wm
QwoO6xYAxzZpTyoZT0LZuIFh9X2tZTX4YsSsCeFIseeLU7Z5+fvMg/mDy2Jb3P8wh/NhaK5W09vn
LU1QPQnz3kv9CiG+kZLS5X8O1zuuTlS1NWx34MGrcgfJfuZLADcKXhvVa1Q/x31BApOG6wGl5Xrw
1T2igw2hjz1qoEghfT/KmHNXFE10u0SdxOTtjbBgoMeoE1y9gwOrrORQXeeW1PJY2H/epiSF1O9r
o7W3QZMxz/5pkQzecrLqLHJE5njix6Inq9KK0wMr6PgrF6GQpLdEXtBuQO0VOJLWBXZF8N4yhU6R
PslydLjoBLANl24+6S7Utnq0IaP3h8euzEggLxUJ8Xos7Tad2Cjdfo0MmWGOyUOpGLcW59fcJ3MK
BoxTyQA0NcIRc3wg2tHpro1bgmS93XVwkBzqr4CvClVVU6l1QPrXA4OvRZswf3H5H8MIBXbmtjxA
+hsWgccHq5l9THI/Ykp0xgQGqFVSGzbKrs3dp2UkbNxdg2vPSMbqxfRoG4ysJ0TYFhMnKBohqte2
q71pVJ28aFOSohVKcdcu07ouYLKvDhGUEAvTGvektruYLiIxYOf1NlVX4bV4XncKrq5JkLr8iQWi
HrxFg9QBWPgHFy+S1fyU8HucSbjW91HcoIOBs2+nL5mTsigkLIwlrx/zOI6Nk8sKdg/GsnKP1LrQ
iKi1Fg+uEKiOLeqL03vIijr/bm+zFIHBLRs+oxuWtjg7QIBA9Gc3J21UryFpkqWdmiZX8vIJz3M1
Ypwq/LjUE4zG+ggpa7Ul176hqq31T+s9xQcc8479Sg1owFbTkF/tHIM35cUb6OctNsVGhznobGD3
cAfZA1S7ef9vmoSTi6W3/UhAcnvgGZnbGMGTuOclV6Wa9ovGvbpFro26yIls0x+8Ri3AzUaDz9GE
kLjEsdVs0pUkF3x5jzQOHxarNyWguFqP+CQeP8TA18SPUzcCwHcQuZw1GGWsNAt0B2+E1Jz2FpqZ
YmWuKtYw1X2k2+taglOFjNSDP95yuJX7G9ThZlw32MkrEh5PBbJp0ceYi6lsvDMi3xTWBpOXhe+j
9UlBcVMMKapsPfIMJGyEm0TqfF+bECmifYw2dys7vF7RT0K4XgKtxwcfxvO1Oo3UPhvdXXnz1mQL
glVtQLYVvd0NgYannhlmR89Y0GHPhch6PwnCgZMnfTZf8iZYgQTIk3E7VQHfqjqIZBEyQoPO4oy/
llCrkjui6+a0pzVz2yUeDbwxoDg2ydgzNZrBrvfWJ18yxcmkFaAyqT5PN3AwuK95DCy6CmmpGPLZ
Zkg/OBaCbEfDxqYyXfpnGRw6hOakEfEt+taMv6Y9rHz1jejz1vvPtHrrnU7NrrwrzhWbefOe9jVl
JdP/4yo3+ifqws0MKqYx8tvI92sUC0xXTvyj3pIPXztJwHDCoZVU8B3w59XhBda2of7PI2v1TGVA
N3e1ExuBakAMzye38ApuYzyQUGGj5fL2UenU/E/vFZjtgDxVV7Nhn8gDft9UfENieecgr4KjtDzU
WR/kAFwfC0gJEQ2lFLHv95ZgpFITkYN437yYHG09yQKtcKh4+34owbg7ockK4jLI9yCViFKnE3Bj
AZt7SVIepVFGS3+OwYDJNMsuALpWH02nGJnONIyM+nnG3bhYzHCZgjcHU1sPz1SquW2tVKe2sU45
ioPML2AvSnJVzbHcyAq1qkfywU7e9gbwH4WSexOOCZ8NPkO4mC8MYfR5oI1ofzQRJAvDVVRJCFG1
pjsHlyoQNFsk9Whf/1kR1sWvfFsDyMhELhCoYLEHpX7g9KACLfnS10KDwOlgSrj+EGFOCi4XhTBY
+kpnmYt2gZmhPPnsT0pzAptZs9tsemk6Rn0BqEMgwouqGf8RRR02IBPnSihVLLC2SqKnI8UZTaxH
vzR5FIXujfYA6kIib3PfOHG4cpNfM4iTYQwrYitN045I8L4eySa1hiCR4ObxVKUvUWEtmOS9Afzq
RNl5h4YJ8NitNiIa+L7H2jq7HtHhmz1MPEVYlYRsICCFJNOuHHEgKTy+r5ySuynwrVNfukIyx1tB
GRLTCxfz/3y0tPFindGvZwjjZN+hl/CoKSNeNLBS6DKTemqA7CG0JrGCsE78IbBsP3jy8REw5RF7
qdjd/BtGIyp/Iw+PabpCzzY1yjzdsoYpJs39ilu1kLd5FjsYLU3YGr5Pyjl5ycOIBv00IkzEBAyw
gMmEwHMZyv9w7SFq3ntYLAdLxKwFSbeTAOV2TLmRxLyUMEUNE6UTk/ZrLs9IVZXerXUDuhzEBF7W
kbF2TZXfaVDM7dZF0xs67yvlItIjYBHzixuqEUPhj1wvrrmcDJDrT39LTYDUxKGYupuUim3M+oFy
clNqiw1aNXkmovew5AmO5PZdYgEvWCRIDlPSc6L49ZMewJlmQbxmcTAJlOZNMNpoaW+v682YPHJS
lOEn69bAnoQkK9E4ytwXy1K0lXTChHEjxXZXcOBBQRJ+SRis5bL//XEYuBVkBO0AaTyjPynxMkHu
6dToHKUyWcxNg/lJ7sesIE+EZGaHUQYvLju7jszQ0EehdbmpbgiGjm07EGbpjOLsn4xlQPFv+osn
uxoeqNBUcsjgVrZBHK3kOp/zF9cfIuLJtX4BU/4Rw1lUls7eKbSeFSSWyrh+Lu0WpGBYUXtmvDvs
GuGyDlz1+3Hq1RTxBwBHDatd0/HXFZVLcrj+6mZauw+VXfMoAfUbAoABy+Z83KqRe4GvKRv97DhR
viyQg7P+0ZszdhvFddVBUfCHnkhcyiUOVSO8IikqOKPwpG/na27tbk9tYh1m0Mh2lIol4Bd7buwT
gHcbN/IrXqn8CN9ssY4Vh4cCeWny4sN3fs9P1U4eYTewmbbT+lfUQPZeHpqIDhEso4Wbm5bGnUkI
KSKJRoffG6/2XfgtR+OH7fNSQ6hZBtIILZaWazimwtjg7rVVggX6SSGn0LOK/mCgsYFYbgMygMyI
Bwv1UsSn9jr1sKP1T3bfcI93xuX1GZwGBEDH+ds8ina5CtQ3Dge3gUt9VdDg2Sz9SsJtt4xdQ+GI
R1/XeF7D0kRjIfXOIUlHLjPQ+DFEiwQCuWQLzBcR2dy74dtlNqXpCYmAWHoG7brUAOkHFvO77RtT
z/l7IsD5jejvQ8SiOruFW2528wGWNdMd/2DVrUdFoNHDV52zsWO22SMh32ep7eHk+9CjHQ1aCQxc
vKEONyYw89TUeizTLG8U9Q5pYjkQQeQY3OFwxCOP5ldYZYKO1LA16x8n+mBqQoYKfFl9cbGSEpl2
lj/8YRkkUryA31hvM4MAlcHBOM8ijVYNkzKgecZOkGVV9MtZp6pKHJ3fyy+Wo3QwmtmUAFLlTg1E
ts5UI6GVO+kRxw5BM793k7WNPPbrvsT1/Mbm7zEXfVsWzf0RbuT3nqijHL+33IZskWt2omGtlu9a
03Gj3f5m58MNnorSTpOM0pGu8ZFqvg2uqBSbPXyqerkWqhrxiMHr1VrRlaK5CCrkAb3ydBqX/Fbb
2oitlbYbE4GsMbgX4P9KbdGDiIE8dqVI0rZJ+nB49FFwOPxIjumv9jDB+cXqvzyGCHiWwL2vQEEY
w6rfnqEXpcxcVPiw2MoHC2yw7HLl/MTSgZpeRDX67Egm+Uoexzyb8unOisyozzvsVzHGr+WET1H+
NfhzsABlPLbAMQvfNycjA/pcobxvf3Ac+5di67/e/MTdUWmW+4dQf4Bv2e1dyI1/Ck5sQ+z2pVxB
Hr7LRG6WhyF35zyI0YZzKlIkp+AK9bp/kB9C64FOlzcxeSR9G+tA8gm1D18tx075LcX9xZ8V0IP6
qNEPzXQxTBEj4ZYh4qLB63BHDJa4PcA/1EA14B5x1doTy0dMbQax5w20AvZcUIzKj1Ac0opyuM2G
iLXtIuoDe42ipCw+YN8uZBw8hzUnilZORgWoXKM01QQYlzeYHDJKg7MMtNYBLberUDA80+dThrPj
XYAjXHK10044diUESpGfBde+11gBY5pLUCl4xft6wjBY877/9p3HUBGhlCW+5UdEG9cDmMua3L6S
I2Gq1tactBu67+9o855TIeIVfFVxRWK6oKQ7Bw9B1YDMnHMrStu/BO32zW+XcTwvSMiYULGCLSe2
M/+qaA+8fgdTCl8+79jRXQ4VkJuwZsHzvX4rB09skrRTujvR7wJPm5mzLODnH6Vy8ruVMhJj7Kr6
y489X2DC85iEITMGqH44f/zQgcOqNQpay+lCYJJWrhn032TLtK0VsAdLEGhBUnZ8w34q9hxzyLSG
4wrxQx2SsNc5pzQq8plinNt06ZbwfaKetxF8eYC67ijZJU4VoGHLYZH4UW4zU7TgPjFrT51GRxA7
p14Hx5Jak+tvAqKiTmhjUWLj8kf+oCeL3oECm7i2Qgp/m0Tik//E/o7rTExyqcLouz7FDGZl9iOd
50Gq7LDU8xQm6YLbhVzTF5sz5OerNQoRdutzQqEfU02UC49yaIVJefBNcBCBa4TdeJDHLLnCivhr
FR3F7as21+1rEAEqa8HBhl2GlHZScQTrBtXdAWFoUd2EMuFNO7E+GlRDSu4p2Wm4MZ9R6qS19Q2F
Z/yqsor66IZKnpP1UWjonTgCEbJ9SY7yQdMiSRdn1JyNfz/wl+htjHmLa86kt038BXiXf6GrS7Yh
ralXgyuUq3xFtnjUHAcKh+jf8ypUjClQZBkAPPfMPEe0VUL4eZKiKYCWqimODuA7qWNxPUl0cG4r
uflPFBYYkwXEZDPda6j4gGkA6HmOU65BplaEe7Vdns+DG1V05vZhhUPdkQ4WRS02lUOCWPMfe00Z
o2ILRqktJEOLkRNgP5ocTBDyOJmpcNu4Vz7Ec2fkwby3Pl0Em0p/QDfV1QvEJXF20Kq1KfYu5Jal
L0s+UXPBSHYFUC6e3Yl/aD01OaKi534MB8QfWOzAn8ZIEaQinO26uVFiN1Nf7iCvmnGRndY1fLOq
bEAZG2XhK6wJZBtywJ8HlOOYIwsbjGlbEyc=
`protect end_protected
