`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Jxuqb805KBajLEG0SJQr1II5Y5LHCPA8UL4Rq6IO632SdMNyHWwCOLxgV9LG/rD4HC+FIaE9r3v9
C0waQHn5Jg==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
CEe9jbpSNKFr2BUtOlsKpNBbrA8+vH5SJ2zCkF+eSPA0jxG+EOUN+i4w0XExqtY3NMFgFuwWLJXq
jGghBslulaSQsGixbChhHmaKVL5ekzuE3l32ZMYINhFFPRGTLn7gxkXU9PZnbSeue6AtM1/wsiHu
+rANp0kdR5qSPux6a9E=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
idtOAGocQhdkM1VwR5KO4DpXZCBxn3WjZpeRut9M+T0iEWqNa+jjUEo6Tr8IhV3i16+fv1qynMKK
KSsgIWpeR5SJf3bJdVBZGc2BcR0VjTSNAu7Md9bd1nCm53tx+8VeOxPBrxXCra1IS/7do7V+FtcC
HkZZypzmEBDSiK0G1sLLW7qj83QotyS5mq+l2+rYQ83mS8TtPwBJku31SOcIpc1F6YtP2+F/G7yc
m5IrSPY/mZgCA6eyrrMYriKnXv+oPQrNKv668bySdNH24YGLFYiplkyo75spyiYfpEl1FKiv1cC2
nBTN1PTJMdyjb/d9IQOdqPYAFyQEqNSCgQiGSQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
guDfG3LL22ImXg0zpQCG7SClIfhukDQYIHlOct/GlF1gFnSc2OlryRDWa8M77JGGn4AgmcSP251d
ziRYJcJFvamxxvsn870h1TG8MUqdJ9yeKyoFHZK2UeG6uEpVaJsyBMeksOyoNdB22Q44bUG3CZdd
XkPcjl+pGEUoPPq5OVh7yQ3Wo8UIMh97x/AfKFiKFjR1cMEdUHuj/s75oPXcNS38oXbvJxvqZvMI
1xBbUq4lU+nCfayD2DObHCt7idRYo3K6YX7BBVLILztou3dmwazcQO27EbZoCbCYtSU7mg6aQ3yh
n+gYSyQiSZvYx55SJ9uxH3MIQ0+2pL/rwhpvRA==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gNO9yFSe7fjJiaVn/nZoBAMWyekSWAhN+Ifm68BkJO6b8j9MBtsVk/nLFTQrJGo/O1TODejzEVY9
JMr7qHu1GbiawsgxfLlg2ZE7DfSo7lbLsMnEGTq0E0tzsC8zo4+UrwrUq4KJHrZXw0qBWJprSvYL
3DNvMRwBcBDs5YGoG69iS/JZLdSJWVwTkK15G2emmUI6HGOaDySzB44lHb7Bt1NZsSX9VcFAzu79
gsWmaTL7vspSiH86SvyDf0k3nfpjKvW6tuFRIQIj4pbr+CH8q9Ic83URM1Rd1mblVFkUQXqxAe+e
CLaLzjf3atgzADBMTABRZicJfoBPkZMp7bHMJw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XEST68kG3xftA1q66RUnxBsWBZBG/tOBaoodLPl9LMU3JkcPTxFhWeYlTskoonHKJOg0DBbryFZC
pGzHiBawznqAMt6iYU4gvntPaH18Nrur0FcIxTQg5AumK1+9srutGK8r1IbhC56ncssgLh8x1pWq
XhPuYlKm5Pk+m3WRLUY=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F2Xsr4DX5js1e8ivWV+fAxDcghqBR6N73XvL3yFiR1noxGJCWGFgQocIuaJuoHHLSxP2d8DVeomL
ADyaSLtSMD3eVplZD/HENDbWAYL7fPB2/m/yLbD4UAQ2l1s81is4u2qE2ell64+tgn08zA10KjjX
7I5SdHRjMtC7ysPx4FmZfMdgYo19rSoMWFM8yZTLwc/+LKrk4aWBgYoxawv1p7CyOtG4Rp3tG4DF
YCKmIm1yWS52hinJARA38F/UYs0YfkYARigtHdbu5gGiqgQBWC9yGGlKcFVtyGpr8P6nh+oPu6HD
6zjECprB75HrRgRkbjFlyjCUdv1SoTsZgeXl8Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64160)
`protect data_block
ENaU/7ZliRK2ASeKdgT+VyyguDD1XPo5AoCG3lZY81lE5/N9DhSn0kq3i1EFAP2pThnwHYnRcKDC
mIe+9jSmFSwXHY7lIL6+1oZz2sVhK5lKbmswrFlP4s1EaoGH0ykoPGGuGp4Z5iSkTC3UdKIAGCVW
XiOD4OPNgo/9DHUmB5hzQQus7Y1p8UGJ4OI+0BaMpjoJLltyiDflfAoCLLUdkiWm/TGB17MiVdPZ
+KZXL8Pw9lIWpD46o83hUUFMOav6oGWPoDPS/wbROrvwQB6X36qYsVP8u/u2yyzlgeWaoDJaeR13
TlUfz35wgxp+j3Gwr8pOnFGicAoVc+MaIsQ3YfgkPi3iEJDVYA1k9G/wDL0WZluJD7ck0O/kI9/0
+daBrphsoAyOWq+W1M7ZGBNDQdgsVuG/VSfTkWnETVO6PzBFIMQXll9x2eXBHfx28e17PKwM+wYJ
4spmRlFqYkV6bxLBa3FtREjY4VPslngu3P256oU6Ul9P5xyUnjlyVC2AGggXmeE+UdzgyN0t4cx2
iniKOwKMaz+i8mNucmj6ihuwkZ8cByhnIKl22i+e7UuPS3tqrwjobmtOaTU/qbDUcG6yCZUlxf3+
zaRdV1DcSXB2bScJVLcsWF6mbakgPLwOmC8F45GomTliBlzPghGqf6vBCVOE3lgjPzoci65WjY8K
Orb3B71Iiivhj4VzVmYBDZOY8S/w8bsfS44DUnLejIE4ADKtyPk20bzqdwBC0kREeiGoT6KOSA7Z
yVPVkp5hVttLsSj8aM0TolkSCnq3N/RNhiAJHYqAgyb1BA7/sYio+KrOcHDtY9Ri4sf8rTTfmwRH
nxnQoym2X4nOoKUUuQs0AgyBXP/IF5N+dKeWvbzOLaz7EGZ2yp8rswgh2fp2B68ihGlw4GlZp9PL
6zmTZp+jCOljmvT3Z9WnAhJjN15fDHqJej2S9boBDsK+tHwVKmkbmC+gtBc5ZkC8h2Po2/rBnPca
nOjRlChfVonbRVv+LRfll3keN3jMWgNC9kXZ+eBC3NYtiLFlmg9zd71WnV9cTAWw0XhI5nh4xeYA
q5PeQcGy16P2kKL5+j38uCn0uZ7oITpj3zac33m0YH461z12q+0F6a9FdUs6wGJzunwjqU48XNG0
gWcPykp/b2nLVz6kzyoIS+i2lIJUjXmkK6Ur+nKUa8z2OMwGLVs2lAOG5gVTXs4Xos/EJxxuDwQ7
6llOnXpQwQfndJwLMrGdhPEHGzyRB3WDtiDKrwB24YkI+Xr8enBAlDnv4/udwTDsymkAjQEZHlhx
RfvrFJI3Vh9peXmOUctzzmhJ9XeaW4PCBPmH8v9ebtx7dVrxpTcMIHAz1Wi92dR4aUvW889AMjuf
L8HMgCedpCKgPGjojEDsjFLTlCV9K6vCPrJWMQdKUAlclAMGXL9VAbutjb8y0awYCFzHX5VDDv8d
/o9pzQOcFWnPp3SctjjeMfZv3MsgaHLYNJfItYhtGZd42Z/hf+2rTB2PElHWoOlvpp+i6V4jQIxX
T+0ZIJ4oxfWjiI/GBCee4zvIuC4c8g0DRh0dSRP9w/dIEi2qEjSMqbC8tCCG/TzovrO40AG61hjn
NV8gkLhWIb6/Xn8gIg86LR6mf9cHud+jywXBhGH/DLEz4HujBM17reMo/RD98m73+tGrrBd3S6nP
GoXS7XyiGV9F8x8CNmO0Ouy9OPaG6K3iZvWrrsTcpC2IX2QYdg3q0hspXkAPPQzZLrDXTUA0K6gC
NpI8NlOYFFRsimU9FCizE3wFQfxZfh/aJfs4iGGGfTG0ebbrQHehWSpllxsJ32cKrzjoCMyMQO8k
ySUeRYuvyXzOVdrRa54ZciefdO0/JgRd/oyB4B59wv2EEXlTxJWjcyEMP+tAuIQnTaFnXL7ezjD0
aJUZthSohHQrJOogzut+KXD/nW5ETUXMNncDE4SNlSLSFp7pyoCjWYKmlkI9UMlRxPwkxF6S1lym
dWv2NVHPjU2ZToM/qIeaGB0XsNuxbL3lc93tv1wmehFX0V12O9dk+PHZbPu9Qd2paVRoF2WvXhgs
HdomOGj2IuLCPoCNRTtJtLT0pY3guetWaiUsFeDQIZ+xLV4vvS5Vuq+UcdGraAVTyAUdWuGqoCCe
IoVbsXJRzYFmDSdvz0sUDBWWTaEE6kDO8oaqZyXv1IifEwNhSGFspZRkf8Vr2YnskqnJ5kS+/hKB
LwVpeSoKU9EYcZeEkKAivfLAvgxeEdudH1xISK4jKZ2Zmw+TRXuHyE6iwxxeNnS9s7+3h+PsAl1e
Ggcqwd7E0HpwDlmFpB7r9drHfTasRtEY2W8+oOhiT2TnGDyqa7yLb7LwrCb4ZyBTUMlQYSBjHRuT
fqYJGQf+nuXmuwiWiUrdnwBEVYlgos2aoA2bwRG0BBbNK1FVvyWza2XLXchVoBswNiwHOhErsgpq
1G9gBxEIbeBrp5co1TdiElSqjbx8L/K9Vu61e36QHRTQWd5XzXcyV3a7ze0O6qx7D6/Zf9amTOTg
UlFylZv/X0N+NeGSbd2Vu8IsE3RTxxA2SAzGi2iyO5APuFItk3KKlXrcxqLPvtRtfL1b9IVSgPKE
Q3etQCY+/x1G29/BSEjDsf128Ou1ziICqDcA5bqe51M61LecOMLMmDQiRs0goySf/F58LnrGjcG5
z9FKy3EMlKTvbVeNPo6UDvB55malJu+RIFfrNbJVWDM37d0zVQNPL8p3OIGPgKE7LVTRBlmpjplo
u+GbFL3+2sA7C2NBnXDsQehASQ+ZdtHZUu0E/IkcBtyRnUXSMtbhMweagIu1YE1oTCV38to9e6IE
t0739URppYPTQk5/bq+V4KVR+8+HuKOCS7xON+CqnpmaWkZm028Iz5JV1OzGCsaPMGDo/lqQ9Boq
FjLCDenQs7OL9Gj04TealFt76DQ4fYu6/ZvNhapMzDSquNsU3diyfKuNXa7yqOlsHXdexj9hBXbq
UORG+CXqW87r9rzkdbwLIAXiDVsg6U4uTVjyGrrj3/1x5mX06+aXBNl6lTqRXnoo6A6RZzNioMZP
WkzNC9TvHNL9WmwmDQb4wGHiMFzgphwQ1Fjg6Q8DTvueTHGjqE8TwvBfFxebYlmdtNkczsoDbBn0
PtPrh3Me05oFCo1lW2yarWO/RN0xtKiPCmfoHpaUFqJPu04H2N8C8y8+pfCo4zYsp0ralPAowPcx
tAs0e417SOUxAySweFhoBIJdhqiSnFeCJ9Cw7iAAld2edog9rYA2RkkXmdMBU9eVSaEGDbZ1yIOV
ZHY5IysnIVgR/TkTCGfC0USqk3K+fje7pf8RK43xnfRTPTfZr02SfLFL7JYq+srHNRtKkCo7Xj7K
NfiB3/9CYR9UUhL+qpDEtE5zfa9in5jr+O/k0zn2dcXpxsQBYFraSewvhtS7gB4FYt3njSJc9Yim
avze0Lwj7QWAlmHxo5Q1LOZRKryY57rfvuWJLxzfPK51aITlhSzDV3vH6RKl3Z36Q13ehVuPtPY+
PO3XNuchxNFlEXc8g6b/SLW//vC9O2Y7nlyHhhvhWcx/KYgb66z+cn4mnKU6oFUpZZ5teK0tz5yh
UL9ZU1EouOZObxjhKbE3z8IORGGJqLYV4jiNBskEi3tjJQg+KsMCz0nqcM/IV+Y9jZE3TQcwNm3j
iVGis69D4XY9GQyk6c9HArq2HTlPy/rxxvuYrrXg1nlV8/8wF/Cfyf+ZaM4MHn8DWm6MzJ1SV+AW
2T3xA3uo8Rm7OhqclCkx1huJh8KwA71VA2kpb/Ryat8+326/VryBVzBcO5KtLztofjEgQ+j2RSb5
P6gQZR0TdfHFjniYBNYFQrg7BUC/6vH9J8cAlElSQiFHWnXNAFIo4l8rXVtK+SKTbB6ByrybYiNQ
tv+0eexOu2bbdMUD4A1Ff9BfAytrFkZOkAJwznYDXUijiGWBOIhar67VDZr0DJkcMpX5sKFovM1+
iOjJ3sTL8JjiXHHtgV0yFzVX98roLbmxGxMcYWRG0S+Ed1Xn0fCpKFv1aaRn70RGlq530VNVJPkc
D59yn0jSIz1g3+IxTERoKGHOM7Eu6Ydlwuy69wxXI0A4+mm+a4f3OYMMqgiSDP3pgJ9Kh31zVRo7
F0x14eoZDH5Wse7HsH7QxisnSJ65u5SPO5xuNDss6HLkqkwSfhgXITx0TpxKcBX2GWaZz31ftwdY
5mnLj6c4VEm7Ime1WYl+iOJ3VqWZtLWJl7xQGbVHTe52DTp9nfJWuh3Un6IMgZqDMqvhx9YdUXqj
WNFD8/Mb7WWZZjoz27gNmQZ1UJm795moVIkurOxMI9phCMCY2kLyb1dochXnYVRurplcGcEfG54T
N/DJCc9YXRvFz9oT3eZTL05DyEziUXNcvN571heqVFT9+42yzQXDRVacJ59Jv0n0Rd7L3pHWT8uy
MuDoMG199BkZ2F6Z+IKxEV+fLvV33Dr7AoS1iAAOobFQSTDTsZGvVFPsbzJrRQVUilDo5ajNdf8e
oQPNW5MM7Em8ahzXMqhmoBWonisALzI7/b9e67rYNX2XLjvSgK5LHCNg8/hx2YiRo1UiJRc0gwzY
KXfILFGgobvkHKABJj0nS49OfxBRs2NDxIHwk86bhII9z2K8LXX9c1xQLdgqHYq5i9UEpuASEDnE
VgJWc1BpNYVS6RInb0EQ1GF42F91YKb54ClOhGfrTq5e0U1K34PluzWSaQIFuyLssKT0FFgVKDz6
cV2mQ/F8uZQE/ZJnYdEePWT1ST30eC9U1wW0rMw9eHbU8NrxkVHD9Vn1i68BhMGNvGgQxzwkTMcy
74zfcwJLatgyR0Q4BNT/Xi15XPGeHqHNCxc5WlpIYx/eivkwedhyqLf/STvlSAbBXjoM7er82swY
IdN06oebe1DBnar2oEOrY32daBTSw1rIuI9wpMVfMEtzRNoNY/VC2jsuegzCKBNFygdympG97f3M
sMSmPvt0A8NFJV0oQbbRle214JhpUONRgljpQ225vRSPaVyeyh8BnBewwvpqUowtT+Vq6sWLtBU5
9WDvKkHjmMoLJFxfnim6nxV7W6rKA5wiGkHXBhF11kMRWsCVvWHIjTnL86xLc7WXf7RrL3GcRCWO
XAj51V5J06iKicTUy7nwSB4XWxq3ZdZ8y9mR8/9j27p/qpEdtqvycnzgP5z2fMs9pFyx+frN9DNC
lkdchOr2w+e73NFNNzqIp2oJEV3FURVK1NYQUKJc/u+wcXY9MOsFUTqPIBBuWmroBnj8BfvqbCDJ
T1uFiFUhqUcC82wGZzgvNfHzUnJWdL68a/AF57M8DqoxQa4A8Faksa3nN/+2ZUmuWWHPBvZSkU3X
Tj1XvUk9WPghXK9BXTnD7jMWdzWEL6xzbqwpeBqiPzTkldVhNqXCL2yJVrZjbLNb7eInA3X9zalI
/WHkDGHcd+7fKEFvHFdiHLTK4r79kO5UjhPCgaJR7lXSXrF9qLHJmGlSOZLrPEgQ3ZQ+INy6oFU1
WSmuhsOoopgFveb+DtBzq86ZYohrzq2JLZzn6y+0AE0VSh3weFyW2QwHnBCzbS4BIUG6zXkpNQKp
daKwOb7xV+ePWR3FlCsxYMV6RRsWi+7Mvqb4obibJ+wXmBhb61eXp4Yt2wxBRmtU8E+/B62N3qdp
98VetB4fmnIGLZ5BNNRHUt68wZCkC3z1NLphDqNp6jfedy0JAh7d0YvqGTRzE95zSwSM0L4GpZzc
k0Q9epLBKvnDCn/5p5gQkvIzGP5m+lBsl4Wnad3yjjjndZvNuEEGhELWnPnowIupKIV6uJLZcF44
mywFx6PDiI6ipdpqWe4xLfwRTkMfYmGpsdetf5RqjkHM65fa3nC+rDWAiiDK0OPcOquTHRAVGT0S
I1Y/NL9WN69HcATzfq6hfYjuauZZF+s/SpFEMqkobF6uTxOV9iz92ZIgbrblpYJ/+wI8pgxWjQdR
Fb9EPpBYJd1ezuCCKf2fqPWRWVm7E26p+tn10osJLtRMa7JMdNHIqEVqayAI/dJlcxujezLLuTx2
y3l3NgHJNHhfXCN+B19scUU2k5xN6ih563eHBQwSwTpzy7HjJ0DDOockFG5le4b9/5lOQavWPDDq
40uJFPpXcIK4pz2Ba3LpNwnhbI7N0UJLrbQDht+o/apcuXbKzjQ/xXwjXMC40tGHP3aKD7W9dCbD
R82xWuJsZ32jng+IpQvzDqbhrBou6GmorAZQGyImWBwNK9CIu2tT8D/1YHI1M2iFot3epeTR1Lwr
8VMM2JqPQ0GVH6PwIKMspCuRmxW4+QX8hPjcH2nxHEpEXgHqj5c02s3/ffCUl246i08HRJPUqMfE
IKvz8LH1JG6Emhf5QcPYGl/JJAsWQemWEo8JeKszP75EpAt+VswsIRyLnmyUnmC8QBvji0fx/TYm
M6ZUPEMSpPTHP3NtLCV3p+vY2D5xR3IXggvDjH/iiQvXW+jn/UP8OPJw3hVRYkC5aNqQvV9fMmD1
tfGQDZ3JKCRYJqgBnK6O8v/T1J1RigvA+BwJSI5DGqYvHvby+kC92eMRiLbdqeA0mGLy6f0/XspJ
ELZgZI2zDnRSWgShcyEf7wIurcxp/uktgmnWwR3OYU9U0eCBqSfbLi3bnPqogr29tLtjgQJQ5BEW
HWs20p8Tsuwh6RjJUz/GUf3z5hASxrjNcVxhQtWJwzJDs5AD3s/7wN75afOoeguN9yrwhyTp8aSn
+gGBlMFDEU/47dbgaHLE/oeSE2A83gtEtCRfxZzCoaG/uM8heXqmILHP4m0LVnKXhDNtS0sc59Cj
bXj26LREgPXBSELxWuWJOq57cmt2B2FaBAkGH/T8+zmxWjLwi5BcJO9FBR5AGdpnelanKrQUrrAF
cPHIj6IH1bhZRDdY5wSnSJ1kRgF6ef4R7b3AJEjqDAYSIq4zszLIU6PDzC42LatgTq1CMejtBjZO
5vULywEm7lG7IFh47HgZUSbwIoRPj5k5du9SMjbEKAXx6FPiTKL/PiCk4opoiNhn4+uNIvVuykSA
7gNrnEjxs07BgDP7g2UxmmVnAxQAnHVbYlzTzyvDIiTMQwBWD4ALSI64BAilIs+InMBpyGdU25QI
MJ2uiZr8EowGsVyoUcH3pOs2x+J3ahmsHlAcM0R8L8mN3lQ4KohD9sHJ7C2xkTKCh86gCU2vUUq5
KlMFmmlSElZgPMB/Cj9kFDJUv7dHGqGrw/bVNTYSqCInRC+u5xlOIo/42pkqgsPROoLC4wIH0RRW
99+sw+1ZjRk86/NM91VI8GF+VIBQVghEv3/T1IIj737v4fFxhD4xBsSWiutnP1i+WKJFgNYBSYFc
GPRT1UAymoWVJzDK08i4da8PmXNoQA6W1nT5mFdvZx9uvr7dEyI/KXn8c63Q2ONfrWrZ9cwX1Y47
/zBNn9eiaBNg8tcbcRodKQnOVl4HIKHOeWZTc8VsWw/o+9I4kq1O1HaNRqGElGzZJAANsq3fab0F
i41oorCgtLcpEl7RWQntUpJ5luLsEwr3sdOtBSyl7QWJivp/QT2reJhZ5JfEOWVBbBQPt1EiUM3x
gEqwJJ/FwM49tsLrxKLcyQMENIUwLzqDI8nT9IJPR3TjoSynqqU5Wa64L+Rz8000b65VZ/KfF9Dd
0/48uXcmvSbpzptYIXsXjZiasxei48sC8qWu2cOR1Sp8n3bq9SVbiRtJ0EcA7UZU8tYhVX/hkiyC
VBDHJUKWeyCxg1IRAV712j7FXJQp2Pts0rxvZc8dTB0ytZ4dAhbiiyn6o9AStnthMjj/5edzXyp5
olO3LbtcTrsOKZUu3P768/ZHIHUAsLl0/5kTj1pAfTym5hkEtefS1Fp74jYOIt4WDI4nXb0X1hi2
npJiQ0AY/T32MVyf9cl69XQeZd6FNDPLcs+Kmuq4m+IlMnFtJq90zT6cscK7mmvR2L6rWHnGY2Zt
RLB4aAVh2aixBSbvm/YyabrXBOzMEo4jIwnwUIbDuLRlTIMGFPYvjJCjpFyyLFH9PYOQFDwqm9Hc
ypX+iDJF/I+1lUxtIHED5wShaSsGoGv/VPxFQZYU2EdOGc0smvtU79UkZyiNjHKM7o3Q8+NDqBvk
Fy+J4D20REULq4vh9nG/53uW62dAw/8wnEgwypdLHbdIZsEk4AlE9kr0Xpkgeu2qMi6wZm/dCb3q
Z8HyY5AIq1pKbk4vg4XXXpWaI5xMkpqWtqoip9wmWrUlj4emZ893FICZagq9kIvO5VnuHs8fRjr1
JOH5j1gveQ/iQXsRk9D1y7CxdG9ANkq+QCBqxfdXsQM59s5o8VARoGAy1zpp3uNamzSRZGTFhYHE
unAswqKnHNXzp2Yzw9XxV7tT1ldkxEo4YE1SJ3nww0e313clro8fr93qG7GPrJng/vgvpolVLVrY
oLsJ1ui2WnjhyNrdzeIrJn5rAxcNr/tQrn0n4CGgl6jQXMb3Cju7qC72C1FoJV3joN2ugmw70cJj
qaauzoDGc/orDYvb1K4JHrx1pj+aXuwx0borrDvGutQALgfoq2PyMmg1ESHpHyC5GOkMCaF7maIB
qe9x/MzKBytQAOHia/zvhZeX6Cm9mnQEq3itfi/ZkxuajBGzOWUqLk3XNu1a2H2pCppx+R3ridXt
/h1rQ2STq/dNqFE2WpYzXuAiPjR2HG6wJqm5mb1Z3jWyFRHdAfSXUKKVgFrR1WleLWNKWdJadsn5
BjzWZSCwQ5qKj+lRMeGUjeA9J17iMy5/5hCoLMlOkvWGO1NY+ylGjfXxC9rwrx3KxZwLfYnhM9tB
Uv7/BYPw2v6fw/BhX39+4YDBXSQG5xM2jToIsQcsDNLu1ke59H0lpPY5hRsnudIlMSC05z4JetDG
2yvpnkIMPg3BUk3eqIVKw7yHPLD+Je7N4H8Wi99SSYtN6FroJcuOb/st4n9cGyzyVWoegsLlTceV
3xYiu2aVJfZ1WRIhe6AjxOsPB0DQnKB95uVpxp6tD9rt8/rxI9TDh4BLT/dP9TgDeBanb/afKT0m
sLr6Zi8Rj7hByV6unBhF/SUL4iCgOS92jaj1L0cW8475wM/z3s20/Ogk82JRJzNF27ueq0oLVcxc
KnNuto8wV0s1N2zE8+1aoFV71fPGdijkAO+I5QOHctR3Qu6lLdLTwA61k0/xtDQzb+VOgGI3eZPr
iylRbFjnH6topxXWTDrgIxjktEUFYWD+FBm8tmoQ4scEjZO/9x6o6KFzoekciSBweBzmyYvIKKg9
0y8BXt0EGMcs3VhrEMHckJiEBtl7ovnca61En7awsj40j58AixWO+tomzob0IZbMLZaYDdcvOJXT
fsk8dYBdKq/OzZsbwe1Mcpa+nHtyBuDjpnVvbbVxNihzl2Qxkje03uXQ5w0yL/WZ2grs8K9mhHF2
LlbzuKE61ImYVR4a+tDL4mf4dN86kR4+wlop6G/yE+ED4ihK7q7/NLMQha7YH50OKcJJ5M55TvTF
atkPjnW2+S5CmgukIRF7nFLOlmrFdTBVCTP7iP1ADbbw/SNTy5ML/N3eNcb3G8tIgi3Z+zdKUhjE
oooG5eHhKIUJcd+ehpWrIqbXd18WkYTsMrEN6qKr+r4TLPC5KafvW8t0I9mDL0EcXRtl8mS0p5ke
fpPg5cLQi8V/lgN/y2ciWTse11G6v18xW7b0UVkK3feOv581eZT+eg04BzmsD6aouLicbTs8qgRX
Dt27yTpa5PU4aayUR+SyoPYZPh5SgYyT3V92f2Qz79A8Gew57y2n3uARvwittny45cbIZ+u77SbD
pfcxvh+26aepbHVVtAENqOUJhIZz++rY6h/P3+Gm2gZcnvxbH10TTSjx13YQc+gi1pVHLaGEs6fB
bM0ACNWkq4PAAh0MO35ENmtgiZ6kG9otIntqAOIc9syrd+oTE1xMAIiONpf0AAktnqsEEl6j2WEi
JyLPojVNdKk1pjXxI8AL3uzEtJ+/fZ+4xEBApzmiCkDg7U31880Wnq0ZX7dgeENSt+KKPZ11fTji
dXo1JDO7eKSPRaIRfy3SN6o6xnI/JJgAExJR4cMJ7QCnuYj+7bjtlu5HEvZ43XppFZfOqZN38uLa
yG+GYwcview5F5Zuqx7Me2XEFGWZAB3Ylp+dH/JIkXVoTd83oSgH41CbSGRDt5ddO/2R2aY2HRuc
fKHSXpQyb4cwt0NMSl087TfXMY3FbfNdTKpaSKhMuQcqTpYRPXfcJsG1xFM4KR8C/5CTmpyhsgyH
mIAbHj8aWsshupaFrto5og8ESARcJSn1uM0OH9ifkNtkDrLJ4OGD7ApVND3v0CJMlQHBbauPDl9D
nlk+H8OBouEcYPhiczxxToi/Op17MhRqdPa6kULo2Hnn7xTIA0yFJJSKMM4gn0N8FwCgXtiuNjBJ
97VNBxy4bSmmdiyMII0bgvHs/8uUmQTVNVfv6jImu0PKwKWc/ZXXOTAtXxaeTuBqDRP13Z3+goGm
c/VSrSBoqDNeF0ocE86YoJ1JTWlMHQCmeaUz0ef79D98QZ7bmy9/EQM7+xkLtABYQn/+V5AGjbyv
rYaIa9yJ1q5rzpSa0OF7QzJFDtJ+VVH90FVBO8n9sQo0+3aRGSzByZJGIfj6uvzLNpmFEvtjVk0D
kjGGwUSZtzS5nIeScH2zu7Xw1T6CeFsIXnQmD1g6BzxWtTL7ti9e23SgIXT4Go3eczuDPTjE7/hK
2KheJ2QcbZkMCCFKN+wgNS0FJXpqNvnXZOoSKP0eDlW6WzV/3t5IwvJU8bHvdGakGQbJ8sxFtp2w
mjp6rO9DdblsxBUZ/z91ouPFgxzeKzqaBmRTezlM1VGVuHfExgnE36u4p/1OJQv99m0S/9szLwrf
49QMT7Mc2CRcE4LTcRG65ozHsMJz8IYywvOCsRO2EuTDRjFC+QK8fUhYI+xyhqnCxt8Cg3HluKLQ
erhcn2UBGO0jnNHPsWR1TxP+Dr0yw9ZRbZADacdppFkoI6J2/D2PR9bUxt4Ldxsi+KupbWaPAdNP
D/Tf30gcojpeJ3Xd73+Yn+Czd4KxJR++76zOmVbGUvRRRCR14s+hEopeKR3ZBRYgtZOSf28XI+97
w6DjgF4Ks4nMF0NpdgHr4fMaLqSEuz7aM3L7IslsECszwz/bWuhx5vaNiBPn4UtPMot1ZeM7IoiH
8pFdcO/d7wGx04+YIPLSX0MixQzYAO0HjEN71k8eJN7TzIVcXR0l2MeIHwbnnI3a4h79MmaGzcXW
Cc2XHIhFYNK1tUPM9sx4Ox9XDJcJn/9zjsz1C9Q2euNwxPpvnmPtS7RlTx1AACEXk/CviOlv6e8g
3nLtN7MLTzwz5Z5RLCGdXPdV/7CI10vlTJfeFdqkewHFfJajQVoiSHcXlDnGFURxl039Wlt+Mf9k
aplfw/XEC/KL22jVKWxFqvePOMNy0y7l8goPOjYQZ8TKvpSh79ENgetmYIYv/e9OrJYwLKL/Qtv6
y7kB/ItMvDs3154fg2asz7ogQxGkxoqYntk3Ve8vQNc8QicfePqo+Zgv37vnYGDcvmRZ/bFoS8AO
68BZAaJUzjvmjRKIGvaJenX79Z3+dvPUu4G07ntuhPk7/bryoGhNZBGYaBjW/N+RyhVYl9LSsA6U
kfy2DIB1jHrZqcV2UsFkQeU+ME17qxmUa76MMyFIVld8jOclqWHX1HopbddNPGEuELs3uP1nmIdq
hJJi65UI8UIPNH3JXzOIkZxV1Iadj3UoPbO/lMow2BfhTdrgyx4ZlEsVu3ZDsTJmh+MUvkZFVBGn
DOMlV1GRX5J8QUcmEzxOfeTE0MiMFXuEs4ZRt6+NOUbNCCzNyMh2QfrXVaSXtg++hp7o4qQ2oE7o
dErYMk3Kg6XQsW1VmF4/nToZa+FgJfMfLsCYp6qZfklemMhi5LabuIdFqEVDS4mx7yjpD6MltRg1
1poAxs8vMEIYuRxHPbOF6OlViKzR3atc/FbMHesVpWjezje1OSNbZgnuwjg2BuNwyFooSh3OvTAM
P8PDB0eGttc/2zwAam6mlAOkMyzrMI5OFUOW1nWZ8eyT74KGVLsItJLr7ptHa+4ATY8jNMN2kGbI
tBfcGihMTB9R0U4OVHSCc7Su9FFp/3D37zZU62LYUWs7Y9Dl3T8fdTvGpAsQsfx0KZYOUsj5LFeH
z2zqGuyv2ULCY0zUEj0M3ZELvYrVFAHQh5W+1K+EDroN20VLllMVGxklQxthmEnA3k9taBjr1vmO
Vix+Nuo1q+QEy66GV4y4X/v26g82BSMXvacPEiacJyuPCe1K+9Aql/561SbN9oNpfFqxRFbLZe1Z
nNzDVDOEAcFehCE5YH0SKk4YQA5gwNsuRRF/Nzvuh4x6SjtmTbc3IJATKjIKYT4IuHPbHkU4PgvM
JMJcWS5Y49QEvNC2EYhaSf2HBjq2tCm1BfWwaOBd70fSWZJQ4z8Msgo8u+f0JpdJnTnzrRCHoufS
yr2LjAHsMQXlcaVdgqhHvxSUqT4pvO2grLRQFYpZtschMz6JXxwsXpN2pXYjjifL4RRSVLcBmdTh
VkGAi4iV4AHcEsA6wj1wT3TTlsvQJTNW1hCsGNObmE/QbnekWjAbpMARtwhWrA91YZYirwQzhxDw
IIVX96mSjGA8BjfyC/SMEl0flz50rf+97x/uYVh3MDlLUsJhvA5Wkbbumfk4P+4s/1sTFx01ejRl
IFAyPDQawzI4FMswm0teVKQx256lUGPmbZpxpcCuaAhohBxJIhwCJB7rCeT+MpIsX37j0n/ZG+iW
dx8f+PgmktWJ+Iy6n6DteE/5ZkeW3Chgx03yFTHxB11OeqpZdJDztFLfQwh3/jcbYEMBc2NHRvzB
lGPqcVEkHm3/bz7eQ7YZkcHhOK19CyzH3ID6Z11poJmU/ICpn7jP4O5mcsX3cl5zLvlA4YdAALQM
bcRWKdJZ/+9mwgvL4vVLy6GOnkCooMTp9JQSmkDp/1Ye7eQRi2eYON7ZDpm4KU0u98ZAJW0jz2Dh
xP6VKCyj6uUGJcl+Ee2BmyU5oCDYpo++OZhZolPFtThxQVjKXIZS/GecJlnksJVC4ja/ggNbFlNM
g1VABY2QCe2fgGnqTFJhCDIefJucdFZnUKq4O/rnkOf1I4Aplitw29NsSsQ6U5sADAa6+hY4uenA
rGwLlkE0aJCZlYrre1eLCprBFZSuNT5vrthVIlE+LbvYRFijYaEo+HIhdWsajoYWrcQDO3W5op29
fQgVPuWGobxeJh/r4xZOjJc8PrltrTDoKmp46GXf36f6Y6O8ZngYr4QJFNiG79QFsFpACGvbupr4
uRHe3nQu/seskqxtjRpLHJNqKVmL/y+t8+yIqmEOPZVlIWL7EmWKHe4+DWgFM7JL73vrIcqv1m77
NBPBkZsnd30c46eYvkvJ8UFqCF/VSm6jOiyLEtMqdsPENrGU2Uwsh3wMufCXzvdfrb7/G6Ez2AW3
aojSqoRYPtN4K/2TgjB54iWEYHgo8et81faQ83KcBlV+QwMEsbJ0E7MMvIE6l3hASLyUr0L5fIkm
su+eBwlVlvyFF6qFW36zctuRX2yAN49mDVAG+N4V0ALcqilT7nc+MHkjqjx/GrA1Di4g38UAMsZl
IV6P45Q4wdk2JX7VHvxXFKCXs2GN1AIPD5dms8wQvUpVLhR0KOFogtWAVqWj3yLwGp5CCUx0PjCA
ad824ErhtZmazfCiRfbNXawDFfLNXItEiy9zPRJLj3cc+1+JAs2ohNb/vXQuRbDPtVbgW/yfyHKW
hI+97eeIakt8urKwxdjx46/97RwstCcxIe212PFkvMmPHI3JaoqaFErZsVfBLdo+lQ7anxEbtE2R
XFvRl95mZ/anm1h7Tz0C6OCGOaM2ThQ65PAS+5HrHFMppGWh1mhtKYqvRIt9GtkTbZR03dPX7K3C
tglsyyC9ilB7Bj/jKmzQeQ05KIbDIhP7lLgp0dUz0BFOLEYMB7gVA3HEhFK1kllK5cIQW5y0JlnQ
Z4/vp3eX1tlxra+myuib6BpDxxnVnHO3ZgjOX5KaKsDhqTCGVyiqOtGkVZqUMC4i/t3E6ipbE1Fc
Q127lYnix7Rj6TIK1xBViaJMocNEEWCJd8uiC4FKYDz8akbX0I1/qQxKMlXr7UdPNqn1Eog/GHfs
DR6CTkwtLcN/tEaISMrL+qIhKQyJpJlScKOctp9/beWsatfB1NlFOzfTmhMI9WAShZoyzDHfnQXE
5dpkTdO8YoccNX/apxU0Ri8CCyRZx4wyOVocJUyVbqyPK5Ki1wddfHDkplh+gViO/5b8hpMPrwNw
cIGlfY9bU1f1LiIdoto9VFrmFW57apMiOJLAS59e7cnL8zF0yhfYbCJqdawVVQ19dCrun0Yr6hB8
AQ0B0toI0M1AyFp3DXtLPbs4Q6H4bcT6AtdkqRByArq9QEpMdvCogMA2mWiGOyDXlxyAOEOe1Vl2
LXqfJ8Q075IJFlcRKndE91dap9AZbW1CUqTvoKAvAEgLIr9xmttUwMlDCzjuOnnZPP60XlUNPl7p
yqxoURF+oG5XSoeLiNL5ExgYnE7v3eKc4raquex1424vnl3fIjKI2EBpegc1cOdTDn27ENDpdWR/
8S0D148pdEsYLEyHq9X7YZHt1llVl72Ywj0axvr+7lEk3qP2+6ezvHM41xhblb7ou6PqagWiSzhg
ri4n33fAaQ/8qYtCdT5VUYmmbo6CxAXMkmThtoe+DS8O8+2vFAplvAB7X26eomKmFjwg3/p2HY6K
WpZZGwxhYpXGlAXla7XtRX3Y2VB6/VrYspsbK13xz77KFIQwAAXeYAUOARiDq+U4GV1i4yq/V5bz
4ZtHI2ufQ8eJqPXHFk3KZc4tgD03WzSr541kM3VORb3wi64lUviM5Njc1PmFQKVU5CeoFOzxc2J/
TKwUx0MXV4tPGguQcWioHH6ciAZ9pg070Z+84ZIqe2Wa1Av2OJSUnNoGRsHCSG07pkWe54ZtNeQR
ocL16BajhPtKH+WICTL2vPfQoTGmugbFIHlnblJkdZ0cmNgh+HW14se775eYmB9iAwMYlso5LbnK
BUD9lKZRqnu5dBt7zcmkej6LHM142iZXwxn+QZAFh23DeNVpqLD9IiebNi3JbqlYyZyT6BQHnBUF
CiVcoiPF1hoQAj8YtZL4FLT0SLNIoaoAA6i9lzpnhIDYQ65kV1qY0ZgevIjw2CPB57xeCU+RMs7j
9KyADxdBTvqtjbRfC51jbMMRTisOjl+gqNGfEiRGOMb6GLn4m9boikAEG2/iZownsVfCFc48KMXh
PbLYwFMXGPq20b+iMhdEDmaLOYQeThMXC+xaEHjS7OmdQQssXxEAXVe299JKaSKAa+UwTb0P7LsW
Jl880LtZBEwR+zy8urgKLgZOdYLqrKxHRLG5fffqWL4wOnuvnK3B9+nMcklrzpFrtLxTjCD3jh6R
AK2OyAMWex/ozZURZQoUFte09vtwtY85XPF+PLUfsPsGRW5xYoU+SwJbADsI2LQm/syyrn5/m6yV
fMGe/r7Xuef2tqyXzRzrf+Gync1QAtnZ8BJlJjy8BNFDQeTEmsZ49VlBDHigiNuevM31mN2qZj79
K2AvsCGl9sgpS4iofxya+PiP2LXHxyTIHn9UZ1pQeD6PlPqrFDAtHDaaYb9g2GC8NqTDmMTXJ1+V
5Pyi1UgT3fzN8Yv4z/ZW9cahY4vBk22kxcq9NPBwjoYS283P8DUcACPHfJI37v1JQ+8PyP/wx+n3
qct9Kc21wfpnfEVMAweWXWoKSZe5yyDqTacZ978zEeYfVk+rKnXSF1NFEqec1ymFfdysIAMNNFjB
hBYSteOdN90tmrlF9bXq88hOIn8RXi6IyKK+5iqvVc0vgIUodHt1R2C+IxiiU9ntYX9Vs8NneRj1
8LjsNJ2CkX+5N1XJFEzMKwfkfI+6lLEWvftWtw8/LfsfDtXtVPq5+genA1ZQjK+ys6mjYXPIMICl
8dnnWyDvDTSkrONtFJJ7gclfS4lp/27oIkUNZ0V+hszkwPVUTQsf57TTqMzU+03pOMhtCii73oFx
LyhK+oHFGYsbysuEPIiwEHIYvlyGTnkpT+yeflAo7eX9pAPlWgl7DpT9gHZCpBFp3owm6ONQaoRu
2y+ixPqUU/twMR8GuiQD8FFwyvUI3iE3oAp5tIldZDPTAVRoPtXK8ER3z2lw+YxTPv5BeBBhUCrg
X0mZTepcbXeCZ/YmyX2c3SwnowMhKwY8caBWVSW5ge3mdHmw8CEkgYxIeCborlb7E4FAkxwgfn2G
sL6pN8lk60R46gCuzXjN40Nl7jKPLP26YklPcNMWJXcUctxXih8zBY5h4uFgovZXDiN3r2TcETfS
daG5RQ1WjhpHZ5YC+F+9IDLMi7CB8BB5N6nB9DgNa/EUXBR3/rd2tPVD0pT/e/th6q+CtVNKhRok
RBrWJMCgL3uId1pM1DHJdemkDqx9rUE48PXFQX3WZZswrENo5SwbQ64V0UitiYCKETd4TwurE54t
G6yywuymOYoQSPA/qnEwNr0Eu2dp/+k/sjV2TwxuRP37TjYgRyrnq/XSprPWJPHZGhsUGsTC6F7u
aDTUnggbxz3Iqv9s5/dOnmISPpFMl5739SZMYYYzp+JXbznwmWPINbEP/GrKq+IFrO1GQyf9j5c1
cfAUwaUkmwPMd/Rb02B7whQjS2qGpyyTn/zrVQaARLBT9vWBEQnBSIwyEf4zX9C36bai31Z4epAV
HztFDO8HWgIupsrSyWJaRsPr3fKOwcPgAUs5zOkdQQ8U66z7wIXFh8ZnP6+nVW5VIYjbnMPvHDJa
gFOJgVGD1jre/WF8DH53m4rPPDyCxhazDXjRUWsL/IdI5ae7dF9eUvVG7vn0Tn7mt78/fIKr/xJy
XC35HCfWDr+RZCwf3/r4K1LCM9U9Fknq4tGqM7MSlLNfFvRZu6B7D8O/lXEl5BNKGrvpxImb+oxn
mPGH7QNwiKKn+KfTwsuoxoVELBz33jX1GFjOmWrForJq6FeVB73c7N+6oQoTOXsaRNEFaFWPUBab
JEAa9Gd2x/EdrIpT/t3q33t2cEpwl8XjGVB2xkSx43QoS7nqiikPdiTuSGKX+V3JUmvh1ahgX9uT
fvNgjhAWqKhu/fdWq0FH768pN2U41X06ebTinmmjQYhWNwrFZOd604HyJYnDYZc+LQZd2tyFCq9i
Fsj9CQIPWnzWApwnez8+tl95d5mN/5JTBO8V8TkSVcpq4YSN24CZsxqgYSvbP/kBMlshK3qQBE3A
lpmMrGshQ/WukCDE8AEBcEurMaUvJ71jddr6z3TQDS6CgXgfV5rMtnrWtjHM4FFHEj5JREMNtsyw
ccNR8n6p6DboonNcuzBc1wFgjSW8lXrA6H796mdJAZDpqIO/U5zV0TbC44RryrrCFOGBN7fELZHY
AAYBzqf7iIFbIwn6Ah6mOZeFv/iZN8OXuvgI0BLttveEHq89zt02/sSFZcx2tVN4S49R8NFQXxi1
lESG1i80yK7zNRd0m+KRUiV5YDyCsHw6Qfh9/vV/DVUAI749ViE0kjKPYQgwUWsghLGkNc29kUyM
0vRN54mNowyDW4QEmmvN+sbr6/Cpp7o1GmQzlX18otu3TCl0kiJ1BKb/rr0SKDCJWYGOj1mfka7a
PlZ5p2xEfT9467wtdycJOUt4EGy2uu8K//9K4iVz2bbNsCSVJun0zrGWZk7SYGoJxohmC//O2uFK
ETsL5pLKLFgog0f/WdxvcI57DUjxzsMQRi8ee0ARlX4Zeg9e7ouNVNoG1qPPCwkA2fwa2xL4XmOC
+aRbYjuNmHBwS4daSTRBuzPKRRUUiWVnXWCUUnNrtb2g8uMGl++Ojd8Us3KDDFo54dtp24szhtfY
m14YVGJvGlOe4lTPUkSovv1uCGq0FaXD5im4hTEyTxM8BxMZJPnkoUKnWG5O8kXs9xk02v4O4Ee+
Z+CL5SurBh+VVueWi9fERrgpS/yJjfnh3g4DxKbCQCXkLe+HVlleGUErWTZma7Dq3PShOA79pWA6
uvXBi5H/1ADo5MINcYyRhcjZt2rT0PU/vcd7TZxlwlypi03N2zEjkN4GQEVQ8e69Pe7qxkwY6YWT
om0xeo/0q1cBJCwMR0SiLudOkGVFP6CCpKaATM7XRWih/+D3Ew2dvxhCm6v36zYU0Py5nlA4WlzA
UQVB48G+jsCvNW95NwqH1gcu77QyWzg8n/gROGuykrHGB5VfVGaHtG549VbufoIzSJ784KfdBSaC
659gDoAZ6ejiWla1rgOGBbz4JfFRRnOougM0jfMK5Cm062u1j23COotVTO8T41CleHPJse38rjoE
AhK6VBZt6W68TCHZLqfzFZ18x9vN8fuq8NSM+Wwcq/wMI5qac4qoGpeyn9jwRUXItMlWHK8/Tq96
wYi5lOWqHpyUs6JNWJVPSOxW9SvVPkZPFwqxYHGzgwVLXiUk81VYy++/gvth+PozvTP5BxJmajJk
PyzHLpONj+19wwfBpf98oESAVCZ/NIDmWkU5GT547/KmKArvXT90mWaFdwJw46bbKe3JnNPav5ft
68UTnIW/JWYXMkwmw62xYsEIHWMc66bRlrf8k54jCAgwnoaKaTm+RriXUCdHeEQT8nBVaXhJ0YAy
OEk0SjXhmdPR0wzGullWHVD8U+XMIN9zOz/0Zff6LIyEZ3Ax8ZWrGsuYUjBBUE9/9aCtkjXmyzpB
0e7yxkTzyeaXoFxOf/5OMqre5EjoDZ/bWIiv5X36Z6LMH8xdf2bUez9Reoj0gda5SAvrrhbnZNih
rfHv8x2qpXqUztVHtoiQBjqVbDD74Bvsbbar5+/Ty1tgbmSAunUp1VpLOxop+TiiPgpKGH5HVAGB
3pEr7dJO1XbcDSu8zyRCcSZGKmDne4aW5fKuoHbRtTXY+pHNWley4sQdzOv5mCIksRMUym5oSHzq
xNCXTo8Nn19uC7NLRik3VCVnpGJMIj7RRMWFmrNOPXUQY9CUkoFvVDfkxfHRlcEfFa63jTwNLRX1
9d5YWHdSKIICj5zhV548e2cZMaT5/KcXUu/LZ2HdDkqZAjJhOpxl68Zuox5wnDfxV53Kv8y2006H
GyrJ1QxYb2tm6qovM26crd58nAUQkBSMw4MZrqLMxMYSUGM014Cq58DbC+U1qBzU0jLlSkwJRKwY
TPT9pCwifS4ti1KzEdCR+1a7Zgymnz3S7dkiihlXp1AmZIPhDzIWJWh+0oEUnSPIdscXAbhdYbaB
D/qxDizADx7XvszkaVHWkZoXDrto6Nl9LvC0HO19Vhg4EPaAUt+Y9UqZL/P8wt3TWAsHleFftZwL
Grop7Re+ixBi5wRVxTGg/ba3cQ6dHFEedMeLis3L8zl5fJCqoxc5M6+s8kquPBFx7lCh0fF3jv7v
9JEAI8s9xXGrJqz5NfSThpmxP5AqOlN0ts/d1dDM7pJfCuc2YD8moX4hNKb4SdAnBiz73r2+HRBf
qECycZQ0EPAMRSL2KPXuB7sYA8mM+jqDUwMRPIO1RWtUGeH3XLp37UrFNhN3txbTVgCPZraj9lVr
8ZjZ6tyG9YZbpgivH2hcXdZpmjO5wM8L4u1pTmtJbAf0Cf3bqB3NxYVqf+T1Nmt1Yyb+HlqYX02k
VsUU56yif9CkyzXlg79PFN7AB8pboIgHAFyvUWnmY6ODWfj6O4M3QH9jwDA+2RahpQIhxkQ4W042
YhFVdlYYXHqSM5H67tSIkBeBvcuxHMokTa2SR8TRMYJ3fimk8XWDNLXuuVVUb2BmXzNRCEKAXViI
Bfw9al8vr19QHfDVKwaYfJri23wTHMyC4lsIVf+hbmbIRtA867o8jjWr4GXSKBaxR4+y4ATDkWLd
XKUvc70nlbrKTGB+7CXHrzxRDQ1bijUF6OXoN8AvRutUdR0jQN/Nrk+CbJb0iS5ZnMnECTx1XQ2P
BO7df0ldzLA/rMit1wCiFSaGfrpAtaCmVeDpkqjw0nY3ZasSLgA3BIYx8G85tN8DPzq0f1yITMye
Y6GriYUmgNhbj+hk67DBlXVskurGWgre6esqMJU29zHW9MoPXpsFRueHQ0YpWfiTduapSYJaYj+e
I6LaJQtvoMo6ds9L+K2NryzgiRlpAUZ7W5v0kVjcsC8eoGe1o25uJVLJlkhUEpPnH40JyTupX2Ag
3KlDs19iQAJ9OQOsxYnXRT19i1y5mu+U0jJdKWrPVJrbQiZ6flBtu+JlSlrIg+x3jTrXubTWsxkt
BEHm3KFA2LNg4bmCiuDC6sutPC2mW0SnMesnm7tbpGLTBVgEE/55CmJDqYSpVFbJ0FHt3sOsmt+S
qHbDn9+0rndncNDWNqRF3IJ2OPAFGPFuuJxSLSC0FYQgqYqgyJSUZyoAGPh6DVvFsGF0d/K/G3OZ
fcUHoBp/WmR1M9wLshMDbdqwJW9O5n+NMS7PbCsVTg1+dSEEZSiikJ6jcE29JW2C8EctfF4tWBae
4/4iJsdqWVfUauiWA2IvXw5ataWxIn7nSH3SjicN62Jk3QgZ2hfhQVC8u3lTLjHHPROAxz8iVvUi
ItgDPioC3xA05RUd1to07IAFCuKJVRfNRhW2u7gJ+OfADpwP1WG2N5i+O64JJFOfthRTMnj8gOf9
2hJR6KAFjMC7slWrdiQ/JQ10qty95kj8wVIGGRe/mcv88fR1lkrUObg1Q2w8j9+9BNs+ZvWjVtMQ
TlJHqJ3Y8XPNS6GB1TRXDqvaaLBmWDypUOl/+g2i91vZHvh4hrukDkYlhgWOvU9hUQ8LJ+6BjnRV
40AXXPEWTCH1G9WHCwImDA9YY4paQqQtZElKSBjOgS+1yPI2eoWafc2ZT5lQ2dV6HUhueATlTvCK
wqMQVMzX7QnDwu6bmcyRSCKKrdwLOoKBlqzGNZYEaJZkJm42ohdbhltvbK2WCJWl72tra29CcsOG
WDwjgXeWUwc+GmyELB0tu5R5ZMTze9+cfzYEnEDn/ABsj7PDx/kfjpUfjuXA+k2uugiTx8ylb/k7
9QQTEPW0LHnsco1PsL2s4EFeM0yO8I7cAz6vhXkt1jVpE3bxY254lBhSexUmYcjXwOAONBgy8pml
c7amXAewyPeaFPDwGisyb6s/HzDeruaH6upOY1EJX1TraZqhlvNp9ns3QAm4CcCSloBiARxlhEDa
4aXiUZhAgv8zjSbqEZf9ln8Dph6tGyVg+Grv3abmVZQuw2oAWC2RZNCfjPOdzrTYCop0JFazIsKH
hyXLE1r5SHHwE9G+g/jII1z+iVR52P8UuIBNf2p/955tgdVU5uiFTFfJaADHnPMQBvwbqyAggL7D
OGCUIq8DnLV7fV70DqgC6roiJ6+IpoJRfR8thtPrzsb/jGBmiVb79p84kwtJRrQeYXCFHHxxCvDG
z5LQCe6TQFR46pemYxGO8GJL4HJ3fKuf5xM5XgdjBKtcnoMLo30uN13FaWot/yLYKEBqEujCaHZc
8T07sasarenWRvIqc9eJmq8lW8E8W6sB7uv2T2UhPC//HdM0iag3Wmg4YXkl4P5emuMr7UF5HTPG
DCkrs5VzfozBupGJsxAPbNLK3RVn2mpripsOMGHTVGWL0sKJKUZtVPdYDzoKn3RRwLzCiFTUBmHe
T6ZNKrVNgmg4OohtFXyufgc/DTnrIrHje/mQKGmCF6Wxu7biJnE8ezrGIPPhTFAY3Egu9YgSopnw
YZthKKhHmXBrHDsca3LYIEmtQNid/V1jjmUrs8xL/rzeTv85K2OCqRmSqrmevxc1DLQfpJ0XYIfG
TzRE5ha0PQSWEqXVa0VeZqPhz1Y5OafbdTAqiBHy4kogFSX4SLZBWDXFnBpzzFcwwDAdEgkld+MZ
ualWDuFas8KswvzjBmm6tfAewFlsID1zUArakFgQ1Y2Hdrp8+QABJ5XrFQB+1BpKxJvYGXE90ZQo
2ED6bLGJF7Tgg0FuH0H6A3wcfmQsr5S8B62UW6DBYM5zmNGbGQNbm6dM6o1ey4RBxrcXrWzVEGGP
aM8JmSzdXI5i+Z1t2MIXaMUg6feIpryKjhJ5+WfzPAdIr/Xb1EyFNIbnmBjr3kgXvBTIR6lH2oyG
byme5AxAWHeXRweQmYZRz89sNu6r0SagQ8gRImE0gWda/J71YXzeWRnUg+5pQKn7xCKhRL4QygMx
BTgEfxhVYhLlK775wzvTIoh46N/tOv0wuqW3jiwbqkvwVGwpsZwCHxhhjM9pYj6U+Oq+nEnYAqYu
q3RrBTHBEdXStfUTxF0Kdd6Pui+4UTXr9xWDQVlv1qXA50d31x4sijLJQ9Au6GHCXr/v6ONfBJYM
qZRs8YP/I2sT7eNzRIkKWcF2QncDgVznwzIH6bjyk5ySzUPrnbNqOX1lbg3NXEPCImnBHqI8iNBV
+HNIfxf/f1kJEbIVdkt6tX12syqWfUY6l99sowLnQEZ4f3/X87OUWZAh3aNz9RgxIunWHux9vGBx
y9PQHXK/9bC28vA2cO/uYT8E2V2RYXg3dRAY3D/GWTGuTpq2/Lvu8irzG7FLQNTPQgY6cKGMognN
fLqvRMLZ3Jyk3WbA+7g67YW6ohye5du79bn0pEWeSRFYVcdMcDPmJqEijKS5Vm60dWT93ANKvZ5c
jI/fJCp8wvFtonojmEeJ45/VW8/d+qlyrvS+nVM9KnhMTasQhu+H/G17RJVLPfpmC6Hzxg7U5MKY
z2fpKOxj3t0qfEKLbvzWSe855CkUHd8T3ubaxxumo3BXzW5bu9R4iwopE1uP27AcOOwoAKUUJKlx
jRVPOUodV2bWs06YTW04sPV9BMrlvDwErFHinBU7o0u2sx/nGX8vFqFBOLzuccN3NuFTUhEa8MQn
M23h4jQ1ZjLB21kO+JJmZW55vH43hmtIOgSrkZ5NdS8zW0BUlDu41rWT3AHN7TWhObeiKNfZ1kzP
HWdP3Xj431+CCsw9jg31FlRRtpqzOQsG827Lhi7Lp4M4xs/OHsk9w52peYsspdcwL41oJMJuVyWP
3cjirWTFuQhOkc80o6tGmTXztj6M89LgAA6Sc2KWyKMJ5JFaeh/hMNaoRYu3+HAnLj4OUowAyTP7
6/GZMLPt3mfV4pxZ25K2RZLdPHBr2VNPdTgAWm3LkryBG/s/vYjHD1ZUQ9qOiMbzFHGTa7GKzEC7
n4UJegKPi/K6Y2fY4IWsFTii39OxEJt8hPGaIX912mEDAE1XQvt60lOBIEXJNut+P1/CUWxrTuTM
+8w7xe2f31BCpdWCqNikVqpNsxOj8dIEK7eOrusNd/x5A6J7WysNZVGzAmLhWOTGAQ5/CFlqVHxt
91fo74jELMKIowFoqym73zgmA2MOrjgVxekJuIEV8h0WKzhzEBMwyaiHelcAbvi3EZWFSR0zDsnG
n/rd7RfKS2fZ2+GDzvmW0xaEWJD1hRNmZ+thw/zHMnyFq7Ba/qkuEjFgvW8Msj1fOBmXjqAEqYaA
+OIHZvULOnuOVJwEyWXmJhr6DzxU+X9XkVr0D4kNpMU1eEMJ/FEPxL/0IQ/8WR2qixTEHfOPJLSh
V22uOWb+TzB+m5lFASlHRC66YjtzDS/7QfvKB9yCFwoioHVxN4LiUjRBdBjbFWSne7GPflIRfxG6
+lS8x2xtP7aPzsnk1Ysz5CKMoofc8tlV6o9tGsmKf4UNvmaWo6YdsLkAJpd88wlfZrUK+D6Qno/d
oAljWxddY5v/gNyQJI1Uu8Qh6LJEFS3oEkrItNtLXcSiCbXQ6EJpcgrJ34rSpUsbyet7K/+mL73w
iKrWTbeJqToKS5Bda9dE47R15yXGQH627/TGNAzQxNm1L2oKPN1qIZ5oJwEivLiUg+7YbP7e1RtK
XkbLlMdlMmudrtlfIiQWaG3/XLTBPakcZneOSQl8bQ0wMC/5426zEgPVKvI4eLIeALdzIcigsqra
UtROd+Zu2ntf7GCNPZK3RO3F12RV5Qc1ehZ3Q8ab2ABGH4Uz+YA7NXnXBuwsIsiM6GrbWd/JNZyT
VvDljwXViKlSTeGLfoOz5cE4zHmP1jZmN3B8zJQn3AzQJA2mslmiBRNvQnbi9oMS4AyqFYPpf0vb
11UnRsiKSA2OVlvKB+hIkd21H9hi1PLB2Cu+PFnwX5nMKpqT/t34f7GRVujFBmKyqIBcJlOdoDvY
K1f8G0zC1KHqN+dX1bCJeEPpOaE/5FQL14neFgRQWXQUeFcTqAUWkWxQIuc5OEWss7816mC73jTP
3wZBg+u+FB9CAag7dXpGEbEQ/I6BYu7LwoF4HF0yfU58lmTeBaI4lGVt4uKYfLvmm7uOx2Gxw2Gc
dSw8A0yVIRKmZ8AVxHo2c4NksRxmowE+iw1BcDH88wYfEQSgYNyfS6zJfRmOThyb6rItwkFbVz5P
pJjbCev+HWZGtn8VGqxxBpW5pY0iN8V7qlP3gN/D6KckBSmRWvPVxXm0SgYJD3wXUQPlTQKijztE
78Cn8zLPcuhWI5zTYignbf2AatezlSiSOQQ7rQVzitsQIi48NVQ0YNMqgXpnzlp5DQo2+ZQaFBXa
jQ1Ojc2iF0ttZtY/8txzd1lKqgQ05qmJNRa0H1W0xlBkzAP6x4IP1TFNAJeRyN+XXAizp6thHPIq
zXGpLjxooRZWPGGADgnfBhp8rYQXiUO+w07oOeSnylEVqporP0iSUB3ZXd8uDT3WTh//MWQmadqW
1WnjE3KTEBbHtQ304ROHHtXFaAoHrAgQanmL2ib1C7uKLzmxr6WdIndtO22Xuw2Spwwbl4FfkuUp
rmPAPDciMDZeJzYeoHR95nf56PQ1gIiBjJ4AbeIUaUyp88LGa3bUN8g7BisOUm0XHOZykyL9v+IG
0cy7N82qvaOiMeTqt6+xrhuTvD+sSyyN/4OPxt2yPO6XV8Kx7yGFmbNDwTv5qSnQXqNOhDLe1Xh/
2CiVzJYqynZ4DPJK3vy1JTspkY4o7xhlbSfMg7mgs+Wy7QcJKScBm6qNYDvgyzZ0Q2Had38+rxWc
pp8iVGMUEvJ3RipdUbYsbo4U0e/8YnB6/O7q8OLIlmY1niqygCF63i6mW6DQH+8++W4Z1TX1rPcm
v9hJlmHpHX3BtXd68JVNHdkgR+FIx/NhbDytk4IxiG/pSwzHqSnMf4jCe8REqm3lXoZB8emd/+am
So/AbfrVntuBB3rEhHEibbMZLE1Rm+ccpilTBC0d2MNwA/P9IYHwlignbBZosj+Vh60Ne1Uj4iRh
LW1xNDWcKn5EkAEPrwV1yLC3/oDcrFrteXK+7hgv3Xh2shRCSIRl2KgsAVaUH1ZrWHUkS2/vqJjc
sVTOx0F0XREg06irYbPMVep+tRCIbIH+RbU3juX7QBT8DlNRyQtmKPKj8iZkz0k1HeHO/jBLR/2N
bbFLu6Vd/LpiJyp1aQj9ekMjheI6MNOMilQwYIDjgb6J9hJurWTrHkzBHDCzEdp+/eN/3NPnDFD0
yCK4gvFprZPZ9YVKnc6KV3ommuVUvezyUoPaQxetZK+0B3hW6w/V2KJ/ofKsWcdAH8HVw+LZQK9k
nVRoTwAoK0/vAkRzvMFUQ6667K8bk0/hX2iEWhz3NnuGCo5cE9MuGLZ2G1CrdK+QfvixbRzUJeck
C7sCzQydTdVr7Mgion0FGxhOwfWMmvTUXOO56Lm0H1DbF668Xsn/10/ewoSOywQkPJCKR38KDAmg
t9cgkg0hlP8V+r3jkubwSRnpDfngrctc6L0x3BLukWw97nCMiU0WtzN0oJ2111o70B2DmysRUCAo
kqc54301zL6boV5O5aMf10aMNL5n5bSVCmHxU9fIiD+lrkfGX61NnqP1Zi450xcc4zedFMuaqoqv
Udz5HtqmeySHB/7x0RU7sgNLFIj1vdVRL2sVEjULeYJyoxapOiCIbdmd1OZjG8y2hmikP77bwzwl
qj7UevDmrusjYBQ4xJofUJA3AE3BoJR7i6PiZIYbRmxdowvGqKIZ43SHaIqSLGrS2CLJx+E3MDo3
Ebqhi6b7A5C0bK/4CC/YyGLjpV1/oGjod+4AfLrnPyFRLQq72m6D+eSLWCWl1SR8Ii2gbfSf4DGC
d6MF6R5YmZhu/DMY1tR7ShsGineO8h1MV0YTlMhyUIXsStQZbNjl6glYo6W/1JWbOGHWwWt8s2mb
n4sdSj3Y0McbvSGGAT0ifTuOM5VAk05TRLWwqRMndmr3JJV4MIM+BDQQvNoXVGEFRmqI8e7pzdGq
a5ZBFYcwlK0INGIfTgCIOrOH4tEWCt1jZ0PN6U1sGXQceGZInhesDWwbw2elqPLZxo+jWRYD7gKt
4FRrHGum/f3jwohjIermnq1f7WOMg5nNKokpepWsbwnpg+lwuXsurk5gJEyv8hlb7exeu/McHnQE
xrmesPtyOdklypKUqi8kEPXcOI/dSapjn0tZ4YaVfYfpDAdw2nG6RMnWznwFtQscAruNDi8UEDUy
8iOv/wY6d9WyafPpGlq2ym4EEYZIj1N0PJC/WPwnp/ZmkNA7eUiSfu52CB8MgRNVKncMgxLOL1gY
+RtuVXhEFJnUOBf0GCHE1bwQ38g8TgImTQQO2npa/duMtYqjrwAimmprbiOR5NPXPGKeb1YhJRkR
4keVpxJjXsuA/O8znYtV4HJmRO47lffELGPbzM1xAuJPuyzHBIVVnlPN9daP7ZUiD1KBHWRlfyzK
3z7UXVih4VWDALbYvqV8bgGH/ZvP6HObZYOnJgC+NjDhTN5GcvG79R6SlQZnQm/6kqjTSx9f7+5c
/TFUumDOTqRZvHvo7FvG76D91v0auJCOG6EqZRi4W6xgE7gYHjkafvc9Pl7NmJfQR6/zKkTzDJ37
9/LzRqdunYVwThNwrszs383GZq41YpXJu3TZ+nn96XESWxZNHZ5bRBaf3iw+30Z4u1pDNRVlUg0c
t3qlax+0/xPGeE18fzJ4T3JA3Mttf61GT3X3Aa1jO9ipkqun/fJ2B7blTc4YvvmtUZGRqvXtiUGg
e48YqoHpF+pu6Am/q6AT+dQlt5aQAgGcaKxDq49pD3uFuoxLKJLVuZnFq2Q8hTITjU5VU+/VD1VF
CguR0cWiuYcStwWjLOtFHvzbACnXcIsWk+2ZlJVc6TwClULZ9mJEUty+tFKW2Z3cgrD2YE8U2yUn
Lre+b6aJm52XiOFYgPT5+/wI3kQncHCVJ4R3JijXPECXjL+haNYun0F4jXDRP3Jlh+eINSu5rFsy
o1Jvl5No+zE59v+0l8aj6ux9s+YsezgGKgddHDMM3kSukqUDmeQ26Hiq0VM3Rms3eVzsdMqUtdDT
xGJOyr7FNWN5fxalff4gMt9rOQsdHJaPMz3KifN12VerWUeaReDi/vtZ9xAVEQvSZuliKwSsLc87
ZM4fDhBd2E3gkKLgTNIlG6hQI0nvCDBVymJF6mxQRNSR2vfFNs+SrEh4DeJeCbaxe+/j6n5ocQTe
dT7AVsbs0adgBOaetlOXNwMldDFOrdfAVg00qyfkdbV1hlct3pnf9TfvUvC37Z4yvuwtZRX9Z5rh
F+oaRT9sDELEefekxFPh75HGLdEbQqDUbfljBOwz953Dbvn3gPKDqlO+u/1Zs6R2kpNxVZybuY3/
GQx/5h1FqFbFDoUPvprg+3535YP5hfFKBHQTTsWZnfJS1WsvCW/nrcIf4GHS5XcYv/+vXNMSoEnk
yKm8pi8hO+NbvaI6zgKBK4ArCcNPMb5QFWaIkdB3ibLEcdWui9yPnrx7yIqXxor/R5e3pGQtpzB5
Fx4Hu11125N8niNxD5Qk7mgtXUU+HaVSFsI62HQbG+OtSdoOhPyB8wvebX4BNyg7ojI5JuZMtOrI
e5D9E2NmQ7+QJL2huwbGkSU71fFI4WzCTN2XK5mXl3t1yFK55JqQle/RKvRkM/9q8hcyI4QVSJvm
GFfjpyINjwsaZRgSg5hQvU6yag1R/d19UVuUvJCMZ6H2kLEFdGvO9yUj+7L7JVXxNBq4L2Yj81YP
E/5T/BPmJXu/7zZP9i2w1iSUwmjv67i6daa79CqMNjokLmNJgjwA9uWl1/l35BrN9SlJboTARCkl
n7bVCwyVE3960fYqQQbnj2Sp/sShCU/j56EdHpYwjhoifgddBc8pHv98+Pidu8TLLpAR/2509tYS
eh9cikK/P/hLK6fshftS3QpvFT2TWNiWINhQUdlpa23EhHd3X+G1jtQs2OBW+EUxBrVEeHCDmvKr
X1xZntGTO4ukxxuE8LGWaE6u3txVFOIFRVDmIyXn+gfxqEijH4vkKRzTHYT5AfBlzIVQy2jdfcOD
oILexu9M793Ne/XJ0xZ1dQ0g5H/FCRWtldSBylQRVI4bNAEAxH9Np+nWmHPktGuuJhqaYgRILm4Z
SS5BsnLl4/pb6GLD+fiP4dclOZGwZGm3uh6bXlWcYyYajAtel5hn8Pr1c5TjbJzszsvPJyB1KooV
dOaSC3Z8dlIx4TK3SF/nH28kzIuuFveFsO4sy75xQrc1JDu7mN7/1xXeQzRlC03zXiSehrSZwSSs
CxXDAf/jDTxmLaIs2Ha4gYd4RCR6M1AT1ZWNWcJidIragqvgaoYbcR3L3M0opdH7QRPqxIROPbAJ
BvGgD1e9sw82HfngZMkKFJLWkvCfyw6CnxRpwbX+3a9Oeq1g/LbTwDE0NXDPqpir1eEJlFmRdEhT
XXpjx5IPJyvOhNADman2Go3XD8+616Rti3Xlt5lbf0QC4fBAVBUc1uLUd3VwWwfS3XifJ3NpNAMS
CHn83u0j2B7/Rw6/XmKYaz2OM4wMpMpiiK5qJGfVRAHi3cAKLrX4PbJ48yVSOblgFnKNkPakF5IF
Bd/tlHAkUfj5r4wzFMbuSCSa1fAuUkPp1Odfo/fTQO8dL8AkfPmGeZ/eVI8Kced7nbNk0oE+FliL
YgFydiwynSICL4XuLd7F7qAHgwCMMWNGwZVtz2iyIbHUwUusQgSF2jM+AJgqlXlbQLGi6h6gthle
Q57uBpfWBIP+m2Wzng4BGgRyQtP8j72c0A2+w9k3W7HjKdcwqUqqyQutJgu2VSvx1PPTPxhdfJSk
xi4UqLhrZXLtLPpU6jLuDHqZ4sfxdSnpbOSsTBVDJlbqnrSjVDTHJxMQ1wCA0YcfHbG8jDbA5UCB
jjHmTELw8y4UU5vy+WoW3VI2+TnVv+UQ9AGK95P62TTs5X3jsYgxF+TsJfRqHjI/Zke/yRL+QOGu
0dCS2+kFY/Nv+jpfGR1TdmZQRpLATI3ba0htpSYdt614eMZGdQ6IPSoORUVZb9aUyfGawlIWVmy+
eTKRuHmy8rgITa2Qb4UORgXuZ+OWZdJgRRir7/65I6ii1IpGIe0jDMkyxe0HHOSxpW5SCJXvHAKU
fNLQRravC9qhwmLMI+UIxb0Mect0Qw8QHR3m9bfswLrWlw+0NGREUQdGZO653+UT/xAk0FHplzqq
iEitRiTXi8q1DTN+3cI16xLT097jFG9ZAmOcsWrKY6WDRgfvLF1S5Lq8lOSgBUtepnCQiER1pylk
L0prTII7Dd58TuAB713NySPsDQPlHt5sCXKWsoc4wPCU0nl3HUUNcMYL0Z/w5ToeewzOM9SJqq+e
5iA8wrQDxHJJEQjivPCYuWk+z9yCd8UKNGqgahB4ZZNhE6rgTbV47SOsjLFRj1NoREAG1S40b7Zq
5UVD8Ilv1Hnd1SR9QpgeZ6pjQkeMFPtYnbnYRCHZDa+u5Ig0/4SUiiN9hIpbGTIL8hWdMjprEspG
EJp/cTWPzgawJL5o5P8Pbk8jCkTK8zFVCZfe24Kfx71Nig3rEeWgFhDe5OufV8DC4AEpjZ+rpOiP
OrZICr+m29HjKK10hW4v6Rf0DQTj0LM54hEK5Gf8lIYhIOoua2DBY4vhbaQxYZthCgNU4UZTicOK
Ig1lfKDGzaM6Vp18HBQwNAixNhkTJTUoBdVevZHSCA7ofAMO4ijJFD5TMx0SlA0tS3p5cGJ1lXyZ
HBotT9P200FGAdsK2K4gG0K4oU8WKXDXiGv/O/qQU0RP/zmXX04XQ432y1H2Piav9+W0rQQo84lP
Xuog58qK2EWZ7KaIMNSgZ/tJP7sOadpzo5QVFzsxqLku4UovOiOZr4dW6ZWCwEWmTJ/xf0Hhfek5
ioBr4Zrpx4mvwqno3J5A3UtnkphjstVIXf/AHUtyEoRbvRMD8bDH76W98Q4iE7nOke3AYEzGCFIO
NgVmZXw/zTCgsGg3wNu1cmDzt5O4QYBUwsGHiAUWpKd/PEKwfiBBmDvWdeZbj0h6EbaPIFvey58C
aouKmTYhqtocU0721aLZzPU9+dCyjmFBl3HyWs76I/CIXsyC1EXKvG6SXOj9WPYZ3gmn9RbdhTdP
mTyLMujYcbInAhu6xls+yd40k8wmhB2R9Vuts4Q4B+cKC4uweVMP6T/mRaMhn3RU4gasXTe59ydS
ktK11S/ullv0h5JApDd/u+Xc5OqgpZ/Xvk85edxyK+qqCAI9klHWj6uGPWGx1PXytslCXN+p0Pve
Nup+dyZl2MId2QzWntlkxGzOPkABneWFgPca79V6OuENfRPR4WnlGhpAdtHecUoNolmTgndSfhB8
zzD4+CN086mf8BOafSv/r4RJDIRMjvgse3U1FiUipdivoxcAS0W/2FlocWh9fGqVTvo3MkoPHdZ3
4H43xbtDIKFH8w9n5clgnIZqLv9LW13vYpjXwyCGxhEGoDj2HP08MDh8ZSC4A5v9WDfHe4GMczRp
uY0CcG7BGyZWYe5jibZUkriphmhf7dgFVOhBKlZMQgZC11sBR/xf0eCWoSvWrrxidAB1P8ON6NJx
6voYmCrI5m74DKuNnTmaVvDzi41FCJSB1SrOO6/QlxabgsjcNI29Vpsbi5dt4Pzd4vUMJLsiIKit
6E1A5dwYhs5czXU4NR5fyl+WvdWWwF19iwMfoqfujzGcaWv5zaJWd0EIhS/MrOY3RfCZ59isWM6x
fEdg11MEY6DN0FicRdMOH1WYm7vGWeh96RSDbAT8We/WVuN1Cgpz0h7KASwgFH0c18jXbbObBNNU
eu4odeDvEz0bFGq9TBQDM3tIwS7lnyCW2c2Rfrv0iuIJFKXlj6pvdqOeopEUErnnnWk+8fZNpjCR
RV29pFYaO3ZGX4fnMu3YjOySV7Vient1uE527Gi/UK1FjBJsG30OyMr7VH0Bt8e2wJxP97N33H7u
strcHH/CZ6ap/+RkCqZsDuqSOc717gvabGhYhgSoltiYDYRieDB9GMtP5kDHGQ0035zJV6GJPXU0
tGGJCzzCrRwUhQXtnhQJVhZIMtEm+/Yip6bC6r9n6a1njGuv/iLvU4lrF19ilGmZIn242lQycivO
0CesUTIJfZbrt9xd4I8WvWJ2wFpuhtlEY0V5uuZiXoeqSI2lpD1Z26RY5+3VuaC0GRY2JYSPVhts
ekOPeG3MZyM4Vz49HMdVZ5GT0YRTvjnKsrobKoWsx6yEMuCie6GRCWSiUfEAZ+2syEUXKOSBVURK
MyhdeB0+LTJT/MUJymU9z34stw6stdsx3iRKcwowyZM+Maj8ssh/006Lx6h3PXLEbRVkGnxnaamC
gB2awm++sf8/AyY8EcRS6v4q9zBjl0unuv6LerRJ35nykjo7mPqyFnZYnDa+oyWuJsT86UDJEhh4
enZUiMLqVnrY9HsZdmeuZvkuEmvSOsPbncQE6Qxbj8xGnjx5gI0urD7sHbSO6wjrC+OYsrNwrwDl
EKVold+rKn01+zmHWegNjA53M45em1gxSY82MNMraPfVd++SxtZefzgSEY3wshN1RkcRdK9Z5Hfo
vmtqe2uNWX0Y4p+uGUDlDYGL+mc5iLASQlaIyi/JrzqhHMw5VO3b8rsGi6fjzcgoX6456OUF8mc9
b6OFEoRuqQF93EcvM0Mc6OxChXqpCEjnqbwuoOD/EJAf3uRMx6+P+S7L9a3VCLbqt35dJ88vlWjb
OQhZ49ltZKVw6x7gxLbLcMufzrRsNwgNKWNU7vwSwWarLm+6O6zLMJit0QKPDe/wAlTnCm8zuglK
fgf7LkK3oMarkhcJttnCjzZyyJGFfaXrV7stXTA1obz9V6E+rVmDbbyHklgJeyLFUro4eIvhlMEb
ANiqyP3jrBMG1HHQsjwnD0YWc1/0VX/fuBeMykjXpWea6oi6+Y5P8RSmqxtk247kyxqbGGh0Zt1n
+OowHAqJtIx9rjYn3U0aRxqFLX3/iSTuQPqaoY/z6NSsAmzLTP5qDLKqkQGnWXqY0APjI+RtKbrV
IzB0ghlw10KIwHBq3v21D5PYGUYkmcAM6j+VqVPjQF8vS2FSopvcbwcKNJWIXWZB5vGT2uvz018E
h03famlM6IC/Nlv+96r/L5tsr8vb4uuF+CT+XGGLKOIp4b3y3RelliQLOuE+yxGiacQ1SGKcaAJ/
qsEKg+2wNhrrY2Jhvxco3JYAIaDv3XVD3BctxzYHgFtSncO8FBgMHTRJ3Tz1w5fZFRQQ7h1uSaij
1ZFEUtyYhV4fHLKCYaVp1zTRUvt0+kJs/IEXg/hlrMlDlj9aB975xR5xTvVuqq+J/PI1ugjnHDGk
Fclj7L5q4nGIN/bHPnHwl4WqezdUZywD1cPpUOoZ7KaxNzk2QVaLW7sfQm//w6QfNE++9cFWen0C
b5tnFJD1W5DAcBC633xDAV/rVsalNoxb0RjtuVO6wZDdcZjKaTnlGy2IBomcmQKV6pzlmAiSxMlf
YhESwZVYnlBIXmcxdIJaKihV7qakA+SMnNNWJr+1MkX2cuZglJJ8lO6hRkPs6YGg2ikcbxjN+0yJ
dfbZrGrKvNBx4ArhLizTH36a+oY2eHg7YfWUttzx9Pn8S/9/60746PlXIJOd+q661FnsTVgO8fy5
M4qumxtJZ/HGHWAfERXhJEsIOZxdH2pdwt2Y5tBo6fFksXo3ShkSy91S30vsY7MyVc64IGWMGoVr
Lar9Vm/ONRPrxUvfLDXCO8TVpbFNSMBsOhSFJ9r+jcpT4DSe2OdN0lyrA2SbO55BqgsUVyP12XVE
1x5EGKPaQcyGtyPHQlsrx10NuQSvlC01nLc1swgvbLuz+N6ZZ9MjCA2CZ6ZmUak9BUJFXGpE4kyd
ShCGb5I4fguFrEooSX2HZ9cNxyGVlibKvm3bk0xkr93jjv2bWjheXdegIGxLWvAoKfULqBAMr72J
RoKmmka5O5P9VWHEkXsVzZ68h4Uw13qYMFRZRQtGVg/InBdMav9c4zUrfWUGm7wHMCxIr7e9A7gN
hJnlZhAehR+KdF0OODZXEJwFI3z7YeWdw11FvDgYC8HwbC65FtD2kbbDE6W0s3m63wiAleEa254O
gdmpQpdDqXUhMkFhQ65pBmh69AXmg5PugaahLuR0PlNHnsDD8vnuiEZjhUp++YZOq1HQLSZyakm3
mkueKiksJ7W5ryQxCT0GkIhH1KXCM/S+2uCSQ0DAvHWLjnstRhKPyNE0cPJe6gHuMjM9bZLlMwhW
XetR6coP1XZsHk1ozGULZP+9HgmrzF7j8DZvLz4kS2HJeOllAwvHaCxH8o2kxOXGNvBkiwkksePM
UZmfpPT9/tXJs0jZrSgCSxZpHeJYAVlBSNT3Dma9Lb/p1f4SsgmquPypR5Uw3mobSKjwY9LB2P9W
t3smd9G/ElghpuAd9EExzOxgimizz8vwFGX2dqHPfdPjZ0cCmW3x0NjtGivrEqq1duT7Q4WYDtze
oE6nvdtb6nEENCZSsvs042wWyRpxEa1xse5sdhgzRBiQ3y/wcl0JhMNUHQkSu+wABsrOYU8A+QAt
TG1nGGtRt6whuW5ZE7WUVGHTvHp1Knby3aPsKf1vzXbNd6x+EqIsAMIBExryDiuPpLkaiFU5fCdC
1bNl1+QvPGwV2Fae0QehBdAvyuUM8wrOsrzcp0MYQLoW6zJWGFMovtlCzbKPEUwIbJY/qUayq2hU
34tl6GQ5/6GBdK+7SVl8Kq/9Y8Kieb5lrIaR8pMJ2yml9TUKivdZnrmZLpMo/6w0mD8JDaojgtiw
Wyd8itBhGZX3QdIjskQvzACLHZ5PSVm+QVfEI9Q2OSFz2FNQdS5DJrfAFM1REIIOjLMQR46bafwJ
kTkrgluVhi37lvUWwFJLkrh+nWdDhZ1Sb3RTIbIWgYRKubn/3UZ9dcSMjZLPxwQlRvlkAWy/8PaV
MZ+MuMtWeCSDBhFhPcIaRNNSzOfTgDu/UrQ3wjorPiRv10Qge9hO8NRo5joZWdzd+FaosU41twXB
i4e4SlIGyf6dsf5N91XsFnMiu7FeGlCFgUxzejRzn6l2KKdTT+YiNUzNLJS3crJYS/B2KxuqxMqm
LhnSXKRXegIeOciDzODNJ3mrMpHnHrpX7mwLqBM4LtMy2QrjhHiwit/d3zNykE7kG2BwdrvUTEjk
p+qpXyJ7JrS9USPE9y7fCKNNDHXY833zZVemUvXV8VeEFsGwlYorFbYDb5O5IEM+d6LIL7tstbrn
bGVsZ7o1eFbZkfrKnW42g06KhJeJWCYfEPWbvFccRV5qaxIKpqdkB+W7NCII54nNvTYV+2moTVZm
WMxZhorCeR8kaQ5V29CZnpZhHbehKbE0Ez9VFLUSZqsTslErvXBIPPN0Y/mQZDDVn5FJTNZ/n5M5
1x6zziDAqFLp24qAH6SojG09o8PheWasHnvefyYhHw/RyRueBKx+OF8EzwlElt7RhuA50vxyboL1
/hvzdwMwDRY/ace2HEwQFOU2LPld58kBM+IoWYlcEL0QAhjzZEKY2f+vGB910RtNt1rc0YIXBAvh
2k7sE8zhbU5wZ8hBIA61skupEEaNA1AzogUicJQUwcLpUG987yHTluXBRbHlwXXOsYYISvsa3Bn8
AhT8bvyV2/YHgNXRJEPcGWEuiLOjZAYYzSlbt63cjAsmM/YORLcbYVvHWAuVJ+s8Vi6ZoRqD/jDM
sq9z5YmQZAHV5dXnir9VAyEXAJgc1dwvGkb9+U6SgpGWI+KCwNe9AUZXSXk5gfz/bv5nUCcdzDaB
QSN1awTs92V/NSB+WF10i05Fdd4SdQoVpc+xvkgGLAywgD5pRloBiIOtQMx7/7Zx+zHJNZqP3j9R
bnpJWX05C0P5HyTFsZrT0grgDqcCvthcEcmEcAYILLOdN83X9Cla3qAg1EcO4B0auu0h2Nhz4hk9
32kpuCqoUdXSWjhqKiSU1dLVBuMbxBX805gb/+HPYsuyXMsuHUSfFsWaxGFFMju3kqcBdRAhRjvq
F6QovWTgXuN0yCa0kenW3nGHCqA35PilFe018VP6Mm/fKeG6XmrAR9l3vNZbFNr/lTFOfjxFYTLX
hDHwihcFf4xvPOAfkThXieAtRoVJ7k8pGWCDWd1h0xPE5ozviyu31MM2Ddp/KGR4/3bzH5+jDO6B
V/Cn5EJyNjqiWPUuwWVXBjQLm7uie+4XPnPS5rVBgMFRQmR0ZrSuP9tZVyazQeTt8n1v2jMMfWdn
/+cjY7B7adYihI+xmMLB8RDVU7+olKAFlTJYFo4w5CvuPQWz6WNSvNLQSKcrEx3W13m8lZSSZxL0
He0S/0ffdtHHVjpF6JzBjS35dFeBG0V3KSMVicgojrRHhPe/8H4FjCBCGLY52IvjwD338xcFv+PL
/DFVe/J1oa4S9kvDolv/T/th+AB4TlyCjKTb/PTEp51E6Pc5V4efWro35S94ekIoVVAypE6Vj031
mNan645tnTq9DAmlIpbd87mqDj124sM10xaZHHsrHaPMiNJJHtvEk/G7qeOJyAKXLkWqgckOnbFR
1mUX8TO00of4neDQYuh9Rkqnj/tF3n0eyayaqXBh+6XMEpZsWFt4qv88B740PtL/KTLEcyqqhZ8G
HgHHaB3rkMjDYOXRPdKSWYpHWR1Q98ixFnNrVanoGDnAw1eFuDHb9wh9E7pjcPOBxCFQalou8Xgy
Gi20ESDkOneoDEfaZ/zDlC4txP8mflmOBKDSl8o9OveWFdX/Hx1RngLSLgJbYq11ZetWROuW7MyO
NsoK7VJzkvkqMH4suoJY4thLS56FinQIJu/zLyD2VMLy3EAqNUc0GHEbknPsbtal0R3H57NYuICC
98ufdoAF5zEO6vJQh6+ot+y7Edpyzpwu7ajqQovre2DwF+U6rnpJ5eIrQlQjMn99SNiXVLNlX031
ESA9T1ThdUO7MYAbHzPgItlkJQ8mYZ5jSz6VvojyKtfPs92+tAYMleTul/vyFexqjReAHxhKCUat
h2frm7ADGxpBkxdodH7Ldbsb1Sqo8/6ZI13VOtqJxZsluYq0mqi/1kJYLgxXW9payUELldN32Sc9
5Ts/l6dMFkW1iR2SImf4rxOs9hfsEai+NAeiXTggM0zp+4JyObaR/blaLjs1NEG1qLu6Imo4SIUq
5c50y0k+DlGKnUOH0Jn9PQHzYyQTdZK+n+K28a5tvkoHwNtvSP5bpxe2Xs5hvGnaUTACib+UK0qb
C2RxJ8tsVmAw6Y9urHTeCHrlpI3xcVBxN6b00rEsNMf5nfNIV4bWZjkL0lLEzsQQ2JSX8a4WjjnD
Pmxpi/rKeNJfH9RJ3fGFSKUsUDyOhcMIrzPT3EewNSW/cpSv99pRXPLxYbuaW2F4yhBfwh/mHWMw
Z/0dpe+FP1PVyKxB3itj6odgJE2/514V33yUM3q/9uPhJq4zBJfvmuTPVZABhvVB5klznD7hUPuG
x64g5eNB3jyePcZJIrqy54ErfDQkyG8mfcZGI2ANT9q/VS1gdN/10eU2WntneCX9kr9k0gosuBgS
Owo692bqBWRo8GFqCzlphEcv6fzSfRu/kRW1Q3DKy7zZpZGPhl6uw7W8f9MXG9cR7yx87Tqzcz5g
DBgvYUzNx2Wx2hkFMbrCaceem9MNqkpGdtouKkGvCv+OdovOAtwlaW+isfIjMIWnzXB3XGOVFvy8
iGLQCr4W8Qb6AJBcrkllyDFV9L2A8OMmsUwjY1nugB3XewWr5xgR3b9M6LI7S7Vkn4iR5hId+A7p
fGTrKDYhGNXlg58PZaRjOBTBBiMHU5v8mS/ysb6Mu+E6dlIMoKCXR09MRShmD+DNpwNQQ7vRgStR
hSrLOhK4geBtbkSEh1fJmFP9jkbn5txaLyzGEW77Qlqw9i9dIjGw3WWEL9jBHCCWH4zRxxTyOLPN
m0Efrey2dgwQH1q1IL4MjBgTGK6XFwGV/+VjFMIASS2B+m2tkodX2DLHzY7/2+GjamJr6Qv4OoAk
TPZ2VGM0fmhcaosgu4Gq6xIRZBtWSZZyM91onx4VjOqn2MNYST6y5lWdozG6QNVT2UMIYEduT5Am
JiDUm9CPgQhwpizyV9VznK1xsePLKfBVRQQZyOGl5i1RZx9d3C0tlVnVS9x3DK9HbdmiKMBnBkls
apve3A6uX8zRezv5P37sL00ITeAJVvLoq/BRge/2LgcjVzUBa20QardNLyGkJ5t2jBh9AG+fgbKG
zTLsJB+MfFBK5o4EQvUAGUEk6SszGydMXxdB1NhMtbIgHKkluFyjmnnCxavuOTmA8rbSD/RX2Mk6
AxzLcRqQd5D9DM/Nq6q73ptz6Xa+GrBfqdktz46ssnoEGzQe6+yyWZOMR7RaCoL5xyl9HJ/8OL4D
KrHP+nxtfzAtKtbee+3/4lYaOIYrTsxRW2C2KttcougnOpsgJIdzPIaCG1tDkvSrCHWewPq2EYDy
blSmtHGTbhhHExk8hxt9rgqGC83A1hthZQbKE066aBTpceV8U2CAIv/uK/E1JiH74e0hvhsTmgjE
NybUkL3+vRzdrqWGCPdfTPiCgu+um60sIxHG+W/zH4KATlvmJDudUNkIHcL/rv4wWmGVi2VKdNwg
wV4ZJYyNBFeaDe5HVmo/KWkB7RybP7T7ShZ8UCkhZxEF1wgx97nu4kz2u9pzCSuAIs+pv1EPsnjG
mgow89/anpJGhwPzi4lrxlgfo5r9NfP/MPgIrBA3yDfwaqjY/hDdKK1bc1CZsIRifLR9WXRG9XKv
rVPYn4gvVM8F7Kqinqx6Z/bF9m4jZcrgzSEuTJJAX2MWn5eh6anXKRsetbeJVFKrh+qOqkLNIVuR
I0ppOKypR2YGylR0tutfp/yUZOukze4J8sXOCCVPdt+RFAhlwMmRUj1cDDAVZsrXdxpNaLU+jhnY
JjoWNQm91UiLd8TWJSdFO5VBv8G2GtDx+HBp9TxN4/bMAl5qkgDvUhnuwUBErrk8tNE9TwH8wjLQ
MZZNSvAH2hgDSEK4Us7cpUW3ZvKxwzMAV1BjC5PolBAcykjMy77DKSukCElLy/TcGsiniL1FiUjB
+1kTHvNQWdt6lLrrZBH37P/YiDzkOmZVPErdzCT+FAImjl5jQWPloRAf/5VTeyu8IMsMgBie/pIN
xNS8a3bKZ3VRPMzL+XKiFiEytHi19IfvooS1G1bO/UUO1NM7BRxL0iZgVQ3e6C0scUTD4HYf9cPv
vPYoLrD4XIHX00woDvsd6JaBN1i3McME82Xv8fJ82ujPns5+9rRoSDJP7Jsyq/vuweA7OAmsrh/d
iEAXoaWBOB/WD8C7F9E0spIQwz5ogOKqjnb1oaOI0FsNX31ZRXRPB3bpnzX1wpvqijP1/EK12qMG
JP6sl3ezVvnAaLcCFNHLW8xgxiTD+aGq9Pfuft7gr6z7yAaonzskCAebgMg+X5Uc1UxljmEcOY3A
mR/UDZT3sDvT0sJVv79UZFiBqUIMw7oCeC12b/pcTtisoSxU2jJcEcGI08/Pyfe1hzltK4a/KFVd
q0YVNyNAbXTT/yDpVjNb3dfafF7b35B74zUPO08EZMjbDB+gGPOd2JdClwpBuYfDiFgC/2sKD/DX
oM9ZmyPsR8bVHn45n6B7UGHNrbbTfSGZB1vW13NE5ZK07gYCQRWLENqlJXVPgeZnxd3n+1wuRsx1
vERd3hv9w5tGdeNRu/xQp/L4IdvEowBtjqmT5o4/tiTuIsMqWLEcCzXMgFdVGV7gVOZUmgRGYWZP
XyO9KoBqAiewBN2LrfwGBhbdKrCA93goQ/vUULRr6K2Cz0TX3ctK9qKabQEmS4Vyan5QbnJ0pgXY
71pIEcKuj9/kYqVmbzh85eu7kynZKaNBgoYYN5BtJj/mkZV1BLiVYmnp88fXZXRcZSaRY9YeqLA1
VowY6DWM+rCK9RwSDQTcEcsyKSNzAYzhuxTRfqPmH9RNOPgMLRlepJHRiYy9qCUgBA7D6ckPLFlF
UGD4SRFecm+RRHQvCMAObVNg8x9zhEW6sinEjF0c549Wz5gAjys0ynxcw7JC1ZYA1ptC6A6W0GB9
+Bdk9kb+uSCRnTWNI/zkBgYJ3DEuSj5ppmRaqVTKOCZjOuZzTkjPthbt5y5cFw0HiZ2C0U93HaC3
LV2L0XaJDIAtHfu2M+hgq4uPWoarorARyyDqo4m5TgU23wVDbMRAv2n3EIbmSh54u5kkzwGgVp+O
dWONM6c6DNbmiRxMDfNL/FZOKmr4SjTYHjR3i0o3yVgz7HFpwxprOf5i3oMAB1oJGAVayG2Dwl0n
313/pI9IlacG93xUL4Y562FoLgBtJcZaCNf/pWD7cwRYlyaEy3K2/W0sekPWPJpvsAGgt5EdNoUs
L6JzxMdXh4B26c2BigizUemF+zMkvRD4aUGqilbnvVWfs+xdvxI3pXLCwEhDAFqqFB+Lj21RKrph
hQ0tASRdL2YLztA1qtzxUmCKivdhOOzhqtAeKuvxN84VKue2dFBdoUqPzaxvY89iaub9+NHHYd0z
iHVkKpvU5ePUKG9zV37ouOCLSdvSeA7KJ6UqdeIXQ/t9qdxnfWdISsmhCwWGcz66QzQ224LVItnY
KCt/WXIZuiZSMVPA3TeXf5LjzGSbmmJhsXt+kXR1k9WwMZFfa3fLduyU/vNU994JNajGO2tohBb8
kMP27z+7K2qZKA2AhTvFawPTG7Rz17WYsCEk83VN742ni3PrKlMxU980GaHS2f58TjWbBHrkk4i6
EOONuwLYr0fl1IBKSeXditaFsRcb6GVtfMpInADZfIWNwfSwq6Olu8y7k2p+wbrfEZDQ3lCwBRQU
KUQn76p4L6V/leq8SaHl6X4sNZYos3gpXwKa5Q8Vo1vc3KLF+vu8upkfD4jtJbDdr+U5T8QHRrID
XN1YV1td4mmVNYTradzMR6L5dkvJY5Xg2FBP+tqV7QO8weGUoxBou5Ggxx2A+oE51Ky4n6amxUeT
YxlsMa9zSAnKIhjg3mmjQ9DMNibQwCzqZ/9DmTJdbs9VqhY3Q7qx01ibHmuBBPgpKRJU8iC2+fy8
TObFgQvGIyk6/3Mym5aLhmNwiBB2dONhG4QcfeAdiH6HuFTm88d/ISepFKBeXmJhXTt/NI+/Hma6
332cWK0PSlsmLyF8O0FSAQDfu8KL8Abv1UjGtvrU/0wyDQ4Pb+yHCzG0jnPddU49x00sdmxq5eZK
oVUV4TGrQSZmttJtrQ8FizYiXMnKOwKiaDpR5ATxS2eMyPQZ/7+EFD20j1JzzWjw+ZQd5/5y2lJs
NV7vJEa50rBrPLWFWbNvdo7k/xcrxc2R71ivsD2mwaN0QV7lGyDjTa/hTu2vG9gJ/zaHkiX3h/bd
ZsuzXY08Cqtrajxu+mMXGs3JOs+VwveVtDTBVjVqkOeJ81ioZzPpa55j/pwZIFqa8mP+Xds8PSy0
HnQgiuC3LB1bR3lTT7NBwQpmH+1CoZ/Wd4cOBc5wqlvCZZtoi9uuSxkXnLx5fH6zPQwzaf9chRuc
AoTvWVxURjhsEn7Z0JfLYtFDr9CU8W49xPIKRH68H8OZXPJkER93ehU/4eM0EIGKSHbbfp9NH8ll
6pNyJOe9xgOL9sVv2s2wCGIsgWofFnDFarMLKwEOESlUuiTya/zloFf7KegV8c8+59lacAuClm9r
F1bX9JMopE1GUcJnE1kTqu/W5QOOnx+9oh4B37kWggRhhAb7Hl225ZOUMOTute1uezd12W0JT+9P
4901TUXV1kVHfvNSdW1lhHfsBl4Zy9bpcWe7Y9G9F79jCnBWg+xPWjrrYXqd257XMj6u3xxPUCE3
+NU7krNJYhWOPgyN06Z1rFLwwD4lYMbGBs0s+ZkqXyRnnAZfpK5J2FcXD7Z7Bfq9Q38EEkyzVZYE
P3TkSp2mXl2WQRUMPrIgvHx7kniMWEZKw9sy7s0xfW2ztuviJeiikvEzsOwM1AcidcdOSyVC+6C7
tNw1NCOwgNhWeU5OWYw9KLo1LNe/VN7CIl9nkpxIELeG2wJeNl7nwYdnl6lKivFlqD0Vs1ovnD4K
uR5E80zc0T+RKATMGbKoq+9Xn3Nxgft51rZtSZd2y2tbe+/3pKjlCrjKvWf2WGpLcZa1x4nZhho/
xWur3np0jxTjL6+Q3iypdmXo+zTC2NNf/OfI+2QiZJ8E64WiqMUycZJnRe7BkhKSN5kSbZTs2Jcu
krWilqiH/0EqxnWoLoEW/OvXVAr/hGECPu1KoawUoGBJ5yRFQmAbl9zUIOAJ87OZl++/CoTE56Ol
DBNQfokDL6QEC+zXareFoWO5Er6bhmmFTzZsmOcQkSUPf6GCZPeN6jolmSLJDpOLepudVj8OdZKz
TFgp7qaJyTf8uZLbDq24tfr3mmw2EiCquCK5bqnHh8fkj26tTgYEed/77BJvHTtTr83v3wo/zEAM
ZAzs+eZDFQ/JxgePZHMmp1JG4xHmuLQBx5Kia8jUGLOYtXOdDGnw8yOBrfnj0x1HHDHRIbgMGan8
01aRHsLRTsvAQRhGFOR+zdO+oQMrveTGGQNov1s0tVAHaAU6MzSEFxugjVl7+58SAtQ2yNbmAdvl
q6BeuDwyhh+hcZmwYhxwYE05qRaMHbphIlZb+qqNIFkjLGnAeXce/+Rc8QynA+YyHZyUkDR7yTVv
ciii+lsK2Wccy5XYFlMniwtSd/b2TjAUr34OEMg1sVpHgv4AF8xnUQJSZI2H44jRmsikLi4ekw2P
dapb+d3Nf211ROlCVYtNMeK02EVhJvZshKvxP5+0J5lr3yQfh2nRUPLDUbuzbSoI+sXZCfV5P1Z1
z1gJfAJ7m4//mKwIUtlnddetz56YmAXGgN7+XbAt1T5l6RD6QVmtEa3joR3JodqnlozWkkCG814W
bSJqSTev7L9pFtLNpfLrz/F3tIVG2hNwfmHL2IKyg8hh0uYE7vJXddxlPHltuQ76/5PaEfsZaKil
ko4g+zRAOXDS7b6ys1sG8PhV0DMOE2+gtUbRFrc39mOqiao39/g0T8/79+eGwsiA4en05y8IITGR
T+w9RWVvsAbs3CrkEGz9tELF6FNi+klc+U1LzNmrqafR5UDB8gO5QyluFRQMlankySJz/lezATgM
2pwXgV4e8X3+gCnVY0VuM/ZsFY5A0IXjpXYmcZgtxePhPd+ntyjlSpANKec3NmxIVBtaRfKmzBqW
tuXbzUm+tHLKNzb9GL8eBfTncMOfDErsDvOLjUHwwdIOln3ocC2joa0t0Kegi8BR9RJmjqWzmE4A
t+jmKaEntlv7yT250lU51xEUNpzj/r3yYNUfDeaQtE8W0bJdzgqdHTRdEkxxuNEiSe36jmI9w3nD
ct7rlPZtrqeYhFlm2CEbAxs6bgx8O7PhQLyedm3hFLxolCU0dQbwxntMJxKOlNWp4gkx7yJo28rY
BbqRI8RSZlgdu0EIiSxW6/k8AXi1ch2zPT0SZ7bmYDWdwpFt/jVeNkfpQaUWhxkaeYxWbcwsaKlQ
zXpM5LjeH3UpsqmjK/lHny/fBcMvGeqydZ1M8whyVi7sLh2aI+8+AjxRpikAb0AaV556KxRR2dZT
K2g4gvknbYZEHtXtSKznmn3vZhXi/C1LCQ/EkAAuvMySUCXdO8SIwFF0xvOzsdAtW0dyPj3Ayhhk
mWodE2vccIkt6t1FxcYxmsZ2Dba+Tqv9YLQxVcF4g6ToUZY0RUyxi4b3KFMo63M5HAu+iBl0NctZ
ymaGTKhKRfz/kXZEKewK59k8CUL3VmdCzr36U1sq6iQgZ9F0NQCtkM90rd6/D7JuO1mhSMXVWDPi
6N1mnl/32PCMXdOUJYdhNQ28n00PPrNBZOKTmwuOecekKB3u8ucNmGSKS2SmNZtf4qFZdGlulII4
jzvf5/c5MrYAEA1vv/2GM2SCQZeewyT2aUrf8plYDxm458/7aVp3QsvaeNMYJ7+NjCCgYaOIeKFo
bv4xuXc6LZiv5q4THL1t9kJnz8JkjbImztIXNXu09YuzZNC+C/4+V+OTsJc8eRFmyNo24m425+n8
iWuycGV2nY4O9xH/4AFiS1U1P3uZW2WoODF9oii8uwikeH+jTe/XRcGkpgl4PtfpqK2jGsJ4Alo+
M1nxCffpVfeUrRGjWJA0DyxGucB9T/A4AKg25+z1Z+EjKdENOkPX1bOgr1mOlJ3CgxDhlT7z6O9S
9d2So0mnqOiO+aKYG37kezaa8zbY/TXwT++do8XQ6HFqJqmUcdmvrODX/Ahr0gXSrHMyGc4oJLfj
jJY+21Jghqnls42hcatajfKhlztU1vqkLuN0O0DYUV8B/6l6isf2Zn+429wWsvlpeE9yap55iASP
DSumPMVuzUJmlJf86S9uaxiWNOayYQPzi4uRxFZm3BUNaMlJsk/gGxklreuKFIyrtMJkM9QGF1HD
FpF50EKnkqsa1DSEFRc2gqOo6UT6uZjKUd58xH2xUwOaJ0QTXrPwhDJ39T6QIVBGhDYIhdiSveOm
n3Xhz35sdcUrLT8+Js3NBHmwrpxfrZ0cy9UlMbVbERRW6nmO87aIzF4esXYBVvbaBm/NG5XxeJ3q
fbAUeB+U7Vrxu0ze+v7dL99u/qZahdazw1yQr4PUKd+mtv3s1BayWFRNQGTL+I7+AJDLT7S/dvmN
g7u8EDMP+6adEhQqYISOzv5/dZJ60PBXkFYJmkeaxa/gSqi8KoFuplURFjQIe6AjwPjNhB34F7IT
zFaVjqH6Xel9hyLqSDfVptPZh80I8XZop1u9T8slQOkuPW6+JJE9dwdwaB8spmmOLNjD7th+WK+Y
QmFr3uEfXLVKxFQHVKYVasdDMT1ik6hELgSX5q87Pt2eeHZEN2bUvzvkMV9MK/u4PKI9pvmRWZIz
WFEd9wuP+flyNOQSiOc/2QCkNNGl3m/EleGgaUQHZ1j89E/6LUt04UjAHvf7/qME7NaEYlBla18F
KcSa4n6BEeZC0QWdYf/lCqRy+8LDZVhJ85cpy0dxBcqQwg/srBnJ3kf8ZZuP325EEaFPeSZL73a+
dr7PLRjnES2MxOtRtJvtjth+l/UXsrDeQzsa4Gyy3z1lls343pDs6IoMJgFbh1UMkiEtresdah07
gHg/MdkOovWTwuXzCU5P+tZ5JsOwkLZXiZEB0/ft4Q5vHsr0t9geaZpI0/sXp0e5WRwxDhIxgNpw
yZWoZ7kM4ti/2Mv4FG1T68LpSsboM5RarVNhPK0eH+PH0afjOpGD2mruKe9WWGgz2ZQfuhc1KKds
byBh5eom5PWtvN8k406AZ2lEtUTgXSQPQpvxer7rhafDtdC3XwEwIQbLYYLCrmVYeVFuoK1F8uI/
5qxQfvzZLjW8pOZAy5+fAZwMbvX1RLvmQDdVrOOkkiMemeCQ7rYAV60tyRVTUAamr0hS1To/EdMe
iMk65O9H/pqfu4o3QN6wpnJ1aDuUcXE3UygcsbdEa/QDEOKt1Fa1a8gPQuy3EoCJL3+/61ijMymg
j2ww00DluK7l9kqVMvYenDAwG5yMnavTtAOTvhTAuHOQ/sy8hIADIY2y2t1CUHEs0QCNZLXxEfmE
HI80uHnJ6PPZtKuvU/zx2Si9hX/D7wXQGb6GdAvH1GeZbKGibeemr1NZKtn6r8bVf0smM94idwVu
zZxH3Ry5dpNblRnZD+JCPiwkSV+IhQgRgAdZx4dXkrHLtGduztRBIzkio2GYlGVeOznCPLUFBv/p
adPo1Xp7AqkjfszW6QNcYprr7ovbUddD8BPEODKJ+hg78nhRn2jOxT+EKLUn4I548d1ahfYUhBQx
WijYQEMS58FyLVRcg2w0Ilun5XusMbSj/AhU85sbK8KtSzGjwd4dQfjqdvUzAg/Jr6YSc4EC6hNE
xiUhsLFzunn3HMDE4jtrFaJwSDbZYDV3Lj6keHK18EiyQcP/phlYLkv5qVpC4+yqjGb6uGVHmT84
JenQz3WIw/GA5W6aQkSoA6yMfbe66C8ypOC5Rvp+JQCjNXnz6Gcyn0BuSSio5x6BzFWl7z9rMFnE
yS5dMJGKQ++3Oicjn5Metm4mqfix8ZNs6+JbnEGB2A+0f9EzNQ6+oqQmTp6kX3cVXIUUh1qgP5gN
Xf/+KVmI1e/gn4ckUonU91fA5GrfIlunzeqJupSUcIZgm3QnXR2BUuW9B3cgfO5CBNyXbfm71gF5
+arzv0DMAqqvfId5ho4FpmeiG8fgV+d2lTE2p2433RSUEZzteXJtIzEZ5a8Qllip1qJehRAlx187
C/VkzZ/nh8B7EV7x3SFgZUtW9QWczcLqpld7GNgHWvf6C329qtX5CkHyLTma1NJCrBW9N2EH89N0
kCImcac9TFvfc5JKDqU28lADU/OC2uYRP7NVQzdCGU0R/FAYYYdPtYo3WRHCpnyFuYsxQ40syC+I
C2GjJZ/APNqiYx+U2xdmM/5ciMHXpnKLEu0liSGW40aVBkaMXgP1zPyXejLhxoGSropPAJkwu7fq
2/GAwTcqRZUmmS20NRLSuPD7Re5T1pycOavEmF2aq3CzW5l+MQBAIcSKLfiyNesU71/1LkA7/FuI
sRIxanzNABSOTPOmv3KkdCfVlRpgn3MW8OtY5mZEEqs+poP40JRbsG7aMhZyMofy20eH20QlRZQf
X6nN963gEh6TdcDBNox68Mr/NDyc8mybhLg8nGTa+AzzhT/DlZHki8HfgAY7i1gKh95KlFoQY1Sl
hVryxZQn1YV74e93wM0aZyNEguxZIq15zOt5ldN82yYctXqbKA41ax4eU2Bs39BrOGxIPIbHYBPH
Gy37mmOUy0JH4CaEnJT1o9NT1H8n4cjHdrwqO5J6oZmYFI19X3NigkySXPNxm25o9Uwcsf3qJmpm
W2dg2DsJXBC148rmu8zDJBKD1SCst4ujCIcznY19iEEA88frUpAuxf9zd8Ec5I94DmUFGDyh5tSH
fN78BHd8NeUnnITYEwDXkqkInFuPmRrUz+7hItEBNw24T41rj/agbUWif1BGmqZiCsWzERCqX4lH
bJliUgDYkkda3wOHFw84faX0lTHL/vY/TTdQrEtLSSGkWnWguWxOLlD6ujZq3G+wsE9llMbnl7Yf
CT9WnO692PItIgxUzJCiN4wm/rgZSF/Z2PbYy7HWz84sfaA6CZgKfYXJgqIHOyxvhxG1TQJdGFrz
5qGkpnQApRg9VEUF7KP/AqsMVf4flrwoU4zQ5nEqhZE6cKwn3ivM8gbzB5H80FuQUww1/gMk5wkK
kiqFQmHT0s5w/j8mcPqxijXJm8LGWAvzgNZ5LnVl9Wj30vpnaHOi6+HjbcWiAQdWQN48Ja1Gy2N+
ujbojvdmvfdFn/7SgLAHmDQ6ElXHuA2DE2S0dctLZYQl5ojOUul8pexKck9KTit6IQ9dhz/TElFq
UY5MDyN8W61hUG2ghJdTVh6qkr8/DYnQjxK7m2ATrHz2LsRA33iEsDEoyByRFVRLE56cdjeD0u8/
RAWo5Zw7BX0CqKk/IMnwBHbObTc24aiwDOMfoECJHaOT1SSR7JVTZh/KL3qkkunQKHv77j4THl84
lzSZJCC1I7/aTvuZZdRsh6YQ2CGTkBPGHtqZqDG00AhN76KgEjOvDO3XBCq0fcz1ODfTJNPCDAJQ
71L2AimAd4kFDqgazZMCs3jqQWw8mmH9gVhUiV++QE06QgumDNPgeHoJVzitWu9dtvhZA5p5Eajy
pCiTrpBuHZvcL3vlBHL5S4Ydnk3QVSCElw99nYHHkk3adYMvuWi0svZo7DCRJdRAreZsXxyBePKh
W5dUZyNBxkjLesr+I+KHwA3y02ijs1dn2a+UAy1dmbrZtczsNPARNzNkqgRAiDGQ1LWAIspuh2y9
2NElRNe0M1adM+44B24GVk3RgBCinz1eRbOc9RLvsWc2VhoC0EYRX+/5xmThtMQz9vWmzjdnArme
qMUTCNG11IMxdTHdl5P/jcifb/DzjaTk6UmWXijJQvop22sWK6ixWd3Me+BZdclggSPzkGSn87+S
OcWCGc/T1gWGFh39kFtP2kCmWH70f/WL1kb2jQgP4xVF+fYijS9wlklgGN9gSmU5cUl23anXhsIn
E+z9nzM2k+D3jrY9IqQUvsMKA8Xx2mG1wtipvxYAbRXDqqjmRDcBnWeevjUUGLqDUnK4n4kWm9u1
xZS9tVSbZMVv81epjoGjrp3nvU/beqpXTnFXVGE6Zj/O9Lg71iXUz77ln+WzARZZ8Fw4ldvY+SYU
OgbYM+y+LmquDRMZTR0jkbP266V/tEpUWNASWLM6pmJC3wUErtQNKnvfkHGmFdSA7+oPM/7ond5E
+mg5Z5V1b0HpbU82BvXbrP1W2P7nUBOanKu4sBuwor0Zw4uS2mNuye+VkHDtEe5LWiOVaPLnO1vt
A46PJmXsjUz7GMsrKQdG74jvp6qTnCYleKqcQHVDFHNQGl1BunmXfeSTuiSxvjA5UnK2r1c/72TQ
k1y8OZtYg8fA63ZMm1c7C25popafZmF7NpwOVR2KOzXFo2jTlphWX4V/wkqWAaIKYdh7fu6gfFQV
By4AbUwRRWa9GqvDWSFQyWpxtScr1EMdBdvpVb5TFUZ/UMxzrErlLaA4MCb78Zg5LNjrmqnI0kwu
GHjfurBNOjSmM5kKoSXMOVS2b3JNY3AdMBcQfjUsKybR5v0Qbe7stle64tNG6N4tjX+Ki0t3ZSN5
NADBlKKhGKpCBLXzx13eLEZ8H2kbWwf0ki3ARDAUTOmT10yEGQxwmExMHNjVXDH07FPYSG7QgIVS
whHk1NBJrV9WXcWXwMNjYt2NAg4zUEEpxgO5gEejx1136F9XStiye94Cc7uxcQWzPkamCX//VwIP
KLlwajdJKogrb1x3g2KcRucclI8oqjjxYFA1Qae0JUfzY69rSzIL2LH03iWTkdivcCR1alfPvDDc
IdNxO8Fb5x8GyJ1BalsAul5JwvsZ9eIuC7gBRf3gmRPdWyMSei5tUM/DOf8REomPNiymSC2wJHTY
VdIQZPIFM9mcAIYwFAHJqRqpjUv7E6KZ4LUnMfyBiWGOAmkSZcgPA82swtqA/o4atN9yChACBUSl
VedD3R8f8V00oMtxkZUbwrAa0ayaBep5HQGlZ+thkZPg5nXy03GYQMWUb1P9RqLGAc2jZsvpP04x
KVbutxIyTplNQw6UEpcOeSYBsFEkdNzBvad+0ylBYFb76Rz5J22AOGgroJmdPGYoIIpLWsLIv+km
j7FCfhY3UO4NzAv1InWISVlIoDvU1o0p/XUJCevDhIwLCPMxoWRfgpw22v0b73junJMSkhQrLmxj
cj5jpbknWYOJ6WxqrnNgAo74DEABAlVSVrThvM6qmCmihbNd4+HcV5Ozl9eHs3AqxlfSXisr0sgH
QQQlKaT+extcHnITxYo4+4DK4vjSLLgvMd0DyKgqbmopnDFSgJ/Tdpw6gOuAPzuiixG5jWsbeiHn
raUxAfwwaN7NIk0EgT8eBE4kIDpGrOiDbqPZA+2o9jKgqUn0qmW3jeo0opk3pt5LtcUfDAyWhmkr
sfvTgoz/znfVCdoZJJT9jDZPiiQUEozxu0p0aKEpfreLTXDAKmRgJglQELzxSgKPeRls6+STOvx9
uQJaiHB1hX4o/pHdCX87IWssJoWiEhx/OnWPGlvzm8sZ9+0aWVMidzg+DtwMaDpyaPSSaYCdrJmL
iYjAUsOdUSMnc3NlM2r2FaAD6wFXQzXC8uIjGdV/s6ElGU3niFONYt7MxlTBxbYAVWupIRZgeZ/N
i0fTxMtkloPUdh6v6Ku/uMt8QgWI7BKzmOxxK1Een7nB7YqozNxlg2iYaOu7EbiYk3MgGsEV+RMz
U2XwfYT5+r7kzEHfqZNbDoHgmfs9FfPTsdvoBCRBCPMNhOFbP/yNx0HzuHc6dCY+h+NJ12x/UAtR
nIWI5EaaoOOK9wplxjBxidr5At/tmp3L6P/g62WVkwc4yvvLGI7Efin5oYgGR1+/JoH8xUS/HfQD
XbFkUoVQZv5nXiBV62Tt+TB/TsSWz5poL4+IPDKz3YG5KalUuEdFXhzz0KjQu5oyyWx297x9Py+W
VRkslWCo7QtwxQY/FLSIuPFHpgIIwLfKtPGOfW4nttqmCJma8ZFIj0YVZKiSHwyHmuODODUIsWzH
mjPZpToEJJ3knYhzYruGLGAvfUt1q1jooPAoF5h//vg8IEmNBgaZRuEbF7A5Ps/BBK8bOJ7vz1AL
X5gcb/s/DCZ+86ZvLxpVwwz9MjZWbEfdoDIPT6xGF4t1vtfFFpxKAeepPf3K/9jypC919w3o66Dc
ALzniCcAZMUwQxSAgUDtXjhdBQQaMuy8GdyN/X34h+WB1EFxzJopVp8o07yEyFU/PYm0l1fiUIft
6iPTP9QKfex6ADBTgzQOxxaXR9yz5HBQCgCqKfcAR9+QpZ2yYS+u8o296NiKyhj6A1JX2ndIcS1p
gpX4rnyYzYacYYclyPh0AHSjZZToJhG8wkbfIcg/v5En8vdmRdG70QGDifxAkNt2aV0wlDdZwllj
u3oeeUwa8A0xQxfwNWpitsW9gFBOjmMx0f8g5qzfo76DLskoY2gWZkuleXk1V4JBUxIx+hxVcPID
WGd4g1vTnnfl5cI5mDmo1RI6NIWcQ432+Svnlds+222OsBndxjxSIRhG/pIMXHEy5hKcYwGDm+uE
SWGufNqPWYEd8ydaWVDLrIkLIkNNp+owTHsmAfNMBaesfenwlVrtAVDTYZXDkqAsYZkltf/69kRA
d2+GBYMyeTGJo+FhbGNV18T1lSbF/UntjI67RD+1cU+sbY8GadbHESSF0/gn1meSbmpbtPBT7PV3
c9Bzk06XnqxQQRjJ/Jzu5ovVj/3tGdlAeuPqj6OBfO2steUAW9hv+Z9UlEoLEvYeaRgaHBLtFduW
IZVpC5NXwpnZ7l4act4Ywakoe77NTOCUvQ8kAXTVpWBNIBkAs55A3u61po6b3bQnA9SVSA9SSdNu
JqWRvk/S9QfDKHj7UGLpMBpkH6bqnCmlrcfVYrzDOr2TJNTBxMuAMN3dIRjd3U/ouS6lpXzdSj2T
G6uJ0AmSOy3hrF7i+LHykocLfD2swmEUYno+9UYprsGFpAR3VW3FFRzl5qQU0HfqHALstKP6crgZ
BksnfYvvQZFldaUfm6D1fZ04rvHkpwdyK99tPf+tC7WtrzJySiezrQZddg/r3sXnC7LDArVVtdAN
JX30rV97t0QF9YfdJ1cU9d87b4NLd8K3kDc77zmf05++6hAd8JzJN7Qtm627VQM/QHZmL5X/M99C
U+Ssi6lRxWbo3k5L+7jvywSbmH7FZ/xEhcIzp9vJHbpcIkvrjxhPvY3I3huN7JjswyKzp+p8NcTo
ctnwKlrX7cFn2Alqe43JjsKcAuQk5Lv0WUJc6iysTO8d/j501ilG2eN2Bf5neJjEbZUsyz1MPpMy
3AX9hIGQSUloB5kukLwRm7pU3vQ4ohzHLDzIK21kAFc1qoHVddtnua5T0ver9CqbTE6le50MH0sP
Qh+NZGEnTefEBHDXPDEuY7KRfC7jJ+DJGt578DlwGhhrEEL6P4jIxzG+KQN5XG20ZI09khbvPpwF
3tub1CbcimXd0U+S1OqrF9TnaOU5Z2WVTbgSNJUCpVm82mpPdJCVg1HcNKTyzKiji4LKtUEOhT4H
6IQIekRG6+eLQa4ZLk9HWWVPm2tNWu+kPpeFBS5/x6LMzFhqhtjvOD+H26FOzNCe5U1bFX5VOBix
HOoaKILHKEBAZR0Yy/Ff/t33MZGqllsgLCzJuwVJ8yh6i4kPsW2bNKgiy4+aLKhsO6kRyxOmdfIn
xB6gGg52/wBUly5+ioSUWRNJu3aS/4yWMk7UOS+BzY03e658xkUaylluF7QxNBAYi+5uj6+wJmgM
R8vTypt4YkCGwN3F6WH0dVr4ofHULPnzkM7UEGduVrE7ZAcmUlXKtcdl8Qo1EEEZUrGXvYsikRbk
F2WGt9FTtxt/2jeOBDREBh6Zuy5jHLu5tQanO52NZnJK1nVVlHo4zrRBLQ4CDouH/mJIvXxPnqnU
VEKN0tcBSbmfOMUdkveSX5jACXU6m9sgnh+M1CquHr+VIvgUSfcdv/c72Xz6NAo4yRFgAiPtDYw/
SfchcdDq5Q4F/lo9wiwAfU1kSj702BoA0VegrES+a3RspyuPKqiiRLGmlAE3P/tNPdOzkNSXepm6
xD6p1Vek+XBrBduqu2GXGhkryXgb/s62PLL+DIz+xsDLFBAWTc1hM2UFp6zkj7EV1exWPu4YX3WY
p0dIoA/lgeqhn3Dx7WI907LfulgEVuucWT1m3Oi7msMdlfEjw1z+r+zzDZ7Kr+QiVQ6K4+hVGbv3
arHsgLN09qTqh+zXRoo1QAlpoMB/HpLnOyijerk6MfE48CbHIUS4I1qA3Udd/ZbEPYWyMuxkTItw
Y/0uxaJ4TzYPt/gF3rHYFlxwVVg+W97iEGAuf9fXpvwwyilUM0thkP9bcCoLeaU9fP0muNkISACJ
U3ZiHyKhnMZR3IMdTG/GVApsgaI/jTE+pi86uCuy6P//OL52a3kRnKFk4P3122Raci0rBr11ojGs
TOM13dDjEuPmqikRbFNSn9XYqihLBcWu61AMyFNZmhgBU3zEVeKs1PJZ43t9AePkKa2EAmmHci9g
YKu9NGaLQTbmCPO8zp9U5sSPDUipmlhlJf2BcR5cb6bgtV8J6fdXcr8hKGFZVQomWX+OX3W+0hRy
e+4BvapHTsWRCC9T3J9M4wGmNzYeFMKcJ+WzO2kEhY1cfyXOsHBtzuiv645l6qALy3EktJMsEC3X
YnLKbSGDGK/LGgvwvCKzQMsROPIHgnYH38Vy1m1LMStcHu9pd3I1eQb8iRFWycQgl+z+WyMBXl10
a+1nykfVvs5fQQcWpLrTLhbRc/uJGG2JzLxqVyYkpS/C16PY01BJ8E0DtYyZovQgyE5A/lmUEdtQ
Mzs1+CfzSJTzkJmQJ9jVVem+3hTnRVs08cLhf7MrbIDTnUZhk3/1MO8qCL1rcv0eiUBPtMaNHb4j
SVzS/aIU/OfWl28bvEVzrRaJ4+ooBf7xX+DmES0pFUXTfPmcge35a6ZcgLIoY7YZ5n7ENidz9LQE
H1erp3iUHj/KF+Z4IVnDfU+rN7ylmfqdolSPeu6IcCg73LCzBbyhuHBkmWBzuD9SRJdQ5wqzS/9u
NZ0S33vmmHpciFGRaQ230hVhgvTrQG2Zrm5kJ5M0IthChQoB817NL4DHpPnFpqZCaaw3W3q37ebb
mr/KsZKBeg/sn7hsqCOe7KQaGJI/NMbfj6l7tJzQvhjur+NnkGkBtDhEIV+yORIiaTmCuW9Q5DLQ
e00hLLIpX4bZRhAA6i8yc4fqaRuVjMios4tWiuVY58FTd+nH/+zykbhlxdSGWWT5hZA8Ki87pnmJ
ghEmbi6HOvdGWQR+9ar6ex3IrZqOT8LDy0jZ/kmKdaMCkH18V5Yw5xSV8zKlCqpu5a4jF8vIe+L/
3xJGcCzo3q6hMweLTHDw7/BGBA+DlTbKWBrQ85Z8ljwi/KX8m9v5M5+ptprgZXR2Rllx3sPzYeOY
/ruDgUm3h9fbh8hw/d5+7kjfaShZlRE+rSw9+oMGpsaq/hss4hlmxaDOYojeL88FQEOJzq1FHZQu
63zxzdqH7IVznxDkafxPbMwtB1fQ6qRQdVmLpUtptm8+hjOC+k8d+3NBXcndOwU92HxYUFj1h91F
oOkKfiBMKQzm1BxZV+Wjs6hAEsz7n/LAcVGmZbCuaxgZRiuYFyf1MjSQCUPZ0b3IFz1Z3NzKNiIX
SWvWPYoMwTNyLt70OnGAQXh6xoplPPBpzR5Gw/lZuXDbkbZ0U2bIcraLJ5xacOX7WrfdmLhZe+wg
fiPoEdp7DFfJHyDD5Qpu6mvoxVMfiKK6xY0hudoNtad90GbxWLtVLchw2taY8WgscYkXMVDiq1ES
7PjW/Z/rbr6aLvNBDo4f3OF9DknNxJopDc0hp9nt5ni1eG3+9D2hshDJD/3uEXynsmxHYUN74Rtz
itYzjHpMPMnBgnt74Q6yNFHezW4ikhWrgEJt/V34ys0ZJV/mv9m2SWC3E/lj89saUYYTQ1NdA4BX
FQ9lAT2acbCE++RLNSumAVvIJ9mBUriN5fw2qsgPWnvXd37pCYwoWt2OQv0m8t76pD9bJ1vDQQv4
A2PlUdOZhgdgz2SIgZBcjRLV4I5ySatfE3v9DZ1SrhXG3cFKQWCeIxPlkT617yyehtRuyFnoAlFF
tfiB5i71xC5vdP7RLyhz6y0IwmzSDhjqNORL+e9cqNftPF5/FdaEl+/7mMyu4v2V/ri1rx/gPnXJ
thX2B4iqQZ0rFZ3aXp64u7wTBwcI9MHXk5QRTU7lgecghJY0jCJj2EWZUC4LLu5zpbZg+lmRn5Bj
HaEMUwfEOwHfV9GUtQ1UYYU5f6fGOnbdCOfZN97qcUGOxKN43Z7wyuH7yiAL5pktwiCYv7oBhwco
LnSg2dWNovqMmYocIW+XkpEhJzbBRZh2843fmUjo9Z09Xvawesu4Z/XsZKpoaZOD4sj3vH4rWplv
o+9stg1StEzgDQoJF44AsMN1zOrKpocSla5vtmXGna1deXQU1TgVa7aK8jrSInUiHHQbId8sZYUU
JfpdtJWSylbyR+LWLPvcRZ37o6daRklOpMuW1LNp58vCs86CNZtxPlu380tWdLsZZJI6sCeIK3iP
9e1i7hv9xte0tNcNmTkxZPjWcHVxMgSgmJeEVw8x+yqvWho0RuGLpLDhBj1JoxhknyHwe9+XDEEl
DIt3lWDD2AniADkdou5OqUpOyKUdhs3csXhs5dDGcLuZnRM9L0jEV5kmHqAoMJ7O4IM6aHq3uqdZ
dsbxessASOI0eMfiXe+4O9HEN/CecvOPJCn+p0wD5T1WvnEypbOZVJVQsfJCeWS7K+uiYczyeabn
8qORVjd9bgcmPTrmJnsFBcj7wocdglILQwhq2KqN0KEnRaPqoMnYZaM2IG5XGUdeX/1arjgs0bNV
ar3wwIE5F5L6xtFuCse12qa/dt30Q7puLUUSD8moX0GL5EhTEa3S0BedUNOfGIj/COl2c0Our1hH
id5lFpSyKIdd8LVeNWL3OjLCAMrimsvqMEfpM/gjoIRtstoyALx8vxVjg3kaDpAtHUj6t/Ouimhv
8Mlr2ZonKzR5E5s07RW8PXshuLRWeqFehUn+DBn45HYN1jdhoTtcmYl+/IY9ukrlPyHpIGzJJv2D
AhVXGIBef7pJjX4TUHG5o20eq5lOoEM5dczFnFXwxMwG0KnOWiO9CfrV4gmpFEWciMLRErHoiTYg
DpXOS6DT9XD4alOKOi/q+VYp8Y4t3hajz2dgrFwCS/Aq9DrLpUK083I1VLthL/tZ+bYg8ylK4u+H
Q5T8KBALenrX866qR0mwGN8F6jXXQFMtTLsVIgyvg41D0GyE+sLDQaB+Cw2/m1OsaOvgTRYGEot1
gUdwx3THyZ1yG4W+g9OIThg/bOMbIrqv4K46C7lRUQLQBhouwZUOk90sUvujhC6UFnrkdig/iZ3Y
q+9Uq1Xc6UJ1IEnxDz9h6Yfhn4YCi8vOD2kXGf8fLq+zwPV8wOW9oDJrpNKw2uAUVXpAsIU0kCyB
Noll3J571yyUaMCP5PBJExGjR7l2bsyPLBgyMwG+47z2uiWQVywCpsdzFJXdP8UT7zJ2srZdBJgH
ExwF6gE0kMcBTTwnYTGMvxc4ZfCoaeDNiTGkQRSzFbYEO8ebwRAnqhy9LKnX9jXNe2S/7T57PKIo
JSYnHzPwQ+6yzu9wJAa831NuYhyFhSr85JqBZZ8AiO8ufok3WoTZtWr6gpIa1SoR9Px08a2kHlrg
+XD+XYQn9HGZG1daa4Zf1i3jL8aPVAptG9SxIpwoVpwZPM+XNFELRh8K4iJAKVMlpMw6Jv8cGXyA
zJ4xnmDgI0IaxW+W/gTdib4I1abNqsJBpmRbp8NfFRqcChZy7cAUWhfIKnJkV3rxZBJ5dbsHPTAW
A/dl4sWrVsqXyJz2iOd3N1FCKa7+598aeHauqr+3uQLcFSHjyNkU4ZB5KyBY55TicT6yhPziVpd4
aGO/fNp4zZt4CVA8I2K4lOTW1yt63Cq3JvLaY+GLObEmaXT70Gt/2KHkVPHvi2zXOg7i+wJcDNBh
/nrE6TO8CSKwTxjPUIsrsfFgvv4CV/4H+IVSbjgSYmFCW3FcfievXGRXaWCEfPt/vXQkJ41bEGfe
at9JGc6sjGZ5f5dE7UO2+9p4HWyAMtxIhXFAOK1jffkoLgln+1h8bClpuoNa7wm8ulI27tX+7Q6q
D/2FX580AFRFQP0djh4u1kLnAxtyVBAks11/iK0fl9Gk0rKYdrKcIRLWiK82RuTMVusdceuXcmdJ
/Sue4JkumStCJm5WJYL28K41aZihuF9AwsVvUNDSzHxBVuqUP7Xwufbx5/21/b0UhusskArH1E4m
zOgKypwBaT1qfzB+55EgdiLjM8akyW9N+lq2dTfrLDdoWinrW2dUu4D6nQwA0REUuviMyKfghRpQ
HstOyXe1R5kN4OGYcc+LDMlqGukRt3uY33ZpB2AnR+f/Qpdd1o6QuLfpjyJ5tsposZCyEkwijCaZ
DITIV7I+jKaQ9+fVwzgYLYtMaqfwICJfC9f3Pf3a7yXWU8ypxPIBciVec2TWYWuOWa3H0X5/BMcq
oxqWiIyCO5GEgUW2f8e60ziR8Vr0girxl8eutz7IQ6sn+4BoHRVceGMSS/z+XPpD+EeKdYF7luHP
6pVlzWIvhxsRQ1QR5GMDfoY2p13IlA/rKdr1QLoZU1DtDljznpWVLSk+dffp0uVHG5DghNcpxO1N
EADyNkXba7lF4zeIlb2zmoIJz64cjA3uKuTSts/j9x+1w1p8rifrEq0dKPcG2WqYUiiDMzQwQZii
eaUN1kECGTXSvJF+EKV3azDqmwWUrdcTuCueZ4eRuqwT7nOZjH7BAA1XnuWBHAtiXTKLpi/jRanD
SPRIkhmN2TJLUCiChOaUKK4jxhrCE3j5dUWtZn3ADAls+ICq1wPasJVcPRzCmdKOwkina83AvQae
ejP89BmyrCEl3UQsaVXLGhm6wFUElatGt237CrmGiegTL61sTxjFHIcUNYcZCsRv1ZTeWpoZW45U
KCtQ/Lv3FQmFxYXl79gKLaLU5ScuUSvL9kImkPvKeKLg+KetZiA2p6WKRBIb7DXWPXiNIcOhgzwe
K4R1zkVIj2Q3LvX+J8aiD7ETayWOdHbof7opuuqnINkfznDE+GW/E602ZxbTL5m8cx434xfJvHTm
Efi3gaoJwyRLyXj0KD8yYn3fHzoYLnfog8duqmgtUtOwyt8ejRXRgdM4GrdLEfF+NWys7a90/X1g
hiNVdKJztimef/8DXglPQMwq7RHzPlmrOwrNE7V6Qjrpl1+ABTMV6Ptk9Eqs0ptimAGnAG0l4EFY
wTPaty/OyFv6PMiFcMHlG/FTGZKcGVdSEa/nkvgOxGSdhCi3/tMiKH5eWVsstcgFrXHvNQOX9vDA
q240RKeaMhtsnhUIHdsHhwRT3tN1kmSgPLGbXasJmYxYD+rwHeHvJxWVsSjhDTc23Nvilz0pxlaU
KBtMORoblus0iquxkEFK5aiQOqtMDeztrLVFS5NKH/GkSmwBCDbRtMRd7+jdJfTw5c+R9qTXQl7T
S2bI7F5wzkXRKxdQJwZVlwpWQslcQxklBNPWCKAnIqvoBqDUB8h5oqdqLwAYL3JZxAfdMqH53yQM
93XDmv+qLy6bG/QRD04Yhohlf9H6e4duwfbjEJ5ey87bzE12vCmJUjW/77SH9EYmzhYDMQy1TG9t
RQTvNLwzT79j2Gw28qGXXlxU/7PEvnKcT1uuAHUc+U26ERznOH0iiicdEWekvoa+Wdnhn0ououja
92qyFUBP25Xe4mKGNtd7Ks6VzPIK3P3SRKcsJ3uZP8cvIcY3P4BPJTqC/Qi8aWES1rKJWIJiO62x
Apo/21W66zUKjGNplwZeeriySWw3aG9ZAZXK/Mw6WqYy0PQ8ZbQBZRn0cetDL0SmlUun6aJjXtZO
SxhjZvnsL5VBZmW0fuUiymSY90Hmrxgkq+ZxBSp1uiL1xJq0F2yF5hKPtvRbR5E5pinzhki4mmbL
/vuRx3aDU7pUAFpElBb3+C07hKPHi1ZJt/jx6cbUBKnS1eT9EjGwhbe4WGfYIDXoRbVlPXM/38tp
u5/L0TByl3myBeJ4wUdRTuQNHKpZq7m3kpM3eEUaSgxGf0Qi/htoj3gtL24EySYpkOAKKNmuPaBl
t2Wsoi43cVf309CwB2mtMx+mu80+5S6X7bGrDfIRzIDLZIGzYyKuTWEOrjcTVqUOx2I2ueq0jVXV
GNWRmVVjICvHXH5GMUT01CNMw6yOgeGXWzDYeOT96KLzPTgicXbUXrM50tZ+2QtjMiulY5n3S/IW
tHWuJN+2h3VWQaE8zE9kk+8xGCi8H6utWmOJQafGOpZW72CFWpakIR/0jcLhH9J85KH7BTd8PL5S
mn/Bbe+x/R4QVU3vTvcBKYhErTaS6XzmFywgx/7I6y3tka5oq65wwWTEIkVQnQ9H+v+JqB2mAMMt
ID5MkfQP6xf/Ma9mGXNBvd4hNrwo0zwGtdzdfgH0z1Sww8LoSEf7FrSFnsMdOYi/UBGoydFAqysI
yvGQs5FpjYKSqLwKJJnSpv2G0nwxOKaJ+hkvRSPINbhslr96bsumJdU6UFAkvyWjYuslIIQhv8OK
R5Ue9jixlcoPFIqqz82CPfCV/WO4MsIpIyAeywMbwuSZ+O0nHheLahkGW/diPILaZL9y9HMW2z6e
vS0X004MvuPVa07qchTF0lQLQH/F7ab8nr/Y0DsQin86le/84/yhdrL6dyzJ/jCV0RL80a58pf/t
sXbxSVdPIpYLISdRSnEroCCU1Ped/tLGV/EDIrZ6fW0A+lGitwuJpnge0e+ChNjow7QB0r7hpodj
0sbDYxMrDkmw0K2XZOeUyVABWX6olbULnYHWfRDznMh+cdF7HzN0CWHfPC0Uj6rRkSF7C3wuVqpw
oATrM3x0rL/GPmFUY5v0sW7+NtVEO4D9BTJDNbXPXjR2/t9SYOgy2xf92EX04TNDTj6tEOhGKVeJ
V335pZPghZFkjwLYyNE81EwCKn5SDLdORYeUMbzTjT+eOH0q5rj0HJnoxR/rFmlc6CiAit2xYAnc
lQVT5kZ38godQN2us6GbV3g+WSfyPdpqtCN1xp01EOrEbwaQ0GTcDCxN8OfbRU0axOx4D6nqx1i2
6rQVfWncKtb+rQGesdcbaI0XH7OM06j8gO87yzvRsBM9yZ8ZYGg3o9qhlsXC3TTGLBYm7O5RrAju
oWltupDL+N2q/TKIAHk0PsFd3LI9+rSv7yxDWJj1kmqHgLh2Domzc1eL9lra/4QKUSGKuK7mtvZi
2Le6rxHEx35LgInF1dBTKX9FZQYYQBW54PqzuRNSAZA4RY5iICRSZWpTt6jWcHKe44AmNd7AflgD
66vTdIiXSNVI+Yt2lnwvmS84pcwNwLkC1hW1GNdHzYQj65mUxGCdAirL3KMhCLdRCqGoitRjzMlY
fZd0Iq8zx8K1WZ0loe1ot3BxySTVYzlb5LVPxjOd/ynL3m3Vn5BrtntdSIS11yvM2PUKhLPzKgck
r1479Zw6W+ftcxHuMC2s6Ubb1GtTo9upngYJJheOxb8HpMMmy+luVrrLmi0a9a+ppiezjdW6D9UC
FmveSfFmEij1nl1hv6x2y0QgWfj5xlf2w8VLBzUNnugdsVProJvO/k3nE/8MiYXHJcOqIP7zK9/b
AtlmN+FpfJGPBQjv/DwyHXYLoApcIQegVCjJmsfRxgltygCF6lJRCI9CFGGCsxy8NMgwYzXGbKvN
eSdX/bC/BQeeXBZMFBYLbUIjALqI6eVQcusSZ9CcrdOOJMwY4V5L7ChZnFBGigozBBm/zOxUqPVD
/4NEZdcz/8nPhwqbR8GmfSrDeyg2k7TIyJMosMawECdF31kiHT/Ek9fgpAYUlOJnQAg1s4J4L48v
BfHSGN84lASB2A7fPlQ6Mlz7LNS/RNxxdNed7KCOw18mcJXI2HBbr+Ccyf54yqePeLoqS17YMXwe
z6/tGIcY1CYdhWVj7rfDjxGtnYknuguPlEh5RdYnkpVn+/5A69SerGvKgRrULYoD0tKl8CsU7gL5
mI/jNqJ9AHUWt7IwDOxI4jGb1Fs+OKhoAsfT+jVvTUedAIU+lzQkvmyn8n8/aEV2PXiJEM9+nHrZ
nsa1k51JnJpG/hZGAKAKr4o/lnluSXXEzEQEGsOATo28hYUW342UmgI3MgrDkpQM02LZpKjazvlr
GMLa9OwgQQIFP3oHOzAQG626VknzjK2g1yqUnLAIjFCywBJYIU2u1fH7r21KeUpFtGKqjuOObWhw
LLKOudRj/Y3HP5x4OrRe+rf8wGaXmBtw9quWPos+WrzZP124ZDAIzkhC/O95KWLkWAPMgu66Ygcs
Ca//YT67VC9w1mxfAQgeyUuQjhc8C7jznlCZyBLlycBdVg5VvuCjE14QwqsDGB60FOajVlYeb6X7
mnckHycn8fmsXqc5yL5UzEhDQv3zHfKudkVOvoC3b1wYWbtlUoTaKw0aUYmJDi3Qec9SORszDCBA
42ngjN0Lo/Ol3CZ3fJx0l0+DS9v8Thce/y4bDRFfwMl/Y9L5woH8poqcrCH0rkUKiFNQaHumRvvq
w1LOU6suyZ/9b+1hnbBaqMANGy3l/Q12fM+cm4E9HQLDcmSLh9yO7gG0OYpfSgwyQdpxW138KuOt
uPqRnl8X4l9HTPNWdsuMlQNG+qd7uKb16efjpsqc4hGcArGKPmSbrpTwetddS7bHoN9DVbaf8gF7
VltU1UOfbQWRPp1a8gEWw4HdtG3BskDHoU7akf58XlkyJzCQwwGPGjc4WlNbh/hb42LuVkQTEtWv
0DzLBZytyMjBR6gSGEwv4cLqNrrYn+kUCxU5eALVHBOzmPDtrQ/BYiXWQ9gPqlqd4ov2DD2LdvuJ
FTGdHO+EiuUoRl4QGruEm5f6Hmh5LhY/mMUWhr7/rwDpJvPN2eT1UHBanlFZrWhsl14ilgBqdLOy
tmESSYPx46ILbWNdvHlaKPCe6q2g3zOH/f7SE2x29II9ugc2kJuVy6fwRDorjp2D8ztMAB1rj7TC
VRqykamWq5Tg6q+NsoJUejtO6hlLvicAv+XcjcagcWzcTJpkt0xtK7Lk8LZGWyJ3jBvVOn5U9ik7
H1pAK35NZv9+ZiAtJ2oC6Wd1FAjaOd5nZpVAPtkt3oAqyAxY5TwdYWhO6NLFriYYVKXDTnS/TWya
k4GLpUjRz1ezxWHYfbY+nnOkNm9bAfSja9oyrKDhuIVDKKEWdOIQIwQvLamaKNGSHmkva0/S5VLq
U6Bc3y9Z+o+VDU5BTH+GwqhghP8tlK+B+K9PnOVLiJLaerwH5VxTtThEDIWe0QTXvtYCKkOLxecf
PLELU2UkHhJURaMpj4dVo20TQiMIq20Fry5d6NlK0jfhyDAfyDTPtO8wB6/nbAZxEf0tZ73xPaM7
l+qQ/9RjGzM53M7QQxPO7Ma9w1mKnjOIxAlDjeTyOTlMFz76ky49Rt2BmKSzd3W8FV2u/OqGkeTX
HrjSwQ6EkxF/h2gWmlcQCEjsFaV/lo33Hsn//HGNIFT0KdUK/T7MIlj7Ww57BwOMiUA0xrfIvnc7
46gK33z0XBSmnPv4PVQveT3+yaLXhyhOvz2tEU14/GtDgftcjMhWOnVqODYKho+qW1YeJ2vBXdED
8PFpNZaaTwFhb+u+8nkGxANTYxBoKbMyy86gAN/vp6XTBZ+ieb6bwdFpJD6VR1P16rhd2BbVxua3
4q0S8C4r/87j4YHPj7jgXs8Q4tEhTucb1hIvAck/wIWL4yeHx9c+xZULSU8S0ylJuDnYX20QFSlZ
O+lW+fFDPJ2qU9HWbdNdwl7bT5fQ0VRQy5x0dPizwIZQV+B3I+AUFsD/gnmDhJgPb3d/TY0u4B7o
l1tUP1gSepQtV5jmIlbE5fzO7xMtqFP9j+1a92bQj9i+C9P5hNfI+Qxoq8wfv63zhe1ObDAeVsgm
RzFmQIau43i+Iz17KhtGdmUO63me6Ri6iAyeeADU9Wg8jbzv37LfP30EgSvLLD5ef4SfT4cWe12Q
4kkAIzvZWlNPO8Fuaam6xzH3459nzN06hRLqur7RiKeWZg46SyvwY+pzAUc8nBrSmYTDyYXIMjnn
AtluBiCHmbOr4GHZ+rLF3hwV5/XyvqzivzekX0iNF/HL0tS4oJ+qGc7hbhUvbpKXSPQiIV6JLTuh
0Tc6Da3WrTRHnIpWQTf091cu7GWO02hP3CIoRoC8yX68b6BFfl/O2msgf06fesmgJMcTXLmt0NHS
RIt2AaY4mIxNzjUd2mHVDulvzpew6XH3IbySeB1HdY41ecOJHOM91HabrrLxkQRJLHMhfBLRHNcE
Kae3TynNcrvhUghEd3iaeqWyHtuOXSmVhufKTGWycRiIjlmBFoFA7iKpfJKKMtlmcyXotdbpaIg+
juaKmy2v+FDmHd/gojX0+Klc/jDpEEBLICPtZOR77wROCger3Bu2zMZ3hijnuYYaC54ThPLx03ph
SkZ8DvF8DcauEiAbkUfNIjvdCGJfs2uOCEof/5MBl0pDF0TUhwkW4r/2AqSA2vURcbwaAu5e8CTk
iOvOni1h4JRYbRrKnA0Ij0rPojBTXlc37DKOuLVc941yijdrKyYCaPQBqzFHTv602xVMThAAynmk
yBY4K3MYhOFB7PfrU8IYQSZpKcIIDbgsdyJiN7koQvc6wmUBxQZoMdvMZl4nUH1t4bKbWx+5dCx9
FwHR9W68HRyYl4oaz9zKsUtnbZfSPvbEdnuddIp+agWppJA99QAvEN8B2/N7dtXRazdGC1QOkFd0
cW7y4Yo+4+v3fx9ZADG2xmDkeFzbacg5azkDgy4kK19lv2RkK1CHNefHlXmbGu0hw6qQss8CP8Tp
XasV/fFhdu2Pdij2+j+ddfpr1MW/Kr2qHjNzHq6lfkKQquD0KggDNotgj+8tQWvVT3+kKUiq6OOg
13ItQH/x57iSeFHFFctivjFxPypS2vyZOPNQbTIrfksf52aOhMH/2GitxBIAWPaYYVn6du89y2+M
I8xQYaJH1FQ0oggnL3VV/glF3NGPeD1Z8+XFZwY8CLrn7VFEfvz61bvUIEwRxQFjOuvWyI4/jGZR
9pKDkecK17cRiYne3SRgDTdPOQ6fMfSt4faDiTKSx+Upc1FLOVSmXRGBmnOMCWi/UbAJjfji4P5c
JRdrM0LB4fzLSyBx4dvnECXSgjfBJ6VDU8twzNR/3f9z7NEhB7k9rY7AEZ9zxnpTvewRdPrQ/OTJ
vVtTa5MyYL05t4ZhmS2IkkhIbRO+2ti2wrar86gjMQAxZGm/SG7dLS+kkrGxKfA+7qUvFXlxJ5sM
6dJclTs/fCXAcviKfOtb+TrhHBW84sghxboII/7WvGUuE4AyDlEx6M7IYfMtpSr8WB4gbD74h8nB
j4lrmmzwEOlmXscQWfPNZep8PjwREdvfL2W+zeNMhAnQJvZpB0T5M+aJ3zE3bQSKHf1Ji0F/PqNe
+dHF70D4WZpF0UbP+IJPDzj7IVuTUd59aOHg51fyMhuOAwXJqT6WJwAVE9xU9sQTDmOINrhxxZIB
r6HosLRBWrrWrXy5EQln4BB1IYWvGi2LOrCx4Gf/yBnd9H0h8536BEkb7O+hQAemOVoRSPVPL8nk
05VGaszGGVS6FU5GyYjR3XXQVUfctsNy375KzKe/k2Ht77T5xGSgIiMxPgcnVeDj5U8b6tiIJIAs
Kx4LUzzbr9KAUCMLiMQ15vQaAX3X7o+WMmTF2KqtSY/zvQO/xEaUGbn/V8AckNW5m/Ne/i11kTBU
sRBKqK2pfwpkGVly94rvQJdfKpIund4nyOtJo5Ki/uaqia64YzUaKhHR798xWPWytHpDWwtxsfai
qdkR8e1dPKDQyYG1Nwz7yqWwqgkbtnmcrs3ZvMSKzQdwFqvKFeSyGjho7ePJjigi8rSSL7kNTvjm
0xxRFJHzDXl1nffHorh3SR6aVIpyoVlqJB/MKULpnVYWgIW18QcUnNXg13v9QJSxbam4M8mGMhx0
efgTTEFDx6YBUZ1IhWo3y9lULMczBN/F8B/+/ULboKV6oW/9GLUUyBTaIp3iA5oivy+Qr0LfGoQe
hPXk7ibBiqHct/Iy0225YJASVHTrIpLC8cwcm1QVPMZBzfND9i/TJsjVS7DGFnofgG+BFFMArSrZ
jEV5AFQ+W9MxkNmLUF15arL4cYy3Aw93Y9AqVnW85ou6sCQz15QMRz6YXFqLGDpFc+au4DLfNGLN
c7jwNi1NyhYaabzHqU6b/Gbm2bNQYe8FFZhyP2gzVCzqPa+rI5nBgN0tY/SYq44P3Qm2/M0l2T1h
6+mphx0QRhk31ZIEyygx1tQQWocKk6YOzL3/A5iA47HHQJ8KiKR4IuuXHsaSbvt/Kt747mYf3nl8
9GO7rooMDbVmRU1kx/5tBNafa5qM1o7g66/QwmGf1VP/qeETtduPqMxsNfU6mQEprjva5B5rRbZ/
pBwTKgUIDwmZtceLJeP+nx/hQ/oda6Q6O8jPpK4OnwZ9AbFxQKaPCtjyT7J6sCbsgxK+aI+ggIi4
x437tWRItdx4pJAmaQwDnx5KBjLU40KHuUARqT0F5iK/DQySOBwAN3vbtrqACcgabYN9nSHflVIh
RseEJKLKKp10oYtmgtkvD11XXTWSe0ZEiBidPgp/iAYuBa51tAhH/Ec8LIwfxfIXHmH5M2LQuGGT
rScEdt8MjRPuL6HdKTT0XTadZgyzTbZ7lsslojSuXK/3ExA9l/YdOpA+gZo/JxE2PjEPD/HP0m+s
ynB94ob53BP6UHXM5MJJ6YcN6FDtd5PTQ007tH3k+a8yH4UcdkVJOQa98ZH32AlVcn2DdfZ45wyE
j9bMtgi4cjTwI5MhAwRGn48XPm+E2T94iDPE03CVUWvIwdYWddthCHbMJghwU6I9B6L7ZRyGVLql
ssuzmgnwU7SSNVMFcY6ufavd2Re0tfeuXa/P8ma/vKFE+KKTdrwywf3JyRXxPudxrE0J/2ZOFuE4
obZrpPWF+naMuOwnwZJWpfiPOv5Kmgv6s67zeaCtr75iJtMH2sqIfzD5qHi6QOxE5NmgjlAEhy6l
z0rUXW2kBGegeghomYEZL7/YLqfciZdLP673wr+4E02H1G0C+MQgMKDSdoHOQtVT6dWKibPfWe9R
4hh1u+duiUuHjyO68bVFz3noCwzwmmxmrtm0+zawKPGj4kU8Za4c/z1Iwvd8OB3kz70v6cRlyPYb
1R21yzrZ1zwAcE7Wu0jv/Eo7x7dusPubsnUD3cbmIapy8G4yqi4zAXrASQgfcVmPJ+MZxTWDq2Zp
VlJjfETz9oLoDpa+GT+PqWbzVr5ZUq8bnrmcZ+5cP/J2Van9sU1TLIXUt8dY/lza5xaT/xRWhY4F
fkxNhiKtEdwWvZ9PmWvQgmIE84mDBMSziBAQqy7f/eeHY9W4YuVnUONMrfcSPuWdra7zODRUnKLv
kEKILjlc3WYgAugwSF9TjERez4/trbEq0NA8ON26oF+QmThXMLIOqDrR6PGD/JuWNkyAxaTFZJZP
2N6MnJL07KcPH75rSbSxtxfbvOStyMM32TzdwIyYUpDCnzDrIMVInGRSloU6NKLlCWHq4ZLvn5PJ
xodgcQlayPlFkBmIu6aaehs7EDPe3ruheMgl4FVloltn3VOwZOTv2dRAdUt2S65UDX53qGkXYqJm
DSFDUQieHWV3LXgJ8VlEr9bb7vsbeTnzTGcC0Zjk7ZE88EJsQbKSeVRzpfX+v/5QExDnK/i4WSHf
Th818Kx9yrZrD1GoiT8JIZBm9nsJYUEO66brBIEMHTct3/0W6DIGV/HPxBdaymhc4/m3DP5dZ0A/
9zLmryLrMZDbkUorGfl84JcZVtvfM9qashHRwsfxTZuMhfE68DYOzxLRYDMpN0xJSE41R1CR8bdf
JoZIxmCOAJNIaYCK2ZMSMkqBKUQkwWqlzHguozh/hiXSFg5Xe5HTX3VEjbB9oe6gL9/dBbQN9W2T
f8jY3GEDHzjawcyxvusC/Z64rjt3n8OPAYtPaZArLYVgztVxMJ82BeOU8BvaNZeutFGlc2Q/ceMS
yMBUJRDThrqKF+ThRrgeXIBGh9DdlKSGWNMHzBC+YuVcaaBG9HzcX9MonCZx1xqpF5FMgMsMfBiZ
k3Iaftj/81/n38H5fpvAH0xX/95j0CJ9fzbN4lDR/2aDxtE0DU/D81njobG1pZICYgkIuRw1cVly
DkXCii9J1m2VHTcJjylX7onReGjvUky6AI/l6C19aKOeqvZE4ukvEPUZCW6D1tplgoI7PjC43GJL
4qtSWKI8JFk35djUNLZhZlay8WZppjmaAHYO08rgdfvn0bRzUPl3tmja9uVVtir0O232zOwfZmyE
9xBPhMs/E7clgI0e7zhjN7Ner/PL1ChyIaNfhIYIsttPcBSeH+8dIA1z+xQXDwyyM72aE4G4fJIX
NZCfgHvu0jr005vKJNtzjdMr9gGJoVeys9sZrEilal8/z0dCVcrgEK53xKMsZXnHB/j84eXM6NHV
V5yDwATFF11IJthNtpB1KXAmBqpyJPzs8b6Xo1SyMJJW+hLz8DX3pGhO32k0Qny6frFWvtHleCpc
FU2uAr8ZaGEM3KFulOc/MrW2loBX+y192ITVqqGSSKpeackEP+OMQnrQquUMqWRSJhwtbfoLTmdU
0lJZlz+KdwKaaQzrTLkkWZcjY3xLN9GMhUm8jXT8KHGUwvhugj2kE5MzD5jsXrTFH3Zxg5vohC9u
8828gjCrEEYWKaAErRt3iY39PKfxOcYi8Obvey7I3kNJ4Tat7KHnfxEw6ur7wxxi4/FztzreFfk8
5wLsnvwOngALp/x0h9UF8FJxHm7RzTlyqNwo7hMgKi6RQnpTms8KbfMqyQwSA9hW4jCuJBlo7zOR
zuTda1uNq/sNgt82WrcXeha0WnDHCw7IPIKvDdP6cJ3MyxoytLtiTAj4WMrvRRC6Cf7MW0TWwKBd
DGwnuJkcXdWLN8iR9YVoQMavScoEbr2xTdQqn+119jFOCfCgkiQeGpu0PGGzI2SvWeTKXZFflP05
P3Wh7d6YEA7WD39q1kC4sLOVd54jfGXAuozUFquj3Is8LS0hcrbHlV7RI/u1xIHIhjMqZUJ4SORj
LwzKOI4g1Qkf8pk9m6foYqD0yDPxFrNraUYXOj1g9v1PorNLPy+LnS2rRgfILSuMsxPe3+4TLAgw
XiC93+dm/ZdF9LDfIRpuTbBKg2lJbZnoHctiOAr9H58qsPWFJJrf1FzaEvE/lgM2hE67Xp7wjtCs
PV1FyuEFky/Dz3QkVu3hriTWNbXpVhze16N4dp9B6UeY+AXLKZZw3/lcKXTx9OF7WiOXEY8Wzw0d
eCo8FSqD/eV2fiMFcWkW9NIQsMlGJdf8B14+VRrM2g7euawEB7dFSqWIUw0Ma1wZ5TTFluBfCYGv
RY4PT3Mgt8mTNtfzr42X8ygjhgtXJii8z1OxFiAx5DZqiJbjvwCVAJDhdI0DX4KdNM6AcuVUQVgq
wa9py0kDXVxcamY4hBhpWzyy0SMhMWwa0wjkQkPXwgOT+vBA7hiv+5eBK4AzxVKhMZmmmsvgY5xO
YGtlEIXtu3NtAmZSU1FQdstVfHDSBqTCnd/6T03JW5qQG2ABhNhyZQY7WCN7CuFV53vxspALnz+c
4tpED6B5+/IPJJPRAWR/7tAShkih0jW3gHZnSfwvvMiSZe5jbKswWxran0OAB52j2IJsCNv8iiUT
OwKnvvfB6oqQzFy8SeUF4di22igKgyTf2BNhLKQk1yvynkmAUgq100hPqlTNXXx/eKDKE2ix50+W
QNOYvp/A8aXrsIZ95YznIcA7ipymBsd6KUthiDCHh/JJeMUNEZY7TZngNRcDl684ZGAKUY+iNIsY
ocRgWY52zDLBbQns3g1q+tGEQSpaaaaXisQeBehqGqdigNrb0tIJDJiYaXpSAnzEw5s5pBvfaAaF
pAgYmsgcXkB6osYYPqOjViliXVrGic/6PrHooiBUe4OhzYC77JyIPVerOyt95FLyIKrTn/0FzAea
ZKpXjPfUkIUs7D7mo8ZjApbEsohdC7Z5B1WOJKu/HFvC+8B1KtWU54xXui1VMMZ6PgEhYDY6oyzB
Zjz7yh7gmKDX8VJNxIROyKdtpvDHWFbeaS/PSyO7zabvP2Fg1As9rak323zzc0/JzXHiSHTgLVPm
k9B9mWhbyJeHv3Ptu+O++jM264Gvmc0ofeWGUylgQVnBhC4eCx9cuqthC9WdYgGy96nw22msDMfB
pjvTM9ZZ36iPwBPK8clU66VPIDIkuimxrqstl3POnJ7CKxJACt7IDUNkrPKxbgOHHODj4siBW3jK
mF81a+Wcjrnp+Fjclxyz0h5DlxqgRM38p1z3X2J0CK1CWcxOGgPIipZOAmXaB44rHsbwuEAHpFY1
KMmr+AxjMfR6va6Qhx1r1N4NBI8Cx1KMQ6dOcSFdh/NFFXNTpOmkOZF4Spqie4OO7qKwnNWh0dXE
eaYff3ysvtYH7D50gMqrlzag50qVwjD2G9SFjMI+wPi/3LcNcl7943jV24V1S+ZQM8JLFYKfQAJF
L+bNmZy7473bU9sKg/jNvBexq8v8bicHsX7PqdK8Pu5KS+gVtoXA50aXP8tigTXMf/u0RCBlwjV/
GrYWj6DIqEGOCT2EJnOy+fLzdRCtHfqd4UvW7woQLpixUo8juxw62ZsPWVWu4ntpTr2bCDUi7heo
Vj3DuccZ0EtQxfN66Yd/6WVUKK0HUT9aXv1Kp7/2JJctK2UQ3anb1vwnr4vS7hgqGXcqSTmh16lx
fl17VNgtMclvjxi94oXyqJg1h09eOaiLo1hQhZoEZU7UOleHvg96bdvN2XJQ7LpM1s0/blUfL+00
BY4V6lgcfN1hA+69zy2Rhy7YKSTZW/zm8nKt+Ixd8iIytT7Mdmph1u1fHzbIDnm3M4OSbKb/y1Sa
S8cI9V6V/sPdOoZOz/VZdJOicKFmayA5yVbG0dXYWrOU4JTi0dfmYHVS2KoJGZJQhaAO5ru/DSUs
xSp/UpAloIWb7i9vmjFu9tRSEjckGmHaHcSbUfOO63YhIc22QxpFC2JX3o80L3X3RJnUtHylVX0l
EGIfHeoZ97Rt9MZsJIwVmBoym6CkjRQT9BqAmQSwzFppY7u20wI34GrzA0AbcLYj9T6SBHTJK8jP
j9C9BZMi5dVeclqvbms4HbvPtPPugW31a7pk/Yw0wKgpFYz9I4N3tZN/+FP1SI2Wzc/Nt5mth5a9
cQ5ecE3MwVOUdyIOCH8M4UgmQ7yHCiWUfChjJ37gEW3X+DkJoMYSqjg+wbfNK/AuuqOtfbLtvIY6
e96dMoLOn10fkfROKL16U8EGXYSHQjhbRx08U09MNbelGL9cGhnoBrGN2LW1LkjMQRL/q5BmojQn
wbKI0VzhUzy3CEsFuFZIDAH1eoSuukwM/udLA0fPcJuGXR0rGUCcRlVOLIP6JJBPxjuCP1CaJMdk
9uulIs2xLdcQWmjBSHe7ykGodnBkHeHQraMyJORHQoDernqQPi0Uu9M9SSeLcG5Rl5oj1imGxNnY
X8ZhHhbpGitgfvOOdP96FvDUFmeDNsukNi+HBfDc0CYnAKaXo/JkO8IqQfcti48qrSqngf14IBNK
N4rJ23AVhovcSSeV0/7+Qgm3QeMwA+4q6TlmU0Z2EiNd+kSx8uPZRhCjauv5SvAyi8TGDevcV0Du
bKJ5r12JfHlqVhZTfYnz63Xh2xvcI/1Dsv36hOWJvvoSJybOmu2NWqUmlLHhxXQL9kxNZk5IFsCs
7O8IkMdGvKG2D51a+7+D378/cRuQBJESuB2JI8UbAKjaF+QPX2k7h5ptEoUuKp/lmIpf0ciHFOkR
Zv2+FvccqKrkIpf3Hejao5wysKZEGSe99ACYphaAX7ArGKLua4uO76+CDYjA4bcl2e4TOP73i5uj
JWP0z9xON2iYCjGhUSuJ3tIMrAFSe+o8fFij1quc7OA6jcRb5nyS2HUvsbOewtnetzRmEWskwsWc
j1S6/3nJTg0HW54OX4PoL/HmaqVu126B7n5u/rOeujT2zYTejQUXdQ1LS+n/5i5ST3kUNztDX8ei
Ydm4swkiTuuGabed+zo/ktNWkv8Zv38CRrlSqfiDlz63ZFZY+mgkmKKu4QLbSyd12WcHB8uz4Vps
pGEs1leTi6y3q9LHazLnDNs8wZ9wFQnzavWse2TgB+WFeVkKs+11LPwduqFSuRhZM3uw4TeOMZsX
iA7AdM19W/bPn99VhrpMdtv+hLZqYLgP6Rr6RWhMABuX2vASI/+qaa8M55Efj70TqFHohCK7rA1G
x4uYcosuIji395CGQ7tAbvGdtyjyeV8JdwNOEDauxjAlae/gW9Fpqjfqf1b6VoNgTT7NmTdo1NHH
hyO1syf+sEQZYasnRmSEtXCrsldeRAhYGnkhtPOLxxO0LDXYfeiNbdHxsnxk8TUxLTr8zxoTLvoE
JU8yqJGTDdb2NJWPzVHDno05wz35ChUOCwrcGkTqC0e3zSNRzMD7T3rqlp5a8PqoK6yc0hRbvdtB
7/+XnArVW6ulPiMXkmUQgvCgR46mI7Lg/q8+lmln9WBh0REf1NlubCkWWswrWll/7dzLgoTIva83
VfI8C9pRGohyBIs30B1tfP27chOxVr+d6FVYHZgBs2LfjO6kNqn+KQ0Vv8ovsj8y0FBrnQpgwMgF
AdeFu2lup4RKABiJBZ3BeaV51uwe9pmNszoqAs3BIuz1UYqsWqMxjSnmXGfTHjy/hEbT3g6SE69E
KOwK48yVYkXuBAB+VmVfqM6yUyDCwwC7NKXjapMNN9y/ZIK8iUhv9EUjiTC9E8L7KlErxHRwDR6m
12nqWG+v8ga2Deo/L8EpRbok91rFOSn6KhQ5SbOz3yh5YBwt0oF5pO6YWWPhfr/JnFXdUMSC/PZ1
0Bilb8SA5gOTbz16fj/MUB8qqdd3SR+V9OJazgFriF8vQI7Wnojw+Ocl5yL1P12O+N3XH/XQoXQ1
jRH94CzBIvUTVHy+lHWhlN6+nTHXDWgIYMm2rPtXvkUxN8A8RTn4yauMsEttf8bVtPuqKl8Y1WR8
xoEN0TRQfU5s8pijFtBWMMcF+Sox5fPDf0ENJ3t/AJ7sACVE2oTpwPZ5PTcCQojSWORYUfzgjIq+
STkFQVCMgVCLPr92UCEe0VkagE6w0JwppsEN29niGSc8wqb+LleS+iwbn7ALeHWP7sCWqL0ZNTIu
Fmnp1ZpCRa0RCUPl3qMRyl2JTlfz/uhT9O91fsFcMyfUwpIZdMr2l27M8zIKU/ur7HfPkGaJeckF
+8688mfszzTZmmfZS4fw+0Re3t2qJ4j5ymdTd4HDB30nfk0GiNHgKdVXbTFYZT4+gB4kUKhaZuRG
UTrvndqw5XtqRfFIxMjyaWeeymQ97s8G0B5RQB1uAsHYOMsRWQgva+PJaW2y0gTsKA40lpOcVE2z
hxTQKOwIBlGvMu92xt4BBUqq1LnO7SiBnfKHjohoyOLS2JsfJhDRpn9y90QUsRntIM38dOWmIU2M
kXWl3blUj63Z2WdIsUIan/cqZkZn+Pd6/AZnvTYU5AbIcPFbafE4ozIzJzO/a4de7DIFUmf19j8a
pvXzbqra9ZZXeC62yQuCdXUnuRINGginG2Eil5i0X0sLDrCVBhi+XiTupXYEx2n8g68kD6qJC0mc
z4yyRwGd0YjdyNgDd0fVtspkeBi6qoUo6N6HWWequu0IBolBosRDT2oZlgRlUd0+bBTeVR+xDMN0
cIuDQgNzzga7qo25ClPGX2hizmrrzI3Hb6a5u+AZ7Wl3JMCpkauiNXvvyNmlvtr4vY/o2FcQlDA8
FLQqA6j0Dirdufsn7cOGxs3JQyyivtV94MLqTNl/kwcYFK76yBZt/jrFKLs+6VknqlsVEur17rUV
hwqz3jQ6LYWh/xqpL2ZHgluwDOLczurdR4mTYKOZfi59TZ3NDvFX+6gPaQpwxqch60R+qVJmnePY
vgP881vHN4BvkZijGPGcVA26o+qr4/jafhJsWfenOt6mq6miXn1B4ARtOn63DjZUKDgRuI35mc7c
qT/SE5tDSONrYe+P2T8qsDpinsozuZAeKelZsxvZd+/EmVB24wBQ+k9dh2DF/DBuLi3pc2ei1+JM
THcjuZTR+7n7Zq8PVm0DC1eZKy+vnrqBSRDA2kh2W1+OBbyQtk3nfC4bsniIqKEDahDo1CSeyFxk
kXUDOpRl6cpRsdfrerWXfKQ2vHl6sivc1Yx4zE9SK8cPyYbW74oTFO4biCRERR/6vvH/zhYISH7g
+5/XU/UhH9RJRiZzYXxiKBnCuJlN5IMOMaUJTF9LizgBEdb+uylri4GJdqla9EeYeXkrSeoD2k6c
kp30ID5SY7zMOMlURuVLovc767DI29pAQ3y66TTPXSO65nGnV9/5v01a3hLTBtpIuVrKFYJ7yNdF
JjrCKTew5rX++oCcP1NVnJSsDu5pA0jfAVU7jsH2x+wvXGanscYyJuIiKvvCVYjlQu16KVyvF5SD
Et1TgZD0+2OOligozizzjYLKAWPqS6704dFT3RusRWcz3a7Dv89aLWUmjC52ElGjN56YnACW0fPA
iJDgnhu0RmzxRXBdPOEARuabzxrZWFQPyXaSg0kuZmanXQnQ+C20KwvKI3BfJcpwEcpRhX1WGGm8
MQT2zCoca10v9ZgjqUxyDfKijD8QAVUjAeXzF1x2T0+6lz9ftUI30Gt8yBvQfv5d/zmhIG2FJZYd
j2spwQIyaLiKvZagFDEtUywp1/CbL1qI9YD9Rwd99BlLRoQG4SI98PapnC+CHcm8tHeSqORdHGSa
6jwpjXz4zMuVgwz3DH+SGE+e17jPnjM4fUo8SiG+eddh8kqkT0wc8+Pj4i8BsmrVJ8xM45yn4mIb
WBDfwTnhVVHoLJUXaTO4ED2HmbCQeYETaJtI3GZbxQLpbTA7qV7E9C+gIxKzc2vNyJqg3G0I1M60
ST27j7lPq0XSZA9z3Y/C8900zltn+hWfuCGQ013HcuNuFPdDUiFsoYp9r7nnhNXuONNJPNjRsznZ
cm3zAfknhKLrCQLOV5Evwj/cTksHsFWWjA0o6nm9bgt9mLnY11NdNpg4U4Wdc4gRgk8hPuOVu5kh
hnxZuMDvfSqU6TrQsn9ZLlMUMPKRrOsBh6ymeErhxqFi5UDeJAQstAB9E4JjnnHTWEoOeLCuw3ju
E56Jhg/h+Y+VS77eGiDCcQbIFkgvsKTLrugI49p69bCNfP7Js8Is3GB9e54xGanlrOldi6Qk16qE
5oGTIsQ39bcuSb/HSdcAVvXwgxRWBHcx8RmB18BkWYdCYchEV0p5SE2ygirNRJvdAN+Ivdf9YpcS
axJIkMz6RsTIKPHAxGsI7TSG/W8BtEGh4RJTNKCGjjJY+py+OjVdnpm6DmiKBVs1r4odK3psF2xN
+hu4/Z05X4KVqR6BOlnrK79KVPO6bqAgXwIkTDbHvnj2ejg4Gwe6S65AqjkwMwMaBXKBWbR98u4b
i/kXVLkmP1V5PhjGbj6q+tGNCZkhvmY4KBK4wUUZTW8E4e9efoxfGmtrznUvVvUfpsrpH/Z5g2ys
pGX8yc3ASLIrXzb+t5pgQScShGaw9O57kInVJy0y0x/djz9fRPzrV4iLihOsEuejuE61LauPq6Yy
LJ258A61WFQSj697TjiQwTsiCrA2GFACrU68R8EINyAXLpRJrARZ8cnWtBv3XmWJJmklbdDAj+oJ
pvU2BXqWKU9imaOJRw/41l1FiZbR26y8yNgJdXQhv95RBGpunAqSNckhjiNg+ZvIzuTiUy8aZUaj
HIEfrp66MeXAmEfP51yZ36rp3Rs9mn7uCNg182T2wlZzpT+my2i4tvxNTUzSmjQjz/iGlSlr6f3X
T1lq4YOxgpgMWEpA3uOGSEAsM6UiFcuDD4wD0qH80zpUueIZB8aq4NQhh/0VXBCt5ocan/KPdRMK
k5RoeJ7EyLUY/qxrkvBvvMdD5t2YM9BUv3RueGureRhuq7/WD6A042ZDE/1xXQsdpcECoBwTT2yD
Gm1Ks+J4kIMsnvpwscxxsicII2ooZxOJpm8q/Dql1Su+GzXXWtvCM+q8lsA+MZppof1JNlkPk9s8
8ienUVwG9DWjXVJ4K3Jad+ouV0UE7t46S0uKdSvX3NeM7qLh2wxbxdm9G2O7Q9bd7y7r04coBImG
HxlmQ42krIaIiZhj/Z0NzmNetG8OKiXREBfad2POev4zn9RJ28zHt7RfvtSdA8dLx5SpzJBtEbS+
H1qpFeUNs8jWrp3uf+fDQHpZ1dZB9lbGyU5vB6qklc5R6N333y8VEaRmGmQDeDVt8+yo37U2ow3H
Jnw9DjsIx6kNli7mqZ1DOpemfAxnyEw3yxFAG5RoGe1FnF4s38onsCK6CbM3ILCVmc/vakkBI9o8
SsJkaN0M8sKApQtLGAk5/Z+zQf9QHIP8UEov76ZWBj8kApxfjshpNuB6YNFsBYBdiM1pCoUpXRtT
EiW51LXmHI/d7Js+9UKElgJQ8hfD7tM2qI6Y6n2k9T2teHBiixvE0PVo3lK14gSdgKoHkMtmp8qo
5DDy7+UxR5Be7OBUURO82XhFJdyUKM9Vzfwew0lbkgNVEvlZ4sAvPwCmnINph3M/6xbwQwPL76lT
en1N2aX2tYltokaIRu16ZPqdPvgYKom72cTJkeF+koozKxSlGf0aUDOu2sWnGrc9E8jsySejkWeT
ZxinCYJqCeSotIpHbyK9sH7RppCqcoP/HRsySbq4vKozdZXsn8Q3vqoJ9Aa2Uf9JocfqJJRiy5kM
jcgwH3GqnOEG3w3X5Hog9tiLtuqrwO4OquurhJ145DJQ36FRTWVA20u415Ayp5Q/cOx7Je5htNAe
4Iz9OXbSqFTo3wyQFIrtx6dffr2Bsud7Bi/lYAR7CBLsUcSSQKrWqKPfLVrGql8mba6X9QiW58rg
EVZEPAwZcMrhY/rIxM/WsVwXh9EMykCaWsvz/rpX9Mp53xaqRi0WwvFBB5PDQqti4VeMfsjd5wII
gmh0m4tCBH4n0GxobGUxsMHhAPsM250Rkf8o9CKMZJb4gCNBqy1FvoTmMlprWmFw+kjOHvXrcc5U
s/ZDwE+Dv1Zu8WD/Mh7JhiV06ZYtc5qtkEySpN3CKRWdboNoRjXJgaHRc8QCqduWClxmjGqkYvew
kF/1PP5VwBCGWL2RdkVhvFLB3Lq1Pxvao/UXxjUhtXFP98mvmSuQLrvj9FoNDLeMhh9916RjUJbx
METP7aQzC4Ws0kckGxEWlDglJmoedco47sY8TuPgZ0qYF2fhcfOCMZ/thywWGY4uVGZpyqUcAlDF
tp4y/YyRjoMrC8tmVBmFrbJuTmmKT03BJsLemTfUZJckJ0eYZZRZ6l0qZRLuXnvZT9Cfyg7uIQRa
CGpC88XsTK5OLck2FTCHBH+0wShA5p+mzrVskSKnG/FF+r2siD+vwmHa2dvi/I8s0k20GoIDb7Ri
MxZDEdMs5lZm4nZzbYIesEclq4Cd1tjkJu9uJ9FkpgHXbJVbPJcekBW5TtR6gDp/JFvjGb7/EGCN
FE3sovDG1YwtDpzAwWNHZpO3AB+GP6lwV5HXQM+AwTjx8dQkmn111JfqB1B7+S6kwJeqnxZSF11Z
jpEv4Pd/4AXAsDln6Aps9yfubd8EXdjAGPT4SJU/phO2ls+33xqx9ps+T8damKl/b0agZmhHzY+x
KnJ9h8+JQ+nUK6OdnmCEH+9jnGo68bQ4/CcgcG6MPrQoiAjb/AbWrtDiHDrnMQSAJntJYOPHgtoo
Ao+MIc4SQgRSac6T/J/WDukcWKw73cZpavvYMfVDm0JK+BfRXQT3MJK1cHyGMwx9VGD55oGbE4pZ
7IWHNVU/9T3cOBoO8bx5wGR1dhrG2AMiiF5vCieVtDLEhQZOVeC2m+fqfItgHURTh4P3ZHLPKhqH
no0aWI+rNsAGtfofy2Or+t/Pc4fTnDG1qqvjIPXOltvhb0c64ayNcZofVAICtpL8UZEVfjK3oYo6
Jz6sE61iQ2fMSmUuyKU+WUUHMX634bEa6/CdJhbd5WkTO4wR0qrFHmyEFhlvFz4U1CugBGdUvLAw
8LYUQk4lNelNNU4H1ICP1FhXvnnli6qwzO0pSl+CCbtyjL+4Jexv5xrZQkxlTfLQSXDF+UbF1rG/
QIJpLzmEnK4tNL0E5WVYbdnwJEabhEjx2ZdDX7/ZgUZIpTIXlVlyTut0eEzKCve2uGNjDcoPN3Fr
oRUsEXxcXZjCbtSjU3vKOkdhY7mmbCNxm50Wxjoj4OFYhNqPepZRtp1Q0BVi2ix2wnoz384K08/w
6OQCa4UokLlsP/sBrbX+CMLPW6GEosj86PvuqEK3f3I9YEIJABJQ5I9QwSH533+9S6Hz3iNp74x1
ozqBjQCBUJ2rqUyxXahFTsqbmLqgslmnta5TEHwyoAv24RUChGfRXP2cXU8SaF4pYEOUKA+2V6Zx
91QT70fzFfRsjKxxHhfToLPqv0sDe4qlST/+IQoFyetHVEqgYnFuFVdKFF5pCm7cC2XekFVie+Ff
hy9JLX9FebuyC4aQUBBGBi+W0EO8TXkflAoSaXhNN7x+hVCqt7gFW8gcHLOkMy1TKj9v8TxCHyHM
F+KuAi6UcDCdRgGFXDQhg5ABa4v+sQ2w/B3sbzEgdj5+eYDld5zERX/kSAqsHD292bNx+bYKBCvI
dW+RGusns/diRzumboEE9nHREYUaF8CGzCa41laZRBMBzEi9CFZMFHK0EZemLnKRH8Mt7P0gR/gs
gAwb9Js13XKEpyPOPwqdoWVSUSwtwo7j2AJtwmjSY4PmcBxMU5M8ZuskoCltngam5vztp1g6N6e8
qMSZwjGDuIOpC06IUT+fMIfvA80bY7KTWb8GuR/xxdi9ZfBnxGfywDfOlE0w1C26NyXMWOClSson
BDMd+UW9AtASz9faNdJ5AwTPLtyWOGhNMjHXaXWMp9hUpaZK2us1C9qQwUTXfeXKSbTH4OhzZuBT
ATd3SiYxkGiWMm6qKRhEr19PzSX/8UNZp7Iqf+I43InAbUHhKE6NaEbGTo8v9YF+TIb87zV5230J
A0YWdikwN2m+6pOwlNWrAGQS4MXb9BJgmP3WKOJ3XdFzYfm6oiT3ENgR8EuUuEdfb9NBk7fp4cZc
ryNWZcIDxlIVRDG0UZoEQXAdvjtQPGPXRDelJzUh3y2uTT5ZAVzM+Ex7E/psM0x1O0HoG1DLnaBY
YJ84O2TrwIEN6QlVVDYcWLyTq5lC24CojQ3cusm9eLDXVaFVbLuVMU81XEG4JeydJJrM7RH11QF2
FAeu7rSKPDVJKjSXQG6Wa/eUMLEfhyW8au/03g71dfJkvdIFXofSzlup3Hm8l84oW5gELlGqh7rX
wcLOTguiay9CVUQfTdUf+zz/yjCsLiiILftufrl1HzEG/AYHE6Jj3snQTdKQqo+rNOujXU04U2ZG
/kJdZ9u2yxs+X5uEfsRXvWyX2dAJQMj4OzhSuJNHz3BGrwErC8eoNEOtf9Rry/VIdKGGNtUDUFJf
EcvpWXzzZGHfPzCc/Sl+tlXG0A7+Is2utqSuZ1gFWrpVv2XpT9dgd2BPFLxRuOwBx3E06I5b3PUw
3qRAEkAVX7kgg5IDb/TlU405Jewvr9q/0X5/5OA+UHZ04E4pWvbpvBuYcXhtpC2/2itMPRa5fJkO
bpL3YRDSTXNRetqNMFzXNOeZczUeUBGVuevO5CLIDgu2Y/xfaGgauigTzc6d6VTC6n+klnY3ElLw
FAkYpXs7anT3wPsz140joMf+e2i0seEpCaQ9cSxYC5bTPGC/nA0rYhbdj3gT2rQGthlaEZ17lwJK
HamU0P0jnkQZK+9x2GKpALEp2+ENwfOH/aFnWCFv0SXu4BaKL540iKZjMt+DGHoRKkj/xQO286Fc
PbISWg39QxfIoqIoncdqO4lCy1swDG5PRZPY1cTRrHCn+5I299XoNhy01jCEEyzL7iYO+QZoF/Ku
n9xG46IBOvAaZGBuI7yHxtg+pvh3DRk5B01fJKzZYvluTwX3y83+YRLO2SYLkgVG3cjaYkPPPJff
ZPQff0oeVN8BMSx9mh9LbW9wh8GTfxgmDzM4ehVLkWM5paX4gYWn2FWgA5z5Nb88y4gbmhO0RRbM
K3nqGaaeFCezDpKQZw5moPJMdMIH8I1Pjx81OHmYJ4muPzECRXeWtaTCIZr5VV+lI63a78B6O6jo
sCK3nO/E/AOKp60CJbf1Td9oY8A8X9wuaYclYwwdEDmRmIT23ihI66F4oP2DFSAAjLDmeTzNUCyE
31KV3VIxrzQhofVdOUFrI9igyM14RdCYsA1jaqeTbkqav8TZEl58Pwr7BQbplpgnDyCOkcE6oiIy
z2nm/djqmMJr1RLztZOBpko8z+8cm1MgnqnRMSNlmwlvN14ZtsEQEhxxhFUZ/hFuowHSNNmDlOBr
iNfNO5RFDI2XuheukuEqwlEWIL041uiITHmZn7tRQwl6Hcs5N4/bxciOnOGT53flpuLQZxov9X7z
OcD//5Hz/ffw4qCSoH9OyP0go3gEjlf8WpNQEOHtb3lIHWa308i6c6uCxt+Hpsi9etFra0cwB/Yz
lRoElwSbYchiCiC4dnF0+a4K3wIietTlIYNVT4lDMBt3my+/+yCBF3ZJo2GyrSMbnrkzyfICLQK1
gqPx1n+qh0WcvBYyasrcga/8g3vBVktkCq+AvFbs6tCrc7pnZlXMsKJ+JT7qJ4G76cn77zQSrC3q
0EldUSn+TzVak88I8mk/G73mVUZ0dA5c6FBDHTjWt9SJSVnb2WuNCnUA5qzyDcWjBZc7UaLGGcrM
RrJ1Jny9Eds0VS8iZDK1vlPwTbsbXBatVJoze7RZTKaR/J/OdqJpuPdAmk6KMDaXlSnLPcZDN/Ko
ZxqKM1fIcpMDK74BZ7WwoAkrwv6eLVMO3s59G2Iymv0yuIIXuy2wL2Y8k2CGKrHiYo3sTsibTI8T
gssGf0+jN5xT+dCRdAqiSgZeBeSUifma9nKDGgpoTvjRZFsKfsTMyWLz7mvTTZNGqAQZGe9JI9O6
XPgbZsBYSIK1cqResKLnvl8KT2UslZtEcX7OJaJRpM+5eQF/X5UpociNjhq0wGvq4UNFi9PSD3Pg
bcaRXGyoV+AOPeLuLqTponQzu0PP6VgF5FCmRxs3jD8EvB/EjuMuzOyY8zWEH6F4Wb71geQsqKgh
7H79Q3eMVSEoj3F6Q5rDeu3Fr1BfCCKoboLINu9M6X1ugXT5t1s8z7vg3sz4RfVydxc6bZ3e+Rm1
VEA7cJDFR+X0Wdoy0qz+/2mXLGxCFZkdA+wZv/E5+TYhqyHQdhP9/K3z0aUyVjzHCZmUd9lB0+bv
8llZrdb1o8fj6C5FFaiVALKLOIq/ZTdhG0IvM8FrXCOxnkVHcri7RPX+26JP9hfM4THizLJCBuIm
FEaY1288p2lnE1LsQ3ajdjH+Zf/zOxRlqH+18xaL0UmapWe9nQwQKHhqENMchfCsqKaD6GbDGvm8
LkXzm0YQ12ZV0i8U3XVTkjUkl+67nnGMh8tbwPg2G2b1rdT0nXMLmGCPLN86+sjL31IH8jEPpX90
zW2vlrkcj5QOzcvtPWfgsG7qCMsJhx/ykBCXsPi1Cv2kJY/OD8Xv3ZyOBRp3V7tFcihH6I9I8YWM
wqKiQbdYhoL9QGr47tpPQrtj5eni3pgPfeosLHk/YpOOkmzS42M8wEPSZblcYjx55IiFUf+xCvts
7hz8z0Y6w8fTuE7rhJEXWiAQRSH+jbvJQ5r4ENrOqGMtZug1/pQTq/I6YR5K+fOVM41MpzYcEc9Y
hsr6MdhiZG/DIycmvDkqj1rL/O6svNyV4UkS9BDGIudJjyYI0cFHmo25S7W2EeozlJxEVkA+nziM
KlUjCjpjabhZoSF77Vtk333nGbQTPjt1AcWHjyBypjNkO7H86VcXxP5jvEuXJEOGMDiJwTdayIUg
jPHurn3aXs6Ji4yhAosBn4vo7xFpksH9xSncWO3O+3Rn2TUjKtM3qgjU7SFTRIpiwirXTYIOBkqt
A7o9CY4QJ49iDSKnac8wo2RKs4ddEkB9I3tIx+YZAlwuBU02D839WpYkLrWzBn4oHtFbdkpCslUX
S57sW++TBtwJKNNZ3XMfSpaSlZBnSazqmCSGU6UgNZ3HtEIpAa9tRN74ZzQr30eWO9NPy1okjg2B
IF/dbxR9pXSS29eM6fa+dp3alCQ5t1WBDXvgGk/aMahPtFvJXegbMIrIeK33nH+z2rvdhYPY3/qT
VqoFk5o/FMFedTOchVE3K9+wzq4vJXNXcDF1/HkbnywNRpi2VkhVtsM9fM2BfbU1RXYwpGdmpIIa
qbnxBTH4gpfs7+5AeuEyyONYriA7FSSlfvW0WzN8gAd52LVwtQVqY2+ZkzSNVGU/wcfTC1LJN+qe
VKB4U4eUbo2UZyi0obvy1PkewM8Yb9Lr5q5KRQ4ioKIuKwcih47/whdeMn+gKcuXaOFPlP/9En2n
ZNwpy9QbLYRnRPAlkHOvEJnqhR+/2DM2g3/F8h9nzuwHFUelZ4MkVj0lDLmx+9aT2jlX9ZC1LoQQ
wfPAyuSW22WzFUFv8RRnd30M7yNO6ENVPjlqtbSHyKsDcsm52GkSloHVwSHYYocVATp7vFAFGAcX
msJSiBernI2IKeYAVisD5SGr+wKGCbCDmGsCaWrYp2f8jbN0WM/lx4hTNtmUhcfYI+U9FXat3gdz
v9kUYrQLhsgflaaQi12yT8YN3M0GyhyLW50jv9yNuAU2l9h20fGAuT/pAybF/IlTq67Gn66/ayUM
z60rwIkgHALVg5RhQj+5y6MO6KjyuyrEMy6u0OqUCTXiYfaf9DEPSN6OktOI5H6ND5cTGO7S5WU2
wE8gfCqzdl9e+dbMH2kuWiNbwtBy3V8taKQuxFyzysjpUsiwWlAVfLOtjx8QCT+RYt7R6/EwQybK
2BawcmX4oXg+jgM78GaIPolJBWW8rtM5NWhE4WtEj27LeHGh11cAyZ28H8C6Tuy07C/XjzYWh0ZJ
ios7ruI3NuAyX6e+OcUCnDzgsHWy/kTDpXwwxPwlKbhRYlJlTCkWoWWKxebHSykpUyY8kjfxeSKx
RqVsgYPxKnbeiOoWPDFqO/MQarK6E41FvxmYYLcourdsmGHhj0wDKDUcx5B1a1mThipRaPgCddPd
b/5yYcJP4GNmdDwykqbAFC4OysiVF0Xz9nQelyukerc8FUxbKqSa2bDefBvA4sS/ViF/0HuLMyd3
m7TprgOJW0OTUdpl/J733rMa/X3MqVJSEcYd88Ec6LfMfYSBkRtqCdtUqFyz2nnU+gICgSby16Ic
X9NVS2LhpyNT6381Gjh0GGtiNL1g3shf1bkQZnPpkEoLloJYvQeNdzILeNZrfdFrsnhyyT7plsB4
MHacVI36gU60wU2ka1czJAK8XXCfsbPdVgLHcHo6fyUM8/tmRu+6OVXcXEt8EUiB8SNkXib31bW8
rHAhGyZUx1GJHilIlTzqBw8GYUyzHa3Ah3UUf3fIbRzPnuRnbVsXtgUAYr7k8FK41vsfNT6UwxO/
9G3SZbCnUPkRmUscXU5uWScDHRZ/7dw12RpVy39b8sH3mJeSH5X3Ut4+YqL9fgYak+Lj2bCLMZzI
KsqvnML1WIsOnDEJcgNXIRlOO16lG1lTSUM+K08M0fXfRlVJNPSfSTc95MDBz4imeCLs0KF1Qgfm
kIU5FKV+7Iq0VNr3TqnST7Dd498xDg4VRfX9B82WMyzfaqVkM9yyoXFeAH7mfOvkNisiX2JgTsQW
uKV5kdyhIlfm3FjSeVsf2EBqU5siWS11XdelwMDUZgIZzCXa5WrPQGMaqpkdMY1kd9n+QUGbkd1u
ogBUWnJB9B6YmFS52GmktFctkS1iLPxBPmke6LzOMmQRgKdqZgcBNHTNAby2MN07MoPh3ZjkF1ro
S+WuDc4JJ7rQO4dD7Pu4SKMkfPKSCRhztv/l+6sk2Hi14Yfr+X7tbvaQ10ovQeOf7ooFL4p7ciBQ
x1gYMU/uyXZDgMEZ/O+rNcqkkyX/uGhqGLW3YVDXqM2ADLpkpboXnH5qvUwFEb9N3btVGhehnxR8
m3BsBW8JNpImuk1cv//xAGIa4m0uk2C0NL+jJO+t6MfRkHcsTLyf5C6wTs4DC+nuiyWa7BK+B+gy
DWDyc1h/9RRahjC8fJIx8FELnPkvmEPjX8qakBPPeSlRmlSjZ7lgN682Nz0x+jitGbMXuGcmLpC7
J4uCK8cAh8LJQdWpfK6jrFkfou+4q8AwngizNfgChU/uFSg4kGlbtzMoFkh26geIHZ3P4dPMRukR
Qr6KZp7+KNgSP8dp2qxO1wDnABKg5YXWMFtDl/IRSuJZY7gXBrRPizoDUa2H9PiCV8cV0canAhrv
aiVOzFbffJHb24jCe8JdFM86prNHab5hMOXFICjClDzmrKNmZjCQi/aEvsuM5tgxRnIz0QdF8q8t
UP8JgrA52FwY5XF6gCnfXQu1qcxFPOePcx1klqdO8x3Lue5TSrAR5EFoBfUX6xolCj9X/T6EtMhp
LrvSPRfxfS27hdtIewGGTS+49oylN5KreUZI5VHwJsiiO1l+0jof6o1MmsWk4qfeR9vdZy5TqyRQ
A2YYoAMPAAUgBz9FwuXFXwfQG5SvCBkZA7EmpLBhud03tAPpcXQhYytE3ljKCuoppqwd1qj/TLP/
4v27OUR8kVP7ONmbXCRk5LVEWgLkIY1CONLQqcXIABwqiohhzSz29aEKkVJ+FXV1PhzsBZxiAWEK
cGZTRIgEcwwb4d5khsr8/dKO74zMKPYXF6FxepZbzYNqqzbmLoz/0jxp/b7a75tVSKpJYzCkwMxO
UNgvbyuLMFNnfQlnaZ2xgnIsCeC/6sT+5K5ORyG4ojsK2hsVr4kIsu5RONlh0VfpxBf5K6EQEu/J
8PfQFNgwAGhg6zaO4JTabtwn4+XNKDxRtIcamh5wKrq+dUhOJ6EWFrTuzz7oncEPM45LoOArkKfd
TxuaU5mvZFvgGHGrGU0FXC/qwJVhhJSxRxKlVzDYFkiy7KhLYswoOZOhVMBPTFfqCfV5+jks21Fr
Nrhxxv1vkyS7Rfxgvb9POeqSFWMS9atkosuTX5jwMd3oVTmvt32QctDAR0HZOGg8KD6VYOdxzcL7
aNtlkn7p3Hhe3nT3OASID4JfLhMzEKuOObAHb614HeVPieJNd0u0XGA74fAQCOqDxXgxBJ6j/RE+
JOy9QLwhrIpqJHhAerAdytmYDAkIEHCprZXZ+VW1L6TBtUSLrnM0bBwwz7Fcv6i9J0zrwFpSUyej
OZwc2qT2ktVogS9xtsjBPeHOueU685BwWo2wb23btuz1bB7+exZUuWq3OWWk+AK+QMk4lR9LTX1z
q3hxY6N30lmGv/NpMK8Iku0ozG52fRD4zoTal2S6tkCvgl0tfM/DUZQ5XrEuQC312L0V6gGtQhP/
NJRGywEaUDNZrcEbTLfj4rvETokzcZuq93EOsWXco3RbQXKHL+xIo4LG3NCB5JWJzu11izalefQJ
cumhXs+alqTUevnVd6Pw55cDVPx0wls5k5+2y/2y5SEtRIUhJmb3ePy8h7yNwJFbdG6UljE7IXkX
r/8npoQxOB6A9vnxcTAj5soMgY3WOIKma4QR4hTK1Yq1/T5GjE1+q1UiCWKGRSIoiqLAFunKNcyb
ICQxksJNslQ2LApZu9vUADfkY7BPIjc3b1PBKpPpn9w361gTQzjjwN/6g5IGgM5kfNb00fndzK0f
SHTSw+ngwuqISwNpPeNL0RmA3tbvmTycIo47GTF4RIbonpvSe1Y4hiGNSPIbMtfnP+pDHA6n/nBC
WGTEiO2u7WSJSvXdBopwtbUC8rg3XYUylaQmBL6YKQwd9K3VnOkRxsfcsBV/dbMJxR5dDcSI8mEr
vb3ddcgp6lBftD7jKNoUVfcdj49M346Pmdmn75hukCiRT5wRtpm6QYht9gh57xozpndvT3rPBZZO
7H3cIH6O6TW/fjWODYbf7Z77SxPoL2UgJN2qNRJGAA94tFvzHtZPtUK3ellY3gBs3Epy/vDopOk6
rraVKb51R2O+hHuebKf98NR3fBwLMjURjFMx+v3RYmsNpsg3o4t1PHup94Ml0PcYcaY4tTWiliFE
tUl/x89p8im4nOl/0CI28+Wi/h8ktsAT2ziTZKcdeQMOnBq5NokxsIAHzjaSX+EB5lLsXpNWwa5o
OSmPtlfXAS2UyihwsVSaxPqZo3WqPlwoWS6G82NrGWMjENsf2W+fBBWIIn5mivQtCbq9FW7VLdUx
a2S9TEHVDdqr7THdY0b5n23MMLPFT9EISEeu2taUfG3hUIr0JzHmspoqkOdykEA44lGzWq2uKPOh
pfvRTwNGG73pVHF7sJEy93vgrJxuMVvqVljs1OY+QekyKfWkJMdzBPdfphNGUT6u8zUpxGdBbiM2
ioFwdKHn0IQ7ZMOFGjWWrJEbkLCgZfpV1WmNPi3T07PRCZLL67UsGE3IiuKIwgoZR49kAz1bgzH+
beRqmo/m23m+0eIO54tivoHLdESELo7BXpbMpDiYjUQvfaVP4ce3u+Ryi7l2RbuEOZmK++1bWz+J
iXHu0Q2oQMx8t1crUoRzLRf88eil0sxFgRYExIUudnrg/0sPve1BbFEoLoMdMmZcvKB63kCPzhUH
g1tRYRMAkCTrq6HT2cdwe+XVC52BfnWlYK4cX4w7/DVjnkLQq98fPLY9+pAZyyeza2835GgDHYj/
JnKbVumlqCys8A7QJVBG/m1nLvLk1K5C2R2M+v9dwMUPFm9/ph6+MOaN9Q/tM0+Md5UdtsM7GIn2
LqCRhFAikoQQYSwf2X51CcFA0Hm7uZ3bU2i2HT9vmWc9eV8kBi1HSM1Nyq+vlLcdmfy6P9hTtBlb
y+oWtt6mmCEeIwhV44AvKMWQFmLtw/FBEigwJMCVUIYSL5s1b5spP5xIQ9OHXq021XTU+v0qFWAH
7moIoTGU3fQII1i/CZd98Q/p/XoyctIlltrzapvF/obA1xNA8FfdTezdi3dt3gTI/1uQlzmYpYE1
Er/8dPaNgdCmZUgiRPISKFDcu3dk8wY5yYNp0GtdLcPdiHQsuhdcq+oUUTguD7uBhZkCDDXeIEtz
Yq1WtBBGlu5Z8TWOZMP9YJSAnpWM/mumgRJro1X6txDPqKJFtbE5hZwAzrv9k+EVTBw9qnhIA5cF
EPytx3sxxb/Jd8cnL/emntq2yHvV4QJ3HltOKEB2VyqbcW3UxfCen8/Ru4p8c4LcZKB3MN5WasOL
6m+RVG3/5sfXeRBZ+3RpAEEFyCBiLO1z2S6WnXq0paNKzYtHm9HN1DsCAStzV0t//CXcXNWZK0ul
mDa3rxFSIRG4WIgCAmxtVcplzRsz4xph2W6+aQWD/AkzGpcrZmsa3LDgxIg0lCkoucI3CxzIjsrl
IdfekrqGOYy6jBNM3uTtjma6/lvQYNNbsf2bSvwnLdJ9Zb8mTix943SitU/AytXPaPdHf6gc0Tuk
1wvf9K4R0ylgavhs6TNARA/I0XHJ1wjPOjMOnXrOeH73p+acDiTvtV75i/SV2yV/bzVaeI90FwvC
i0Vut9mFbsIS4Ar0pLe3sKvpXG/crVOM9SzSkKQ2erfsWKRqHHgEMCGdwfEJlsyLXKQltd7UPASB
3xSAC78grsv9oQ2jaJSSEub7MXpiudTmWa5PCFgJeWZJ7d5pS3WzNkG8XeWfcVZ+yBF0Tsczp5E9
yoFSjL0bPLdTUr28XzoABZfTeZwhs7gHji7N79qJdxkR7hJP2sCIGaM7i8i/aqxWQWoW7/ou9ELB
nCEPOsztrtfmHOn1/ihW0CTHhVunab3SjdfFy0xU3o6gwq2uHOhjRY+pOt6CUppHOXnFyKnEdo45
Cy15brmqSZSsR/VPevz74wBRkgwZrt8rPIs8nPPSYneul0m76pRsMuC899MMeFi7o9UoUN2rBEQ+
SgG02Yl/L4UGRUdFy4uv/XPBBlMu/cloAXvrKfXSfDe51b7yIPiI8cvBsRveMlEdTz1EC/VnZ6o4
KeAd7dLtjjXwd+ZR9pwfN8CIx+13EcSBtjQRnl/hoNx1MTlaGzkX7L+BC6+BT06XAdLhbOc3O7Sr
FeXgF9ur0IO1bKHPVP91wkY89Ojzfz7X5IMiVOjhASLThUXugyGqwblLMxA8iCw62gBctuGICuUo
MAnnAJ9l+AYxk/KuGSNykX9QJE5tfyi8cKZYuf7OiVbY8DsbX7qRLaWZSdpMuh7VmS94buHtO/B9
2K2e38g2njHrrfgrvizJnW0urJtLakeotJShoF+zLwwFsNLjpXPZmEx0rMB/9A6CcDU1hhNE5fJy
WBeu34yvs4fYaOhQrMifj34jK06GSIyV3OJA33ZK1R94U57WfZP2sr2dINfvBc5wN2RVKATBHoJW
Wy+CrnuwXetp+aWPMR3Ig6nFm6MTzFTc8H2xhRjBRNI/V+k=
`protect end_protected
